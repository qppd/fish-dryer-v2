PK
     uK\���v� �    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47":["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48":["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos"],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62":[],"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos":["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg":["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-pos":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-neg":[],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos"],"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_0":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_1":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_2":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_3":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_4":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_5":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_6":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_7":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_8":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_9":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_10":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_11":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_12":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_13":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_14":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_15":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_16":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_17":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_18":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_19":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_20":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_21":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_22":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_23":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_24":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_25":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_26":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_27":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_28":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_29":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_30":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_31":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_32":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_33":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_34":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_35":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_36":[],"pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_37":[],"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0":["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2"],"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6"],"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2":["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0"],"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0":["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2"],"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5"],"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2":["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0"],"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0":["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2"],"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4"],"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2":["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0"],"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0":["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2"],"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7"],"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2":["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0"],"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"],"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47"],"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2"],"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3":["pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1"],"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"],"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46"],"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2":["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4"],"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3":["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0"],"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"],"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48"],"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2":["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2"],"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3":["pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1"],"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3"],"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1":["pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"],"pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0":["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1"],"pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1":["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3"],"pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0":["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1"],"pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1":["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3"],"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39"],"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg"],"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44"],"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4":["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5":["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6":["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7":["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1"],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_8":[],"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_9":[],"pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_0":[],"pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_1":[],"pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_0":[],"pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_1":[],"pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_0":[],"pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_1":[],"pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_2":[],"pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_3":[],"pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_4":[],"pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_5":[],"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos"],"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg"],"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2":["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"],"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3":["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"],"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_0":[],"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1":["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"],"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2":[],"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3":["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3"],"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4":["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1"],"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0":["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0"],"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1":["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1"],"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2":["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0"],"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3":["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1"],"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_4":[],"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_5":[],"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1":["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0"],"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0":["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1"],"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2":["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1"],"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3":["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"],"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0":["pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"],"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1":["pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"],"pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0":["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0"],"pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1":["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1"],"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0":["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1"],"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1":["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0"],"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0"],"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1"],"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2":["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1"],"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3":["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0"],"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2"],"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3"],"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2":["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1"],"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3":["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0"],"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_0":[],"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1":["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2"],"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2":[],"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3":["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3"],"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2"]},"pin_to_color":{"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33":"#4ab036","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36":"#189AB4","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39":"#ff0000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40":"#4ab036","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41":"#4ab036","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44":"#A75740","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46":"#FF74A3","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47":"#4ab036","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47":"#683D3B","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48":"#FE8900","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48":"#9e007c","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52":"#189AB4","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57":"#FF0000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60":"#189AB4","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61":"#FF0000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62":"#000000","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos":"#FF0000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos":"#FF0000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg":"#189AB4","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos":"#FF0000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-pos":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos":"#FF0000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-neg":"#000000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos":"#FF0000","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_0":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_1":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_2":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_3":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_4":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_5":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_6":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_7":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_8":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_9":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_10":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_11":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_12":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_13":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_14":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_15":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_16":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_17":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_18":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_19":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_20":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_21":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_22":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_23":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_24":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_25":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_26":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_27":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_28":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_29":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_30":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_31":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_32":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_33":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_34":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_35":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_36":"#000000","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_37":"#000000","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0":"#001544","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1":"#f44336","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2":"#95003a","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0":"#95003a","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1":"#f44336","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2":"#001544","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0":"#95003A","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1":"#f44336","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2":"#95003a","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0":"#95003a","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1":"#f44336","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2":"#95003A","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0":"#189AB4","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1":"#683D3B","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2":"#f44336","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3":"#5500bd","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0":"#189AB4","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1":"#FF74A3","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2":"#f44336","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3":"#f238ff","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0":"#189AB4","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1":"#9e007c","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2":"#f44336","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3":"#4ab036","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0":"#f238ff","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1":"#000000","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0":"#000000","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1":"#5500bd","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0":"#000000","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1":"#4ab036","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0":"#ff0000","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1":"#189AB4","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3":"#A75740","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2":"#4ab036","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0":"#189AB4","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1":"#4ab036","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2":"#FE8900","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3":"#ff0000","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4":"#f44336","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5":"#f44336","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6":"#f44336","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7":"#f44336","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_8":"#000000","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_9":"#000000","pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_0":"#000000","pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_1":"#000000","pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_0":"#000000","pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_1":"#000000","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_0":"#000000","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_1":"#000000","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_2":"#000000","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_3":"#000000","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_4":"#000000","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_5":"#000000","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0":"#FF0000","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1":"#189AB4","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2":"#f44336","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3":"#000000","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_0":"#000000","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1":"#f44336","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2":"#000000","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3":"#000000","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4":"#000000","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0":"#f44336","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1":"#000000","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2":"#f44336","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3":"#000000","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_4":"#000000","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_5":"#000000","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1":"#000000","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0":"#f44336","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2":"#f44336","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3":"#000000","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0":"#000000","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1":"#f44336","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0":"#000000","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1":"#f44336","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0":"#000000","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1":"#f44336","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0":"#f44336","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1":"#000000","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2":"#f44336","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3":"#000000","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0":"#f44336","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1":"#000000","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2":"#f44336","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3":"#000000","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_0":"#000000","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1":"#f44336","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2":"#000000","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3":"#000000","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4":"#f44336"},"pin_to_state":{"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62":"neutral","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-neg":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos":"neutral","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_0":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_1":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_2":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_3":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_4":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_5":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_6":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_7":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_8":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_9":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_10":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_11":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_12":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_13":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_14":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_15":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_16":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_17":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_18":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_19":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_20":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_21":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_22":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_23":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_24":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_25":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_26":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_27":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_28":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_29":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_30":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_31":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_32":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_33":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_34":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_35":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_36":"neutral","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_37":"neutral","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0":"neutral","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1":"neutral","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2":"neutral","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0":"neutral","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1":"neutral","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2":"neutral","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0":"neutral","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1":"neutral","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2":"neutral","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0":"neutral","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1":"neutral","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2":"neutral","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0":"neutral","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1":"neutral","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2":"neutral","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3":"neutral","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0":"neutral","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1":"neutral","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2":"neutral","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3":"neutral","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0":"neutral","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1":"neutral","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2":"neutral","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3":"neutral","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0":"neutral","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1":"neutral","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0":"neutral","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1":"neutral","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0":"neutral","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1":"neutral","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0":"neutral","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1":"neutral","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3":"neutral","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_8":"neutral","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_9":"neutral","pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_0":"neutral","pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_1":"neutral","pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_0":"neutral","pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_1":"neutral","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_0":"neutral","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_1":"neutral","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_2":"neutral","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_3":"neutral","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_4":"neutral","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_5":"neutral","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0":"neutral","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1":"neutral","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2":"neutral","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3":"neutral","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_0":"neutral","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1":"neutral","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2":"neutral","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3":"neutral","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4":"neutral","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0":"neutral","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1":"neutral","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2":"neutral","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3":"neutral","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_4":"neutral","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_5":"neutral","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1":"neutral","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0":"neutral","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2":"neutral","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3":"neutral","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0":"neutral","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1":"neutral","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0":"neutral","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1":"neutral","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0":"neutral","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1":"neutral","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0":"neutral","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1":"neutral","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2":"neutral","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3":"neutral","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0":"neutral","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1":"neutral","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2":"neutral","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3":"neutral","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_0":"neutral","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1":"neutral","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2":"neutral","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3":"neutral","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4":"neutral"},"next_color_idx":4,"wires_placed_in_order":[["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4"],["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5"],["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6"],["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7"],["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0"],["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0"],["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0"],["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0"],["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41"],["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44"],["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0"],["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg"],["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41"],["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3"],["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47"],["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48"],["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1"],["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos"],["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos"],["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_0","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_1","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2"],["pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0"],["pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1"],["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"],["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"],["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1"],["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0"],["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"],["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"],["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1"],["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0"],["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0"],["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1"],["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1"],["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0"],["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1"],["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0"],["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2"],["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2"],["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2"],["pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"],["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"],["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2"],["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"],["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1"],["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3"],["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"],["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"],["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3"],["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2"],["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4"]]],[[],[["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5"]]],[[],[["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6"]]],[[],[["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7"]]],[[],[["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0"]]],[[],[["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0"]]],[[],[["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0"]]],[[],[["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0"]]],[[],[["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"]]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos"]]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg"]]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos"]],[]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"]],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33"]]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"]]],[[],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg"]]],[[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg"]],[]],[[],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0"]]],[[],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41"]]],[[],[["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44"]]],[[],[["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"]]],[[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"]]],[[["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg"]],[]],[[["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg"]],[]],[[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg"]],[]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"]]],[[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"]],[]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"]]],[[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg"]],[]],[[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"]],[]],[[],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0"]]],[[],[["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg"]]],[[],[["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41"]]],[[],[["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44"]]],[[["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos"]],[]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3"]]],[[],[["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47"]]],[[],[["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48"]]],[[],[["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1"]]],[[],[["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1"]]],[[],[["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3"]]],[[],[["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3"]]],[[],[["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0"]]],[[],[["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0"]]],[[],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2"]]],[[],[["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2"]]],[[],[["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2"]]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos"]]],[[],[["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg"]]],[[],[]],[[],[]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos"]]],[[],[["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg"]]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos"]]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg"]]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1"]]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3"]]],[[],[["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_0","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"]]],[[],[["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_1","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2"]]],[[],[["pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0"]]],[[],[["pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1"]]],[[],[["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"]]],[[],[["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"]]],[[],[["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1"]]],[[],[["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0"]]],[[["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"]],[]],[[["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"]],[]],[[],[["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"]]],[[],[["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"]]],[[["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1"]],[]],[[["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0"]],[]],[[],[["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1"]]],[[],[["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0"]]],[[],[["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0"]]],[[],[["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1"]]],[[],[["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1"]]],[[],[["pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0"]]],[[],[["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1"]]],[[],[["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0"]]],[[],[["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2"]]],[[],[["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3"]]],[[["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_1"]],[]],[[["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_0"]],[]],[[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3"]],[]],[[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1"]],[]],[[["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"]],[]],[[["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2"]],[]],[[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2"],["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2"],["pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2"]],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2"],["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2"]]],[[["pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3"],["pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0","pin-type-component_db3cd3e2-6bf6-4358-bf0c-9697139ac262_3"]],[["pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1"],["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0"]]],[[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg"]],[]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg"]]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"]]],[[],[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"]]],[[],[["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2"]]],[[],[["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"]]],[[],[["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1"]]],[[],[["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3"]]],[[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"]],[]],[[["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"]],[]],[[["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"]],[]],[[["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2"]],[]],[[],[["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3"]]],[[],[["pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1"]]],[[],[["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3"]]],[[],[["pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2"]]],[[],[["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4"]]],[[],[["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2"]]],[[["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2"]],[]],[[],[["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33":"0000000000000010","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36":"0000000000000011","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39":"0000000000000018","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40":"0000000000000010","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41":"0000000000000020","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44":"0000000000000021","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46":"0000000000000015","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47":"0000000000000009","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47":"0000000000000016","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48":"0000000000000022","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48":"0000000000000017","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52":"0000000000000029","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57":"0000000000000028","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60":"0000000000000012","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61":"0000000000000013","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62":"_","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg":"0000000000000031","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg":"0000000000000031","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_1_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos":"0000000000000032","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_2_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_2_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_3_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg":"0000000000000033","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_4_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_4_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_5_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_5_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_6_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_6_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_7_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_7_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_8_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_8_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_9_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_9_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_10_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_10_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_11_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_11_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_12_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_12_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_13_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_13_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_14_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_14_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_15_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_15_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_16_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_16_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_17_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_17_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_18_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_18_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_19_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_19_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_20_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_20_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_21_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_21_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_22_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_22_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_23_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_23_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_24_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_24_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_25_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_25_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_26_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_26_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_27_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_27_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_28_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_28_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_29_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_29_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_30_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_30_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_31_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg":"0000000000000014","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_32_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_32_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_33_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_34_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_34_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_35_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_35_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg":"0000000000000011","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_36_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg":"0000000000000019","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_37_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_38_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_38_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_39_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_40_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_41_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_42_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_42_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_43_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_43_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_44_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_45_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_45_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_46_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_49_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_49_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg":"0000000000000008","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_50_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_51_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_51_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg":"0000000000000029","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_52_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_53_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_53_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_54_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_54_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_55_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_55_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_56_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_56_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos":"0000000000000028","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_57_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_58_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_58_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_59_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_59_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg":"0000000000000012","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_60_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos":"0000000000000013","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-pos":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_61_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos":"0000000000000030","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-neg":"_","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos":"0000000000000030","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-neg":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_0":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_1":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_2":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_3":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_4":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_5":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_6":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_7":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_8":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_9":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_10":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_11":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_12":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_13":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_14":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_15":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_16":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_17":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_18":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_19":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_20":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_21":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_22":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_23":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_24":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_25":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_26":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_27":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_28":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_29":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_30":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_31":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_32":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_33":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_34":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_35":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_36":"_","pin-type-component_721d3748-6859-4a91-8f48-309f28334d2f_37":"_","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0":"0000000000000007","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1":"0000000000000002","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2":"0000000000000004","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0":"0000000000000006","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1":"0000000000000001","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2":"0000000000000007","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0":"0000000000000005","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1":"0000000000000000","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2":"0000000000000006","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0":"0000000000000004","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1":"0000000000000003","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2":"0000000000000005","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0":"0000000000000014","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1":"0000000000000016","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2":"0000000000000027","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3":"0000000000000024","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0":"0000000000000014","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1":"0000000000000015","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2":"0000000000000027","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3":"0000000000000025","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0":"0000000000000014","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1":"0000000000000017","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2":"0000000000000027","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3":"0000000000000023","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0":"0000000000000025","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1":"0000000000000026","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0":"0000000000000026","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1":"0000000000000024","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0":"0000000000000026","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1":"0000000000000023","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0":"0000000000000018","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1":"0000000000000019","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3":"0000000000000021","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2":"0000000000000020","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0":"0000000000000008","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1":"0000000000000009","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2":"0000000000000022","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3":"0000000000000018","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4":"0000000000000000","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5":"0000000000000001","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6":"0000000000000002","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7":"0000000000000003","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_8":"_","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_9":"_","pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_0":"_","pin-type-component_96e3621c-0323-4781-8b4e-eb33eb2c0fd1_1":"_","pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_0":"_","pin-type-component_396b3281-51bc-4ef3-ac9d-b618930e84e2_1":"_","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_0":"_","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_1":"_","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_2":"_","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_3":"_","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_4":"_","pin-type-component_0cc31a1e-63f6-41c8-b821-f4c6defad7b6_5":"_","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0":"0000000000000032","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1":"0000000000000033","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2":"0000000000000046","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3":"0000000000000047","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_0":"_","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1":"0000000000000046","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_2":"_","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3":"0000000000000047","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4":"0000000000000026","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0":"0000000000000041","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1":"0000000000000040","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2":"0000000000000042","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3":"0000000000000043","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_4":"_","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_5":"_","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1":"0000000000000045","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0":"0000000000000044","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2":"0000000000000046","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3":"0000000000000047","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0":"0000000000000038","pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1":"0000000000000039","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0":"0000000000000038","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1":"0000000000000039","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0":"0000000000000045","pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1":"0000000000000044","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0":"0000000000000041","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1":"0000000000000040","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2":"0000000000000039","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3":"0000000000000038","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0":"0000000000000042","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1":"0000000000000043","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2":"0000000000000044","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3":"0000000000000045","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_0":"_","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1":"0000000000000046","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_2":"_","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3":"0000000000000047","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4":"0000000000000027"},"component_id_to_pins":{"721d3748-6859-4a91-8f48-309f28334d2f":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"d5434b8f-b5c1-4202-b31f-205d8ac815b6":["0","1","2"],"4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b":["0","1","2"],"17bf28ad-c945-4b6f-bda0-e3fe826ab5a9":["0","1","2"],"e0564417-360a-4149-877f-c52809d9ef28":["0","1","2"],"cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b":["0","1","2","3"],"84de52eb-d97f-4432-8888-452b5250f3c1":["0","1","2","3"],"fa11e16a-f0a7-42e2-a7d4-599f2d603b47":["0","1","2","3"],"6d2add11-c610-441d-abbc-fd8eae0f97b2":["0","1"],"6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687":["0","1"],"c80f0ed6-f74d-456d-a629-db513543e96f":["0","1"],"50b4d32c-e906-420a-abe1-aa498357d8ae":["0","1","3","2"],"544cf99b-406e-4351-9364-3825fb8135d0":["0","1","2","3","4","5","6","7","8","9"],"96e3621c-0323-4781-8b4e-eb33eb2c0fd1":["0","1"],"396b3281-51bc-4ef3-ac9d-b618930e84e2":["0","1"],"0cc31a1e-63f6-41c8-b821-f4c6defad7b6":["0","1","2","3","4","5"],"390d83ab-07c8-4d04-99d0-82df7aff116b":["0","1","2","3"],"bcf76462-cf56-4f01-b598-ae1e6dd3ec4d":["0","1","2","3","4"],"49c909aa-82cc-42de-ad47-eeb2d04e532b":["0","1","2","3","4","5"],"1ac7d52d-b253-412f-8e1b-4251a9594a23":["1","0","2","3"],"6203bc03-c8ad-4e65-acf1-0957e7d9561a":["0","1"],"7821f33a-bdac-4457-86e4-7ce6064f4871":["0","1"],"6f68e686-1c6d-45e3-a7d6-9788c0bfcfab":["0","1"],"86163d73-1a9c-44b6-a2e1-728e256546df":["0","1","2","3"],"af79f859-314d-4925-8469-848813fd14e6":["0","1","2","3"],"a669ed33-4ae7-4630-b33a-1a8d6006ac36":["0","1","2","3","4"],"fdbea0e9-0786-4f33-9e71-8223031661f6":[],"3706761d-9ca2-45cb-864d-520bef03d29f":[],"06ef71ab-6201-4d71-85ff-63ce83357255":[],"d547533d-d7a0-4185-8985-c0fa1c7271c6":[],"625549d8-f708-4010-ab04-318947e6dc81":[],"ce78d232-d380-4a7f-bfad-f5f98270dc96":[],"a7cb9edb-11e3-43c3-8685-97b305969503":[],"9943bd98-399b-4f38-b938-9ddf715b5998":[],"3d2b088b-f2fd-4ce4-bc73-c68faea65f47":[],"c43bcff6-4422-4f0e-ac52-68d069eea4af":[],"a029f855-aaba-41f9-aa2c-7695dbb49691":[],"82685ae2-a134-4e77-b2c6-b1b7eff37783":[],"50246903-644b-49bf-b5eb-24c7cecfc97b":[]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4"],"0000000000000001":["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5"],"0000000000000002":["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6"],"0000000000000003":["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7"],"0000000000000004":["pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2","pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0"],"0000000000000005":["pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2","pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0"],"0000000000000006":["pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2","pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0"],"0000000000000007":["pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2","pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0"],"0000000000000008":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0"],"0000000000000012":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg"],"0000000000000013":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos"],"0000000000000010":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33"],"0000000000000011":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg"],"0000000000000017":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1"],"0000000000000016":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1"],"0000000000000015":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1"],"0000000000000014":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0"],"0000000000000018":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39","pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0","pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3"],"0000000000000019":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg"],"0000000000000020":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41"],"0000000000000021":["pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44"],"0000000000000009":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47"],"0000000000000022":["pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2","pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48"],"0000000000000023":["pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1"],"0000000000000024":["pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3","pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1"],"0000000000000025":["pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0","pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3"],"0000000000000026":["pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0","pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1","pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4"],"0000000000000027":["pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2","pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2","pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4"],"0000000000000028":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos"],"0000000000000029":["pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg"],"0000000000000030":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos"],"0000000000000031":["pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg"],"0000000000000032":["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos"],"0000000000000038":["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3"],"0000000000000039":["pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1","pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2"],"0000000000000040":["pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1","pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1"],"0000000000000041":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0","pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0"],"0000000000000042":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0"],"0000000000000043":["pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1"],"0000000000000044":["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0"],"0000000000000045":["pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0","pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3","pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1"],"0000000000000033":["pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1","pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg"],"0000000000000046":["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2"],"0000000000000047":["pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3","pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3","pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3","pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000017":"Net 17","0000000000000016":"Net 16","0000000000000015":"Net 15","0000000000000014":"Net 14","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000021":"Net 21","0000000000000009":"Net 9","0000000000000022":"Net 22","0000000000000023":"Net 23","0000000000000024":"Net 24","0000000000000025":"Net 25","0000000000000026":"Net 26","0000000000000027":"Net 27","0000000000000028":"Net 28","0000000000000029":"Net 29","0000000000000030":"Net 30","0000000000000031":"Net 31","0000000000000032":"Net 32","0000000000000038":"Net 38","0000000000000039":"Net 39","0000000000000040":"Net 40","0000000000000041":"Net 41","0000000000000042":"Net 42","0000000000000043":"Net 43","0000000000000044":"Net 44","0000000000000045":"Net 45","0000000000000033":"Net 33","0000000000000046":"Net 46","0000000000000047":"Net 47"},"all_breadboard_info_list":["b62302e1-db31-40ba-a2dc-d3556ee2692c_63_2_True_715_820_up"],"breadboard_info_list":["b62302e1-db31-40ba-a2dc-d3556ee2692c_63_2_True_715_820_up"],"componentsData":[{"compProperties":{},"position":[757.689823,1563.6117905],"typeId":"69c262f4-fa86-6b73-0b2d-129f230d5ed6","componentVersion":3,"instanceId":"721d3748-6859-4a91-8f48-309f28334d2f","orientation":"up","circleData":[[692.5,1415],[692.5,1430],[692.5,1445],[692.5,1460],[692.5,1475.0000000000002],[692.5,1490.0000000000002],[692.5,1505.0000000000002],[692.5,1520.0000000000002],[692.5,1535.0000000000002],[692.5,1550.0000000000002],[692.5,1565],[692.5,1580],[692.5,1595],[692.5,1610],[692.5,1625],[692.5,1640],[692.5,1655],[692.5,1670],[692.5,1685],[827.5,1685],[827.5,1670],[827.5,1655],[827.5,1640],[827.5,1625],[827.5,1610],[827.5,1595],[827.5,1580],[827.5,1565],[827.5,1550.0000000000002],[827.5,1535.0000000000002],[827.5,1520.0000000000002],[827.5,1505.0000000000002],[827.5,1490.0000000000002],[827.5,1475.0000000000002],[827.5,1460],[827.5,1445],[827.5,1430],[827.5,1415]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-105.18448250000006,1738.5675005000003],"typeId":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"instanceId":"d5434b8f-b5c1-4202-b31f-205d8ac815b6","orientation":"right","circleData":[[-27.499999999999986,1729.9999999999998],[-28.928000000000097,1741.4239999999998],[-29.64200000000004,1753.562]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[53.93249950000016,1397.3155175000002],"typeId":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"instanceId":"17bf28ad-c945-4b6f-bda0-e3fe826ab5a9","orientation":"down","circleData":[[62.500000000000014,1475],[51.07600000000005,1473.572],[38.93800000000013,1472.858]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[56.06750049999998,1882.6844825],"typeId":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"instanceId":"e0564417-360a-4149-877f-c52809d9ef28","orientation":"up","circleData":[[47.499999999999986,1805],[58.92399999999995,1806.428],[71.06200000000001,1807.142]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1215.3179995,1728.5505005],"typeId":"b97d5804-295d-4a63-b66d-23cafcd44586","componentVersion":2,"instanceId":"cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b","orientation":"right","circleData":[[1067.5,1640],[1068.676,1814.0945],[1359.226,1636.4705000000001],[1359.226,1814.0944999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1215.3179995000005,1383.5505005],"typeId":"b97d5804-295d-4a63-b66d-23cafcd44586","componentVersion":2,"instanceId":"84de52eb-d97f-4432-8888-452b5250f3c1","orientation":"right","circleData":[[1067.5,1295],[1068.6759999999995,1469.0944999999997],[1359.2260000000003,1291.4705],[1359.2260000000003,1469.0944999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1215.3179995,2073.5505005000005],"typeId":"b97d5804-295d-4a63-b66d-23cafcd44586","componentVersion":2,"instanceId":"fa11e16a-f0a7-42e2-a7d4-599f2d603b47","orientation":"right","circleData":[[1067.5,1985],[1068.6760000000002,2159.0945000000006],[1359.226,1981.4705],[1359.2260000000003,2159.0945000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[393.99637299999995,1368.943631],"typeId":"01534432-bd5d-4550-957a-0d4278d98851","componentVersion":1,"instanceId":"50b4d32c-e906-420a-abe1-aa498357d8ae","orientation":"left","circleData":[[467.5,1415],[468.7592679999998,1384.073114],[466.24073050000015,1319.422262],[468.7592679999998,1349.0898815]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[274.5540309999999,1634.5455005000001],"typeId":"8f8ecf0b-b7ef-4a48-962c-7614bb5a7d82","componentVersion":1,"instanceId":"544cf99b-406e-4351-9364-3825fb8135d0","orientation":"right","circleData":[[362.5,1610],[362.27199999999993,1628.9180000000001],[362.9469999999999,1646.9915],[362.27199999999993,1664.39],[181.73649999999992,1592.1200000000001],[181.9194999999999,1610.5880000000002],[181.73649999999992,1628.987],[181.59999999999985,1647.3185000000003],[181.74099999999993,1665.1040000000003],[181.74099999999993,1683.9785000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1746.6718420000007,1352.7273304999999],"typeId":"1255ec18-62c0-4252-8215-c2ff45234b02","componentVersion":1,"instanceId":"6d2add11-c610-441d-abbc-fd8eae0f97b2","orientation":"right","circleData":[[1562.5,1310],[1564.0075000000002,1424.4904999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1713.3377770000006,2067.3988714999996],"typeId":"6635379e-9371-f184-7e48-a00d3644b40e","componentVersion":1,"instanceId":"c80f0ed6-f74d-456d-a629-db513543e96f","orientation":"up","circleData":[[1562.5,2180],[1562.552413,2166.733166]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-105.18448250000006,1558.5675005],"typeId":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"instanceId":"4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b","orientation":"right","circleData":[[-27.500000000000014,1550],[-28.928000000000125,1561.424],[-29.642000000000067,1573.5620000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"version":2,"id":"Capacitance","label":"Capacitance","description":"","units":"F","type":"decimal","value":"0.000001","displayFormat":"input","showOnComp":true,"isVisibleToUser":true,"name":"Capacitance","unit":"F","required":true}},"position":[794.6995,1737.4295],"typeId":"14d7a2a7-6581-4d0a-a495-63cc6355f7b9","componentVersion":1,"instanceId":"96e3621c-0323-4781-8b4e-eb33eb2c0fd1","orientation":"right","circleData":[[737.5,1730],[737.5,1745]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[722.4885565,1347.074954],"typeId":"02adc9af-9099-49f0-8d17-97b22a4179bc","componentVersion":1,"instanceId":"396b3281-51bc-4ef3-ac9d-b618930e84e2","orientation":"up","circleData":[[722.5,1325],[722.5,1370]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[769.2245245,1613.069966],"typeId":"84de3699-1b7e-4fcb-b51f-13b7bf5839ea","componentVersion":1,"instanceId":"0cc31a1e-63f6-41c8-b821-f4c6defad7b6","orientation":"up","circleData":[[812.5,1625],[812.158,1613.03],[812.158,1600.034],[748.543,1597.298],[748.885,1612.346],[749.227,1627.736]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1195,972.5],"typeId":"c16bfa02-5154-4f39-9ff1-d473663907f3","componentVersion":2,"instanceId":"390d83ab-07c8-4d04-99d0-82df7aff116b","orientation":"left","circleData":[[1157.5,1130],[1172.5,1130],[1345.0000000000005,958.6010000000001],[1345.0000000000005,886.2725]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1784.135347,1005.4810880000002],"typeId":"ef0da927-5348-4d94-b21a-42d8a46ff031","componentVersion":1,"instanceId":"bcf76462-cf56-4f01-b598-ae1e6dd3ec4d","orientation":"up","circleData":[[1712.5,1130],[1858.072,921.1925000000003],[1858.072,1074.6695],[1712.3964999999998,923.7920000000004],[1713.0565,1075.9520000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[221.8501419999998,842.5139749999992],"typeId":"aec5eff0-da06-45e7-8932-95bc26fc4e6a","componentVersion":1,"instanceId":"6203bc03-c8ad-4e65-acf1-0957e7d9561a","orientation":"up","circleData":[[32.50000000000003,1070],[32.50000000000003,1052.3166394999992]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1147.3543435,604.5910745000001],"typeId":"8903b643-ed64-43f6-b56c-46542b1c2184","componentVersion":2,"instanceId":"6f68e686-1c6d-45e3-a7d6-9788c0bfcfab","orientation":"up","circleData":[[1052.5,515],[1247.5000000000007,515]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[653.318041,548.0942735000001],"typeId":"023546b5-ca70-49d6-8fe2-6f4e8641da15","componentVersion":1,"instanceId":"86163d73-1a9c-44b6-a2e1-728e256546df","orientation":"up","circleData":[[617.5,425],[687.501715,421.7864495000001],[616.0660345,674.6406499999999],[691.0660345,674.6406499999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[221.85014200000015,77.51397499999962],"typeId":"aec5eff0-da06-45e7-8932-95bc26fc4e6a","componentVersion":1,"instanceId":"7821f33a-bdac-4457-86e4-7ce6064f4871","orientation":"up","circleData":[[32.5,305],[32.5,287.31663949999984]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[725.2929999999994,-84.4869999999998],"typeId":"28def945-d566-45d1-91c0-cb2676c61db2","componentVersion":1,"instanceId":"49c909aa-82cc-42de-ad47-eeb2d04e532b","orientation":"up","circleData":[[632.5,185],[671.2060000000001,183.82699999999977],[708.7404999999999,182.654],[745.1020000000001,182.654],[782.6365000000003,183.82699999999977],[817.8250000000005,183.82699999999977]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1186.140895,127.54614349999954],"typeId":"b8a657e4-3f8b-4e3e-a2bd-792a2961387f","componentVersion":1,"instanceId":"1ac7d52d-b253-412f-8e1b-4251a9594a23","orientation":"left","circleData":[[1247.5,320],[1127.6169265,320],[1139.5935415000001,-71.10244900000015],[1229.6770600000002,-71.10244900000015]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[848.3180410000002,548.0942735000002],"typeId":"023546b5-ca70-49d6-8fe2-6f4e8641da15","componentVersion":1,"instanceId":"af79f859-314d-4925-8469-848813fd14e6","orientation":"up","circleData":[[812.5,425],[882.501715,421.7864495000001],[811.0660345,674.6406499999998],[886.0660345,674.6406499999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1514.135347,1005.4810879999998],"typeId":"ef0da927-5348-4d94-b21a-42d8a46ff031","componentVersion":1,"instanceId":"a669ed33-4ae7-4630-b33a-1a8d6006ac36","orientation":"up","circleData":[[1442.5,1130],[1588.072,921.1924999999999],[1588.072,1074.6695],[1442.3964999999998,923.7919999999999],[1443.0565,1075.9520000000002]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1713.337777,1707.3988715],"typeId":"6635379e-9371-f184-7e48-a00d3644b40e","componentVersion":1,"instanceId":"6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687","orientation":"up","circleData":[[1562.5,1820],[1562.552413,1806.733166]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"HX711 ","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[271.89804429448094,1753.8900165443397],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"fdbea0e9-0786-4f33-9e71-8223031661f6","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"SHT31","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[397.26190713707956,1489.00097505186],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"3706761d-9ca2-45cb-864d-520bef03d29f","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"12V to 220V \nINVERTER","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1524.050996846438,168.51815453606454],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"06ef71ab-6201-4d71-85ff-63ce83357255","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LiFePo4 \nBATTERY","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1480.677587609787,618.3601797117985],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"d547533d-d7a0-4185-8985-c0fa1c7271c6","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"SOLID STATE RELAY","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1217.868024263463,2267.0705892494416],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"625549d8-f708-4010-ab04-318947e6dc81","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"FAN","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1715.1106813093047,2261.255549878445],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"ce78d232-d380-4a7f-bfad-f5f98270dc96","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"HEATING ELEMENT","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[1757.8089561050558,1489.0573946319537],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"a7cb9edb-11e3-43c3-8685-97b305969503","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOADCELL","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[-26.266679526276505,2016.3138501112107],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"9943bd98-399b-4f38-b938-9ddf715b5998","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"SOLAR PANEL","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[227.43862145758555,-280.3219899869995],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"3d2b088b-f2fd-4ce4-bc73-c68faea65f47","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"SOLAR CHARGE\nCONTROLLER","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[729.3613045369607,-458.7345396378521],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"c43bcff6-4422-4f0e-ac52-68d069eea4af","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"DC BREAKER","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[748.1847473668196,750.7076396004542],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"a029f855-aaba-41f9-aa2c-7695dbb49691","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"BUZZER","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[846.4716786236559,1347.4074421060718],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"82685ae2-a134-4e77-b2c6-b1b7eff37783","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"ESP32","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"0.1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"textColor":{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"fontSize":{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"40","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},"font":{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}},"position":[758.672946257867,1505.5426587423865],"typeId":"9a5a4baa-44d4-4aa0-8d82-488487322b20","componentVersion":1,"instanceId":"50246903-644b-49bf-b5eb-24c7cecfc97b","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-516.73454","left":"-194.42978","width":"2143.67429","height":"2836.30513","x":"-194.42978","y":"-516.73454"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1\",\"endPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4\",\"rawStartPinId\":\"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_1\",\"rawEndPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"51.0760000000_1473.5720000000\\\",\\\"51.0760000000_1592.1200000000\\\",\\\"181.7365000000_1592.1200000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1\",\"endPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5\",\"rawStartPinId\":\"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_1\",\"rawEndPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-28.9280000000_1561.4240000000\\\",\\\"40.0000000000_1561.4240000000\\\",\\\"40.0000000000_1610.0000000000\\\",\\\"181.9195000000_1610.0000000000\\\",\\\"181.9195000000_1610.5880000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6\",\"endPinId\":\"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1\",\"rawStartPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_6\",\"rawEndPinId\":\"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"181.7365000000_1628.9870000000\\\",\\\"40.0000000000_1628.9870000000\\\",\\\"40.0000000000_1745.0000000000\\\",\\\"-28.9280000000_1745.0000000000\\\",\\\"-28.9280000000_1741.4240000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7\",\"endPinId\":\"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1\",\"rawStartPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_7\",\"rawEndPinId\":\"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"181.6000000000_1647.3185000000\\\",\\\"55.0000000000_1647.3185000000\\\",\\\"55.0000000000_1726.8732500000\\\",\\\"62.5000000000_1726.8732500000\\\",\\\"62.5000000000_1806.4280000000\\\",\\\"58.9240000000_1806.4280000000\\\"]}\"}","{\"color\":\"#95003a\",\"startPinId\":\"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2\",\"endPinId\":\"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0\",\"rawStartPinId\":\"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_2\",\"rawEndPinId\":\"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-29.6420000000_1753.5620000000\\\",\\\"47.5000000000_1753.5620000000\\\",\\\"47.5000000000_1805.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0\",\"endPinId\":\"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2\",\"rawStartPinId\":\"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_0\",\"rawEndPinId\":\"pin-type-component_e0564417-360a-4149-877f-c52809d9ef28_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"62.5000000000_1475.0000000000\\\",\\\"62.5000000000_1640.0000000000\\\",\\\"71.0620000000_1640.0000000000\\\",\\\"71.0620000000_1807.1420000000\\\"]}\"}","{\"color\":\"#95003a\",\"startPinId\":\"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2\",\"endPinId\":\"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0\",\"rawStartPinId\":\"pin-type-component_17bf28ad-c945-4b6f-bda0-e3fe826ab5a9_2\",\"rawEndPinId\":\"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"38.9380000000_1472.8580000000\\\",\\\"38.9380000000_1550.0000000000\\\",\\\"-27.5000000000_1550.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2\",\"endPinId\":\"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0\",\"rawStartPinId\":\"pin-type-component_4d4d56f8-ba1e-4a1b-a966-759bdbf2d56b_2\",\"rawEndPinId\":\"pin-type-component_d5434b8f-b5c1-4202-b31f-205d8ac815b6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-29.6420000000_1573.5620000000\\\",\\\"-12.5000000000_1573.5620000000\\\",\\\"-12.5000000000_1730.0000000000\\\",\\\"-27.5000000000_1730.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg\",\"rawStartPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_50_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"362.5000000000_1610.0000000000\\\",\\\"422.5000000000_1610.0000000000\\\",\\\"422.5000000000_1580.0000000000\\\",\\\"632.5000000000_1580.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_60_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1730.0000000000\\\",\\\"632.5000000000_1730.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_61_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1745.0000000000\\\",\\\"617.5000000000_1745.0000000000\\\"]}\"}","{\"color\":\"#4ab036\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33\",\"endPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_33_0\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_40_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1325.0000000000\\\",\\\"677.5000000000_1310.0000000000\\\",\\\"932.5000000000_1310.0000000000\\\",\\\"932.5000000000_1430.0000000000\\\",\\\"842.5000000000_1430.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_36_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1370.0000000000\\\",\\\"632.5000000000_1370.0000000000\\\"]}\"}","{\"color\":\"#9e007c\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48\",\"endPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_48_4\",\"rawEndPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_1550.0000000000\\\",\\\"977.5000000000_1550.0000000000\\\",\\\"977.5000000000_2159.0945000000\\\",\\\"1068.6760000000_2159.0945000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47\",\"endPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_47_4\",\"rawEndPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_1535.0000000000\\\",\\\"992.5000000000_1535.0000000000\\\",\\\"992.5000000000_1814.0945000000\\\",\\\"1068.6760000000_1814.0945000000\\\"]}\"}","{\"color\":\"#FF74A3\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46\",\"endPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_46_4\",\"rawEndPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_1520.0000000000\\\",\\\"992.5000000000_1520.0000000000\\\",\\\"992.5000000000_1469.0945000000\\\",\\\"1068.6760000000_1469.0945000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg\",\"rawStartPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1067.5000000000_1295.0000000000\\\",\\\"902.5000000000_1295.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg\",\"rawStartPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1067.5000000000_1640.0000000000\\\",\\\"1007.5000000000_1640.0000000000\\\",\\\"1007.5000000000_1295.0000000000\\\",\\\"902.5000000000_1295.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg\",\"rawStartPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_31_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1067.5000000000_1985.0000000000\\\",\\\"1007.5000000000_1985.0000000000\\\",\\\"1007.5000000000_1295.0000000000\\\",\\\"902.5000000000_1295.0000000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39\",\"endPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_0\",\"rawEndPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1415.0000000000\\\",\\\"467.5000000000_1415.0000000000\\\"]}\"}","{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39\",\"endPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_39_0\",\"rawEndPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1415.0000000000\\\",\\\"580.0000000000_1415.0000000000\\\",\\\"580.0000000000_1664.3900000000\\\",\\\"362.2720000000_1664.3900000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg\",\"rawStartPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_1\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_37_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"468.7592680000_1384.0731140000\\\",\\\"497.5000000000_1384.0731140000\\\",\\\"497.5000000000_1385.0000000000\\\",\\\"632.5000000000_1385.0000000000\\\"]}\"}","{\"color\":\"#4ab036\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41\",\"endPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_41_4\",\"rawEndPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_1445.0000000000\\\",\\\"947.5000000000_1445.0000000000\\\",\\\"947.5000000000_1280.0000000000\\\",\\\"580.0000000000_1280.0000000000\\\",\\\"580.0000000000_1349.0898815000\\\",\\\"468.7592680000_1349.0898815000\\\"]}\"}","{\"color\":\"#A75740\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44\",\"endPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_44_4\",\"rawEndPinId\":\"pin-type-component_50b4d32c-e906-420a-abe1-aa498357d8ae_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_1490.0000000000\\\",\\\"962.5000000000_1490.0000000000\\\",\\\"962.5000000000_1265.0000000000\\\",\\\"557.5000000000_1265.0000000000\\\",\\\"557.5000000000_1319.4222620000\\\",\\\"466.2407305000_1319.4222620000\\\"]}\"}","{\"color\":\"#4ab036\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47\",\"endPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_47_0\",\"rawEndPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1535.0000000000\\\",\\\"557.5000000000_1535.0000000000\\\",\\\"557.5000000000_1628.9180000000\\\",\\\"362.2720000000_1628.9180000000\\\"]}\"}","{\"color\":\"#FE8900\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48\",\"endPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_48_0\",\"rawEndPinId\":\"pin-type-component_544cf99b-406e-4351-9364-3825fb8135d0_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1550.0000000000\\\",\\\"535.0000000000_1550.0000000000\\\",\\\"535.0000000000_1646.9915000000\\\",\\\"362.9470000000_1646.9915000000\\\"]}\"}","{\"color\":\"#4ab036\",\"startPinId\":\"pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1\",\"endPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3\",\"rawStartPinId\":\"pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_1\",\"rawEndPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5524130000_2166.7331660000\\\",\\\"1517.5000000000_2166.7331660000\\\",\\\"1517.5000000000_2159.0945000000\\\",\\\"1359.2260000000_2159.0945000000\\\"]}\"}","{\"color\":\"#5500bd\",\"startPinId\":\"pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1\",\"endPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3\",\"rawStartPinId\":\"pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_1\",\"rawEndPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5524130000_1806.7331660000\\\",\\\"1562.5524130000_1805.0000000000\\\",\\\"1517.5000000000_1805.0000000000\\\",\\\"1517.5000000000_1814.0945000000\\\",\\\"1359.2260000000_1814.0945000000\\\"]}\"}","{\"color\":\"#f238ff\",\"startPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0\",\"endPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3\",\"rawStartPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_0\",\"rawEndPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5000000000_1310.0000000000\\\",\\\"1465.0000000000_1310.0000000000\\\",\\\"1465.0000000000_1469.0945000000\\\",\\\"1359.2260000000_1469.0945000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_57_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1685.0000000000\\\",\\\"617.5000000000_1685.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_52_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"677.5000000000_1610.0000000000\\\",\\\"632.5000000000_1610.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos\",\"rawStartPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_62_polarity-pos\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_62_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_1760.0000000000\\\",\\\"887.5000000000_1760.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_0_0_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"632.5000000000_830.0000000000\\\",\\\"902.5000000000_830.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos\",\"rawStartPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_0\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_1_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1157.5000000000_1130.0000000000\\\",\\\"1157.5000000000_1160.0000000000\\\",\\\"1000.0000000000_1160.0000000000\\\",\\\"1000.0000000000_845.0000000000\\\",\\\"887.5000000000_845.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0\",\"endPinId\":\"pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0\",\"rawStartPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0\",\"rawEndPinId\":\"pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"32.5000000000_1070.0000000000\\\",\\\"-57.5000000000_1070.0000000000\\\",\\\"-57.5000000000_1235.0000000000\\\",\\\"572.5000000000_1235.0000000000\\\",\\\"572.5000000000_770.0000000000\\\",\\\"512.5000000000_770.0000000000\\\",\\\"512.5000000000_477.5000000000\\\",\\\"-57.5000000000_477.5000000000\\\",\\\"-57.5000000000_305.0000000000\\\",\\\"32.5000000000_305.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0\",\"endPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3\",\"rawStartPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_0\",\"rawEndPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"32.5000000000_1070.0000000000\\\",\\\"-57.5000000000_1070.0000000000\\\",\\\"-57.5000000000_1235.0000000000\\\",\\\"572.5000000000_1235.0000000000\\\",\\\"572.5000000000_770.0000000000\\\",\\\"691.0660345000_770.0000000000\\\",\\\"691.0660345000_674.6406500000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1\",\"endPinId\":\"pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1\",\"rawStartPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1\",\"rawEndPinId\":\"pin-type-component_7821f33a-bdac-4457-86e4-7ce6064f4871_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"32.5000000000_1052.3166395000\\\",\\\"-27.5000000000_1052.3166395000\\\",\\\"-27.5000000000_1205.0000000000\\\",\\\"542.5000000000_1205.0000000000\\\",\\\"542.5000000000_440.0000000000\\\",\\\"-27.5000000000_440.0000000000\\\",\\\"-27.5000000000_287.3166395000\\\",\\\"32.5000000000_287.3166395000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1\",\"endPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2\",\"rawStartPinId\":\"pin-type-component_6203bc03-c8ad-4e65-acf1-0957e7d9561a_1\",\"rawEndPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"32.5000000000_1052.3166395000\\\",\\\"-27.5000000000_1052.3166395000\\\",\\\"-27.5000000000_1205.0000000000\\\",\\\"542.5000000000_1205.0000000000\\\",\\\"542.5000000000_740.0000000000\\\",\\\"616.0660345000_740.0000000000\\\",\\\"616.0660345000_674.6406500000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1\",\"endPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1\",\"rawStartPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_1\",\"rawEndPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"671.2060000000_183.8270000000\\\",\\\"671.2060000000_290.0000000000\\\",\\\"687.5017150000_290.0000000000\\\",\\\"687.5017150000_421.7864495000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0\",\"endPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0\",\"rawStartPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_0\",\"rawEndPinId\":\"pin-type-component_86163d73-1a9c-44b6-a2e1-728e256546df_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"632.5000000000_185.0000000000\\\",\\\"632.5000000000_290.0000000000\\\",\\\"617.5000000000_290.0000000000\\\",\\\"617.5000000000_425.0000000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2\",\"endPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0\",\"rawStartPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_2\",\"rawEndPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"708.7405000000_182.6540000000\\\",\\\"708.7405000000_312.5000000000\\\",\\\"812.5000000000_312.5000000000\\\",\\\"812.5000000000_425.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3\",\"endPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1\",\"rawStartPinId\":\"pin-type-component_49c909aa-82cc-42de-ad47-eeb2d04e532b_3\",\"rawEndPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"745.1020000000_182.6540000000\\\",\\\"745.1020000000_275.0000000000\\\",\\\"882.5017150000_275.0000000000\\\",\\\"882.5017150000_421.7864495000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1\",\"endPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2\",\"rawStartPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1\",\"rawEndPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1247.5000000000_515.0000000000\\\",\\\"1247.5000000000_425.0000000000\\\",\\\"970.0000000000_425.0000000000\\\",\\\"970.0000000000_732.5000000000\\\",\\\"811.0660345000_732.5000000000\\\",\\\"811.0660345000_674.6406500000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0\",\"endPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1\",\"rawStartPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_0\",\"rawEndPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1127.6169265000_320.0000000000\\\",\\\"1127.6169265000_425.0000000000\\\",\\\"1247.5000000000_425.0000000000\\\",\\\"1247.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0\",\"endPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3\",\"rawStartPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0\",\"rawEndPinId\":\"pin-type-component_af79f859-314d-4925-8469-848813fd14e6_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1052.5000000000_515.0000000000\\\",\\\"1052.5000000000_455.0000000000\\\",\\\"1000.0000000000_455.0000000000\\\",\\\"1000.0000000000_762.5000000000\\\",\\\"886.0660345000_762.5000000000\\\",\\\"886.0660345000_674.6406500000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1\",\"endPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0\",\"rawStartPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_1\",\"rawEndPinId\":\"pin-type-component_6f68e686-1c6d-45e3-a7d6-9788c0bfcfab_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1247.5000000000_320.0000000000\\\",\\\"1247.5000000000_455.0000000000\\\",\\\"1052.5000000000_455.0000000000\\\",\\\"1052.5000000000_515.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0\",\"endPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1\",\"rawStartPinId\":\"pin-type-component_6cee0eb2-6d0f-40c6-8e45-a9ca58a2c687_0\",\"rawEndPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1562.5000000000_1820.0000000000\\\",\\\"1502.5000000000_1820.0000000000\\\",\\\"1502.5000000000_1424.4905000000\\\",\\\"1564.0075000000_1424.4905000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1\",\"endPinId\":\"pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0\",\"rawStartPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1\",\"rawEndPinId\":\"pin-type-component_c80f0ed6-f74d-456d-a629-db513543e96f_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1564.0075000000_1424.4905000000\\\",\\\"1502.5000000000_1424.4905000000\\\",\\\"1502.5000000000_2180.0000000000\\\",\\\"1562.5000000000_2180.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1\",\"endPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4\",\"rawStartPinId\":\"pin-type-component_6d2add11-c610-441d-abbc-fd8eae0f97b2_1\",\"rawEndPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1564.0075000000_1424.4905000000\\\",\\\"1502.5000000000_1424.4905000000\\\",\\\"1502.5000000000_1205.0000000000\\\",\\\"1652.5000000000_1205.0000000000\\\",\\\"1652.5000000000_1075.9520000000\\\",\\\"1713.0565000000_1075.9520000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2\",\"endPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2\",\"rawStartPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2\",\"rawEndPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1359.2260000000_1291.4705000000\\\",\\\"1427.5000000000_1291.4705000000\\\",\\\"1427.5000000000_1636.4705000000\\\",\\\"1359.2260000000_1636.4705000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2\",\"endPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2\",\"rawStartPinId\":\"pin-type-component_cfdf6e28-319d-4b21-b73b-81e1fb5f7f1b_2\",\"rawEndPinId\":\"pin-type-component_fa11e16a-f0a7-42e2-a7d4-599f2d603b47_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1359.2260000000_1636.4705000000\\\",\\\"1427.5000000000_1636.4705000000\\\",\\\"1427.5000000000_1981.4705000000\\\",\\\"1359.2260000000_1981.4705000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2\",\"endPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4\",\"rawStartPinId\":\"pin-type-component_84de52eb-d97f-4432-8888-452b5250f3c1_2\",\"rawEndPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1359.2260000000_1291.4705000000\\\",\\\"1427.5000000000_1291.4705000000\\\",\\\"1427.5000000000_1205.0000000000\\\",\\\"1382.5000000000_1205.0000000000\\\",\\\"1382.5000000000_1075.9520000000\\\",\\\"1443.0565000000_1075.9520000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1\",\"endPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg\",\"rawStartPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_1\",\"rawEndPinId\":\"pin-type-power-rail_b62302e1-db31-40ba-a2dc-d3556ee2692c_1_3_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1172.5000000000_1130.0000000000\\\",\\\"1172.5000000000_1197.5000000000\\\",\\\"962.5000000000_1197.5000000000\\\",\\\"962.5000000000_875.0000000000\\\",\\\"902.5000000000_875.0000000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2\",\"endPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1\",\"rawStartPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_2\",\"rawEndPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1139.5935415000_-71.1024490000\\\",\\\"1139.5935415000_-130.0000000000\\\",\\\"1352.5000000000_-130.0000000000\\\",\\\"1352.5000000000_702.5000000000\\\",\\\"1907.5000000000_702.5000000000\\\",\\\"1907.5000000000_921.1925000000\\\",\\\"1858.0720000000_921.1925000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1\",\"endPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1\",\"rawStartPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1\",\"rawEndPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1588.0720000000_921.1925000000\\\",\\\"1555.0000000000_921.1925000000\\\",\\\"1555.0000000000_995.0000000000\\\",\\\"1907.5000000000_995.0000000000\\\",\\\"1907.5000000000_921.1925000000\\\",\\\"1858.0720000000_921.1925000000\\\"]}\"}","{\"color\":\"#f44336\",\"startPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2\",\"endPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1\",\"rawStartPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_2\",\"rawEndPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1345.0000000000_958.6010000000\\\",\\\"1382.5000000000_958.6010000000\\\",\\\"1382.5000000000_995.0000000000\\\",\\\"1555.0000000000_995.0000000000\\\",\\\"1555.0000000000_921.1925000000\\\",\\\"1588.0720000000_921.1925000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3\",\"endPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3\",\"rawStartPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3\",\"rawEndPinId\":\"pin-type-component_bcf76462-cf56-4f01-b598-ae1e6dd3ec4d_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1229.6770600000_-71.1024490000\\\",\\\"1229.6770600000_-92.5000000000\\\",\\\"1307.5000000000_-92.5000000000\\\",\\\"1307.5000000000_747.5000000000\\\",\\\"1772.5000000000_747.5000000000\\\",\\\"1772.5000000000_923.7920000000\\\",\\\"1712.3965000000_923.7920000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3\",\"endPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3\",\"rawStartPinId\":\"pin-type-component_1ac7d52d-b253-412f-8e1b-4251a9594a23_3\",\"rawEndPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1229.6770600000_-71.1024490000\\\",\\\"1229.6770600000_-92.5000000000\\\",\\\"1307.5000000000_-92.5000000000\\\",\\\"1307.5000000000_747.5000000000\\\",\\\"1517.5000000000_747.5000000000\\\",\\\"1517.5000000000_923.7920000000\\\",\\\"1442.3965000000_923.7920000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3\",\"endPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3\",\"rawStartPinId\":\"pin-type-component_390d83ab-07c8-4d04-99d0-82df7aff116b_3\",\"rawEndPinId\":\"pin-type-component_a669ed33-4ae7-4630-b33a-1a8d6006ac36_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1345.0000000000_886.2725000000\\\",\\\"1382.5000000000_886.2725000000\\\",\\\"1382.5000000000_923.7920000000\\\",\\\"1442.3965000000_923.7920000000\\\"]}\"}"],"projectDescription":""}PK
     uK\               jsons/PK
     uK\����  ��     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"ESP32 38-PIN","category":["User Defined"],"userDefined":true,"id":"69c262f4-fa86-6b73-0b2d-129f230d5ed6","subtypeDescription":"","subtypePic":"ab296a80-256f-428c-a4e8-e177cdc61bff.png","iconPic":"c19b89aa-68d9-4a98-b509-123aa1ab0169.png","imageLocation":"local_cache","componentVersion":3,"pinInfo":{"numDisplayCols":"10.11813","numDisplayRows":"20.61563","pins":[{"uniquePinIdString":"0","positionMil":"71.30768,2021.52677","isAnchorPin":true,"label":"3.3 V"},{"uniquePinIdString":"1","positionMil":"71.30768,1921.52677","isAnchorPin":false,"label":"RESTART/EN"},{"uniquePinIdString":"2","positionMil":"71.30768,1821.52677","isAnchorPin":false,"label":"GPIO 36"},{"uniquePinIdString":"3","positionMil":"71.30768,1721.52677","isAnchorPin":false,"label":"GPIO 39"},{"uniquePinIdString":"4","positionMil":"71.30768,1621.52677","isAnchorPin":false,"label":"GPIO 34"},{"uniquePinIdString":"5","positionMil":"71.30768,1521.52677","isAnchorPin":false,"label":"GPIO 35"},{"uniquePinIdString":"6","positionMil":"71.30768,1421.52677","isAnchorPin":false,"label":"GPIO 32"},{"uniquePinIdString":"7","positionMil":"71.30768,1321.52677","isAnchorPin":false,"label":"GPIO 33"},{"uniquePinIdString":"8","positionMil":"71.30768,1221.52677","isAnchorPin":false,"label":"GPIO 25"},{"uniquePinIdString":"9","positionMil":"71.30768,1121.52677","isAnchorPin":false,"label":"GPIO 26"},{"uniquePinIdString":"10","positionMil":"71.30768,1021.52677","isAnchorPin":false,"label":"GPIO 27"},{"uniquePinIdString":"11","positionMil":"71.30768,921.52677","isAnchorPin":false,"label":"GPIO 14 (HSPI CLK)"},{"uniquePinIdString":"12","positionMil":"71.30768,821.52677","isAnchorPin":false,"label":"GPIO 12 (HSPI MISO)"},{"uniquePinIdString":"13","positionMil":"71.30768,721.52677","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"14","positionMil":"71.30768,621.52677","isAnchorPin":false,"label":"GPIO 13 (HSPI MOSI)"},{"uniquePinIdString":"15","positionMil":"71.30768,521.52677","isAnchorPin":false,"label":"GPIO 9"},{"uniquePinIdString":"16","positionMil":"71.30768,421.52677","isAnchorPin":false,"label":"GPIO 10"},{"uniquePinIdString":"17","positionMil":"71.30768,321.52677","isAnchorPin":false,"label":"GPIO 11"},{"uniquePinIdString":"18","positionMil":"71.30768,221.52677","isAnchorPin":false,"label":"5 V"},{"uniquePinIdString":"19","positionMil":"971.30768,221.52677","isAnchorPin":false,"label":"GPIO 6"},{"uniquePinIdString":"20","positionMil":"971.30768,321.52677","isAnchorPin":false,"label":"GPIO 7"},{"uniquePinIdString":"21","positionMil":"971.30768,421.52677","isAnchorPin":false,"label":"GPIO 8"},{"uniquePinIdString":"22","positionMil":"971.30768,521.52677","isAnchorPin":false,"label":"GPIO 15 (HSPI CS)"},{"uniquePinIdString":"23","positionMil":"971.30768,621.52677","isAnchorPin":false,"label":"GPIO 2"},{"uniquePinIdString":"24","positionMil":"971.30768,721.52677","isAnchorPin":false,"label":"GPIO 0"},{"uniquePinIdString":"25","positionMil":"971.30768,821.52677","isAnchorPin":false,"label":"GPIO 4"},{"uniquePinIdString":"26","positionMil":"971.30768,921.52677","isAnchorPin":false,"label":"GPIO 16 (RX2)"},{"uniquePinIdString":"27","positionMil":"971.30768,1021.52677","isAnchorPin":false,"label":"GPIO 17 (TX2)"},{"uniquePinIdString":"28","positionMil":"971.30768,1121.52677","isAnchorPin":false,"label":"GPIO 5 (VSPI CS)"},{"uniquePinIdString":"29","positionMil":"971.30768,1221.52677","isAnchorPin":false,"label":"GPIO 18 (VSPI CLK)"},{"uniquePinIdString":"30","positionMil":"971.30768,1321.52677","isAnchorPin":false,"label":"GPIO 19 (VSPI MISO)"},{"uniquePinIdString":"31","positionMil":"971.30768,1421.52677","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"32","positionMil":"971.30768,1521.52677","isAnchorPin":false,"label":"GPIO 21 (I2C SDA)"},{"uniquePinIdString":"33","positionMil":"971.30768,1621.52677","isAnchorPin":false,"label":"GPIO 3 (RX0)"},{"uniquePinIdString":"34","positionMil":"971.30768,1721.52677","isAnchorPin":false,"label":"GPIO 1 (TX0)"},{"uniquePinIdString":"35","positionMil":"971.30768,1821.52677","isAnchorPin":false,"label":"GPIO 22 (I2C SCL)"},{"uniquePinIdString":"36","positionMil":"971.30768,1921.52677","isAnchorPin":false,"label":"GPIO 23 (VSPI MOSI)"},{"uniquePinIdString":"37","positionMil":"971.30768,2021.52677","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":true,"componentImageSvgUrl":"https://abacasstorageaccnt.blob.core.windows.net/cirkit/4546d829-0f3e-4357-ac32-46d75e79207c.svg","propertiesV2":[]},{"subtypeName":"Load cell 50kg","category":["User Defined"],"id":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f6e2a5fb-4294-42a3-957b-9521668fdddb.png","iconPic":"8fef4bdb-224a-4a07-91a3-222e74c30575.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"10.56604","pins":[{"uniquePinIdString":"0","positionMil":"442.88333,1046.19855","isAnchorPin":true,"label":"black wire"},{"uniquePinIdString":"1","positionMil":"519.04333,1036.67855","isAnchorPin":false,"label":"red wire"},{"uniquePinIdString":"2","positionMil":"599.96333,1031.91855","isAnchorPin":false,"label":"white wire"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Load cell 50kg","category":["User Defined"],"id":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f6e2a5fb-4294-42a3-957b-9521668fdddb.png","iconPic":"8fef4bdb-224a-4a07-91a3-222e74c30575.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"10.56604","pins":[{"uniquePinIdString":"0","positionMil":"442.88333,1046.19855","isAnchorPin":true,"label":"black wire"},{"uniquePinIdString":"1","positionMil":"519.04333,1036.67855","isAnchorPin":false,"label":"red wire"},{"uniquePinIdString":"2","positionMil":"599.96333,1031.91855","isAnchorPin":false,"label":"white wire"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Load cell 50kg","category":["User Defined"],"id":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f6e2a5fb-4294-42a3-957b-9521668fdddb.png","iconPic":"8fef4bdb-224a-4a07-91a3-222e74c30575.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"10.56604","pins":[{"uniquePinIdString":"0","positionMil":"442.88333,1046.19855","isAnchorPin":true,"label":"black wire"},{"uniquePinIdString":"1","positionMil":"519.04333,1036.67855","isAnchorPin":false,"label":"red wire"},{"uniquePinIdString":"2","positionMil":"599.96333,1031.91855","isAnchorPin":false,"label":"white wire"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"SSR - 40da","category":["User Defined"],"id":"b97d5804-295d-4a63-b66d-23cafcd44586","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"2b856d38-88e4-4759-8ee8-6b01c1d6fb9d.png","iconPic":"9aa3d03b-0c22-4f62-98c6-f5f844a0dc7c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.33938","numDisplayRows":"25.44036","pins":[{"uniquePinIdString":"0","positionMil":"376.63233,286.56467","isAnchorPin":true,"label":"IN-"},{"uniquePinIdString":"1","positionMil":"1537.26233,294.40467","isAnchorPin":false,"label":"IN+"},{"uniquePinIdString":"2","positionMil":"353.10233,2231.40467","isAnchorPin":false,"label":"OUT"},{"uniquePinIdString":"3","positionMil":"1537.26233,2231.40467","isAnchorPin":false,"label":"OUT"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"SSR - 40da","category":["User Defined"],"id":"b97d5804-295d-4a63-b66d-23cafcd44586","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"2b856d38-88e4-4759-8ee8-6b01c1d6fb9d.png","iconPic":"9aa3d03b-0c22-4f62-98c6-f5f844a0dc7c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.33938","numDisplayRows":"25.44036","pins":[{"uniquePinIdString":"0","positionMil":"376.63233,286.56467","isAnchorPin":true,"label":"IN-"},{"uniquePinIdString":"1","positionMil":"1537.26233,294.40467","isAnchorPin":false,"label":"IN+"},{"uniquePinIdString":"2","positionMil":"353.10233,2231.40467","isAnchorPin":false,"label":"OUT"},{"uniquePinIdString":"3","positionMil":"1537.26233,2231.40467","isAnchorPin":false,"label":"OUT"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"SSR - 40da","category":["User Defined"],"id":"b97d5804-295d-4a63-b66d-23cafcd44586","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"2b856d38-88e4-4759-8ee8-6b01c1d6fb9d.png","iconPic":"9aa3d03b-0c22-4f62-98c6-f5f844a0dc7c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"19.33938","numDisplayRows":"25.44036","pins":[{"uniquePinIdString":"0","positionMil":"376.63233,286.56467","isAnchorPin":true,"label":"IN-"},{"uniquePinIdString":"1","positionMil":"1537.26233,294.40467","isAnchorPin":false,"label":"IN+"},{"uniquePinIdString":"2","positionMil":"353.10233,2231.40467","isAnchorPin":false,"label":"OUT"},{"uniquePinIdString":"3","positionMil":"1537.26233,2231.40467","isAnchorPin":false,"label":"OUT"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"SHT31","category":["User Defined"],"id":"01534432-bd5d-4550-957a-0d4278d98851","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"245bc533-66be-4bb3-b22a-43c007a581bd.png","iconPic":"51c64262-e188-46ba-9658-f0d60e053320.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.10530","numDisplayRows":"12.00840","pins":[{"uniquePinIdString":"0","positionMil":"148.22254,110.39582","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"354.40178,102.00070","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"785.40746,118.79095","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"2","positionMil":"587.62333,102.00070","isAnchorPin":false,"label":"SCL"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"HX711","category":["User Defined"],"id":"8f8ecf0b-b7ef-4a48-962c-7614bb5a7d82","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"7fb2f62e-2fb5-47b1-9980-8ec272392bae.png","iconPic":"2db9ecad-5c51-4c64-ac4d-4ae785eb4e5c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"16.48980","pins":[{"uniquePinIdString":"0","positionMil":"336.36333,1410.79646","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"462.48333,1409.27646","isAnchorPin":false,"label":"DT"},{"uniquePinIdString":"2","positionMil":"582.97333,1413.77646","isAnchorPin":false,"label":"SCK"},{"uniquePinIdString":"3","positionMil":"698.96333,1409.27646","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"4","positionMil":"217.16333,205.70646","isAnchorPin":false,"label":"E+"},{"uniquePinIdString":"5","positionMil":"340.28333,206.92646","isAnchorPin":false,"label":"E-"},{"uniquePinIdString":"6","positionMil":"462.94333,205.70646","isAnchorPin":false,"label":"A-"},{"uniquePinIdString":"7","positionMil":"585.15333,204.79646","isAnchorPin":false,"label":"A+"},{"uniquePinIdString":"8","positionMil":"703.72333,205.73646","isAnchorPin":false,"label":"B-"},{"uniquePinIdString":"9","positionMil":"829.55333,205.73646","isAnchorPin":false,"label":"B+"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Heating Coil","category":["User Defined"],"id":"1255ec18-62c0-4252-8215-c2ff45234b02","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cb669bd1-12cf-42eb-9243-39a8a80a0435.png","iconPic":"1be29400-b52e-43b8-b531-83e2df2121b6.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"17.53053","numDisplayRows":"25.27840","pins":[{"uniquePinIdString":"0","positionMil":"591.67763,36.10772","isAnchorPin":true,"label":"Vcc"},{"uniquePinIdString":"1","positionMil":"1354.94763,46.15772","isAnchorPin":false,"label":"Gnd"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Fan","category":["Output"],"userDefined":true,"id":"6635379e-9371-f184-7e48-a00d3644b40e","subtypeDescription":"","subtypePic":"146a6d58-0553-42c9-b8c7-03425202d69a.png","iconPic":"d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"19.68504","pins":[{"uniquePinIdString":"0","positionMil":"175.51732,233.57781","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"175.86674,322.02337","isAnchorPin":false,"label":"5V"}],"pinType":"wired"},"properties":[],"componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Load cell 50kg","category":["User Defined"],"id":"2c3f3b4a-c088-4e0e-9d5c-77a3eddf6ffe","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"f6e2a5fb-4294-42a3-957b-9521668fdddb.png","iconPic":"8fef4bdb-224a-4a07-91a3-222e74c30575.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"10.00000","numDisplayRows":"10.56604","pins":[{"uniquePinIdString":"0","positionMil":"442.88333,1046.19855","isAnchorPin":true,"label":"black wire"},{"uniquePinIdString":"1","positionMil":"519.04333,1036.67855","isAnchorPin":false,"label":"red wire"},{"uniquePinIdString":"2","positionMil":"599.96333,1031.91855","isAnchorPin":false,"label":"white wire"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Electrolytic Capacitor","subtypeDescription":"","subtypePic":"48caf11c-09fe-45e4-9b76-5b0bfa123a56.png","id":"14d7a2a7-6581-4d0a-a495-63cc6355f7b9","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"48.90000,0.00000","endPositionMil":"48.90000,-140.00000","isAnchorPin":true,"label":"-"},{"uniquePinIdString":"1","startPositionMil":"148.90000,0.00000","endPositionMil":"148.90000,-140.00000","isAnchorPin":false,"label":"+"}],"numDisplayCols":"1.96860","numDisplayRows":"4.82660","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"16bd2965-d7b7-4d97-b402-ac1747e7568c.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"buzzer","category":["User Defined"],"id":"02adc9af-9099-49f0-8d17-97b22a4179bc","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae99f124-1aaf-4a6e-8177-44087bd956ce.png","iconPic":"f7e3f572-2cc7-414e-8b58-58f37a09912a.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"4.72400","numDisplayRows":"4.72400","pins":[{"uniquePinIdString":"0","positionMil":"236.27629,383.36636","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"236.27629,83.36636","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"plugable terminal ds18820","category":["User Defined"],"id":"84de3699-1b7e-4fcb-b51f-13b7bf5839ea","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"98bdfb38-4044-46ed-976e-d2b53bff2879.png","iconPic":"1a257b89-3953-41e9-990a-6c271080df8c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"6.02496","pins":[{"uniquePinIdString":"0","positionMil":"621.83667,221.71444","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"619.55667,301.51444","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"619.55667,388.15444","isAnchorPin":false,"label":"DAT"},{"uniquePinIdString":"3","positionMil":"195.45667,406.39444","isAnchorPin":false,"label":"DAT"},{"uniquePinIdString":"4","positionMil":"197.73667,306.07444","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"5","positionMil":"200.01667,203.47444","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"ADAPTO 5 VOLT","category":["User Defined"],"id":"c16bfa02-5154-4f39-9ff1-d473663907f3","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"d6a4f4f6-fe0f-43ac-893b-20774d3ea628.png","iconPic":"c7b8e0ca-67ed-4237-9266-7527aa3ce92a.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"21.00000","numDisplayRows":"20.00000","pins":[{"uniquePinIdString":"0","positionMil":"0.00000,1250.00000","isAnchorPin":true,"label":"+"},{"uniquePinIdString":"1","positionMil":"0.00000,1150.00000","isAnchorPin":false,"label":"-"},{"uniquePinIdString":"2","positionMil":"1142.66000,0.00000","isAnchorPin":false,"label":"110V AC"},{"uniquePinIdString":"3","positionMil":"1624.85000,0.00000","isAnchorPin":false,"label":"110V Neutral"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Outlet","category":["User Defined"],"id":"ef0da927-5348-4d94-b21a-42d8a46ff031","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"fe816bc3-a1ac-4496-aca2-7e46c72bb630.png","iconPic":"559c8cb2-c573-4147-bde4-a0b817dc20ed.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"14.17323","numDisplayRows":"24.01575","pins":[{"uniquePinIdString":"0","positionMil":"231.09252,370.66142","isAnchorPin":true,"label":"Ground"},{"uniquePinIdString":"1","positionMil":"1201.57252,1762.71142","isAnchorPin":false,"label":"Hot 1"},{"uniquePinIdString":"2","positionMil":"1201.57252,739.53142","isAnchorPin":false,"label":"Hot 2"},{"uniquePinIdString":"3","positionMil":"230.40252,1745.38142","isAnchorPin":false,"label":"Neutral 1"},{"uniquePinIdString":"4","positionMil":"234.80252,730.98142","isAnchorPin":false,"label":"Neutral 2"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Solar Panel","category":["User Defined"],"id":"aec5eff0-da06-45e7-8932-95bc26fc4e6a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a0bdb5a7-9945-4126-87cb-dac9f24142ab.png","iconPic":"68998569-73de-4f26-b1b3-0b6c45f8499f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"25.99688","numDisplayRows":"42.32704","pins":[{"uniquePinIdString":"0","positionMil":"37.50972,599.77850","isAnchorPin":true,"label":"gnd"},{"uniquePinIdString":"1","positionMil":"37.50972,717.66757","isAnchorPin":false,"label":"vcc"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"12V 200Ah Battery","category":["User Defined"],"id":"8903b643-ed64-43f6-b56c-46542b1c2184","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"a003a845-706b-4c0a-bac4-0f60a60b44e4.png","iconPic":"8a348e4e-00a9-420c-8c54-2da977db0968.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"18.12093","numDisplayRows":"18.12093","pins":[{"uniquePinIdString":"0","positionMil":"273.68421,1503.32033","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"1573.68421,1503.32033","isAnchorPin":false,"label":"12V"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"AC Circuit Breaker","category":["User Defined"],"id":"023546b5-ca70-49d6-8fe2-6f4e8641da15","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"9d915518-60ad-41a3-8ee2-5a1cc2d88e80.png","iconPic":"a652ce68-b987-46e6-8408-d5645582d4d7.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"28.40524","numDisplayRows":"28.40524","pins":[{"uniquePinIdString":"0","positionMil":"1181.47506,2240.89049","isAnchorPin":true,"label":"Live"},{"uniquePinIdString":"1","positionMil":"1648.15316,2262.31416","isAnchorPin":false,"label":"Neutral"},{"uniquePinIdString":"2","positionMil":"1171.91529,576.61949","isAnchorPin":false,"label":"Live OUT"},{"uniquePinIdString":"3","positionMil":"1671.91529,576.61949","isAnchorPin":false,"label":"Neutral OUT"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Solar Panel","category":["User Defined"],"id":"aec5eff0-da06-45e7-8932-95bc26fc4e6a","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a0bdb5a7-9945-4126-87cb-dac9f24142ab.png","iconPic":"68998569-73de-4f26-b1b3-0b6c45f8499f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"25.99688","numDisplayRows":"42.32704","pins":[{"uniquePinIdString":"0","positionMil":"37.50972,599.77850","isAnchorPin":true,"label":"gnd"},{"uniquePinIdString":"1","positionMil":"37.50972,717.66757","isAnchorPin":false,"label":"vcc"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"12V/24V ออโต้ 20A MPPT","category":["User Defined"],"id":"28def945-d566-45d1-91c0-cb2676c61db2","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"a27a8979-5023-407e-b6b7-e8628572ca80.png","iconPic":"5441ee9b-7343-4a92-92bb-e3ea11bfaf7c.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"47.00000","numDisplayRows":"47.00000","pins":[{"uniquePinIdString":"0","positionMil":"1731.38000,553.42000","isAnchorPin":true,"label":"+ SL"},{"uniquePinIdString":"1","positionMil":"1989.42000,561.24000","isAnchorPin":false,"label":"- SL"},{"uniquePinIdString":"2","positionMil":"2239.65000,569.06000","isAnchorPin":false,"label":"+ B"},{"uniquePinIdString":"3","positionMil":"2482.06000,569.06000","isAnchorPin":false,"label":"- B"},{"uniquePinIdString":"4","positionMil":"2732.29000,561.24000","isAnchorPin":false,"label":"+ L"},{"uniquePinIdString":"5","positionMil":"2966.88000,561.24000","isAnchorPin":false,"label":"- L"}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Power Inverter","category":["User Defined"],"id":"b8a657e4-3f8b-4e3e-a2bd-792a2961387f","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"10aa979f-dd42-43c7-9c2f-b8fbfcd42f21.png","iconPic":"687e948c-dc0a-4fdc-b588-e952ae529de1.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"27.72857","numDisplayRows":"13.86428","pins":[{"uniquePinIdString":"1","positionMil":"103.40279,284.15330","isAnchorPin":true,"label":"-"},{"uniquePinIdString":"0","positionMil":"103.40279,1083.37379","isAnchorPin":false,"label":"+"},{"uniquePinIdString":"2","positionMil":"2710.75245,1003.52969","isAnchorPin":false,"label":"+"},{"uniquePinIdString":"3","positionMil":"2710.75245,402.97290","isAnchorPin":false,"label":"-"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"AC Circuit Breaker","category":["User Defined"],"id":"023546b5-ca70-49d6-8fe2-6f4e8641da15","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"9d915518-60ad-41a3-8ee2-5a1cc2d88e80.png","iconPic":"a652ce68-b987-46e6-8408-d5645582d4d7.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"28.40524","numDisplayRows":"28.40524","pins":[{"uniquePinIdString":"0","positionMil":"1181.47506,2240.89049","isAnchorPin":true,"label":"Live"},{"uniquePinIdString":"1","positionMil":"1648.15316,2262.31416","isAnchorPin":false,"label":"Neutral"},{"uniquePinIdString":"2","positionMil":"1171.91529,576.61949","isAnchorPin":false,"label":"Live OUT"},{"uniquePinIdString":"3","positionMil":"1671.91529,576.61949","isAnchorPin":false,"label":"Neutral OUT"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Outlet","category":["User Defined"],"id":"ef0da927-5348-4d94-b21a-42d8a46ff031","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"fe816bc3-a1ac-4496-aca2-7e46c72bb630.png","iconPic":"559c8cb2-c573-4147-bde4-a0b817dc20ed.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"14.17323","numDisplayRows":"24.01575","pins":[{"uniquePinIdString":"0","positionMil":"231.09252,370.66142","isAnchorPin":true,"label":"Ground"},{"uniquePinIdString":"1","positionMil":"1201.57252,1762.71142","isAnchorPin":false,"label":"Hot 1"},{"uniquePinIdString":"2","positionMil":"1201.57252,739.53142","isAnchorPin":false,"label":"Hot 2"},{"uniquePinIdString":"3","positionMil":"230.40252,1745.38142","isAnchorPin":false,"label":"Neutral 1"},{"uniquePinIdString":"4","positionMil":"234.80252,730.98142","isAnchorPin":false,"label":"Neutral 2"}],"pinType":"wired"},"properties":[],"propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Fan","category":["Output"],"userDefined":true,"id":"6635379e-9371-f184-7e48-a00d3644b40e","subtypeDescription":"","subtypePic":"146a6d58-0553-42c9-b8c7-03425202d69a.png","iconPic":"d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"19.68504","pins":[{"uniquePinIdString":"0","positionMil":"175.51732,233.57781","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"175.86674,322.02337","isAnchorPin":false,"label":"5V"}],"pinType":"wired"},"properties":[],"componentVersion":1,"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Comment V2","category":["User Defined"],"componentClass":"textbox","userDefined":true,"id":"9a5a4baa-44d4-4aa0-8d82-488487322b20","subtypeDescription":"","subtypePic":"c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"text box (click to edit)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundColor","label":"Background Color","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"backgroundOpacity","label":"Background Opacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"textColor","label":"Text Color","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"fontSize","label":"Font Size","description":"","units":"","type":"integer","value":"10","displayFormat":"input","showOnComp":false,"isVisibleToUser":true},{"version":2,"id":"font","label":"Font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true}],"iconPic":"d3694a2e-5bba-40c3-8069-8db85c4c9209.png","componentVersion":1,"imageLocation":"local_cache","propertiesV2":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     uK\               images/PK
     uK\���)G )G /   images/ab296a80-256f-428c-a4e8-e177cdc61bff.png�PNG

   IHDR  _  �   �D��   	pHYs  \F  \F�CA  ��IDATx��	�$�}�����an� Y��[Bօ-�r ��!��Z��!mlh-i�v�c{��l��]�$^�	$4���p_b�a���{�>���>)?���Y��U���������ʬ������jj�>�������555�_��Y+++��~����fDE�?���s�]`�B9�3v���M�U@I�,�~L�4��ҿ_)�|������~���k��U��o��ҏO���������7��E<J�!�.R���5��0=�����������������`w��O%�>���}yy�%����h6B!�NI�\T�qQss��~�7~����x�]w�H�9����Ҏ���}�I�-!�B�B���tc���K|gyy�3?���}l�URx7�>��.��dLKK�ikk3�����.��W�?~X�������	!�B$]a��Go ���υ��raAآ~��[�[�I���;���컢���:J����_�4v�Ż��Lgg���0 �����@	!�B��������F{{{��t?sss��@��� ����y���]���;���B��+�rJ�����J�{MF0===� ������m���fjj�!�B@tuww�5kּe�J"�Ɔ�gzz���̜$�J��TI��}�M7}�$�"3C#�«�!���y�� \�}}}���V ��P�rI
!��DF�4�+�_��cǎy�?%���sssw�t�o�u�]3a�*����/4�ر�e&��Ɂg��D�"�̄B!�X] �R{��|��Аg�������}���n��w��b�B�WIx��ҏeq��Q�Y����B!V.�)k0(����<ndB�������o���$�n���������*����d�X�`B!�hl^X�򬈅�6������ϕtՏ������<A|}��-	���E�TDP��˂�s�,`B!D�B^�z�"e߈>�uA��J���M7�t�? ��URk�/�pS��,��	����8!�B«V��i���sll�\�������~���-������^�Z��ի�pRp{>|8�>�B!
Z#I�Ь��F'*/��o7�p�W�瞽�筣,��?-���A0�T(��}�{_��y衇���rxG����B!Dc@�W�Ц��_�K�aP;v�0o��f���>T[�{:K��.��_��'�n����B��L�����+���oL���o��<�쳱�.�Ob�TL!�h-��{��322�j?��o�f�ﾊ���4����-7�p��q�=�Lx����>Z�e�#�I�8/�s۷oO��;���{��[n�`�kP��~B!�Ɨ4������������}n��f��h9���Y�����>\��5k.�ScP}I���$��_N��4�%��B�� ��W^I��$�ۭ
�~����z�M7��>�]��$iX�7�~�E�	!���ԲMa��--+++�������uff�%uV��J�z�8��B!�.�<�ا%������J����$���b�.�{�˗B!���Z�#�0"um����yY�]׏O!��)�\"�����bg��{Y�YW!���ր�c<�>��9ESN�B!�)�\4���y�'��Q���AQ�U!����]`�1�"�2�x��q9A�K!�(6ij}�M�Kb�����)���Ǐ;-�8>!�B�"�/tWfi��r�֗j|	!�����CO��-3�5??�5�t�O!��a� s�vg�����Š�Xҁc+��R!��}���+�df�������֯��.��w�;�~����&~O�ɥB!

���/��~�W5�{v�����B��ii���i�����Uj�>;y�פ�m��!
�BQ|�d1��Y�&�{�[�nM��$��SSS��T|���yooo��|�K_2_�����ѣG���p��MLL�.�B!����������/��/���߿�lٲ%��7���̛"�)g�z����ڵk�>/�M.G!������q�����kw��m����ʔ,'�0�;v���s�H966�Y�������͇>��L�[��B!D1���[�����k����ev����].⋠3���ࠩ�P�2�B��e||�3��+�����E|������+��2�B�0���	yՂ�B��!�#��p�aˣ�6���B!V��G��F^�v�vs�|e��e�;��,K� �A����B���^/�]���P-hDW�d���6::���k-���E����B����c(�Jr_-Ag�7�ē�E|������E�"�/� �y��%�B ����Q�+}A;zCRZ�&�,��al6E��(ǀυ�r���B!�z�`���Ok�9�d�A�`=�z����/?|9���`��η�jK�,\B!�H��}�jtڂ��,bǝ_~��l�h	!�"+cy�uV|	!�B4"_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9"�%�B�#_B!�9��jmm5��ͦ��Ŭ��x����Ғ9~��B!��t������5���%N����v�����d ���"_�`,..���3;;+1&�B�� ����<���]a`�Ak��ϛ��������/�����Y�����E|MMM�l`�B�8����=#O�&�6���̌�Uc����Z�f����:〥l``�S��B!��}���g:::��,?8���i��{2�1�:��D(�B�����A�<8>>�jP�BQ|0� �ʅ1��5�رc�>��/�֮r�p׮]k�=�ņ	!�bu���ȓ�Ř��+^���*�2/���aO�,'�B�Ɔ�hhȴ���O�`��[r_X��^�/'AL!�hl윟��؀|ܐ��E|�V�e�����Q/ _!��s}=���3� qC�#s�e�O�nI�A�0!�B4i�HdU𴕋7�\|1�T�i��V�~8P1��`̂eB!Dc@�5?�q�F�#WG��j}�������{M��/�U�5����S��g������o<X��(RbB!�$5C����،����ϫ��jv��mv��i^z���at*g��T|���;�H��ݛx������w�mn��X�M[�6J�
!��8�vAIٵkW������������7�\�h+������ �~��%��T�"�%�B4��i�������h��I�SX����;Lҫ1O�)�Q!�(6i�^yA@��=�����K!�(.��YZ�QZ(3���`���'�B��>��z�%L��L|U�ƙ5��B!�S���c���쨳n�]-��B!�S��q �<7����H|	!�Ŧsy�r�^����F!�ť���Ff⋝��HWT�^!�(4E��Î13�E-����BQ\�P�3Lod&�(*�r
�ėBQl��쮁0W�#�RS�z��-�B!�C
�/W;�Di���;���b�#'�u�,�B�ʠ7���Γ���knn.V�%�����o�9�x?�����e\!�łV�I�M�>�x_I�cuP�������%����~������B!Dc��P�����������Tƛ$�5��13_����Qp`۷o7��ǫ����d=0EȎB!D<&''���p��>��C�C��'�҂���� �~jj*��Y����zG�~!��������GP1� !�B4)B��x����C5*i�F�b/������7�WT\U!�h8����H�}��\��FQ��,=�
Uy	!��1��r��Q322R�J���K�[oG܏T��c�5���
!��� ~`CCC�0<}�;N��\k[�_��8�xIx	!���A�����9$�pll,vB_����r�}}}��R�'����!�B��F�PX֭	�Bo$�)�]|�hL��qAp��TI	!�bu���ͩ�Pk���w-M����/�/ˠP�����&�A�@TS�C!���(B�0��5�;�V��^动V�n��B"�A� k�4Q�'��A'�B�ǆ"a�Ag�7�q�"��֨E8S�ŗ�806܅�/ܑT�'X�n�����ZB!D�X��^0���V�!��lv������c�YB!�Y��"L��JN�/!�B�FE�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G$��B!rD�K!�"G
#������ʊB!���d�7�_�������fZ[[MKK�[���Ғ9~��Y\\4����O!�B�8�-:::<�a�Fss�	�AkX���`��(sB|񥻻�MWW�I_>B��b���4��������x���B!���~@7�Y��]�@���Zރ�B��5�Yu_|���>o0��D��������B!�'�0�*x*}z�k���DjV7񅥋��k��(�cǎ���Y#�B��	!L�����yCCCfnn��I>��/T���`,�_Zt6�t||\��B!�*c޵,Ag�g������B���*�p�k�@�`P����ѣG�B!V	x�zzzr�F%�KXr_/��y���'&�B4>y
/?x��
�\�n@*o�e�>_E.H!��1��X�eA댎�VtA�"����=TO���I!R!���WY�x�cϑ#G�z�2_�]����aeB!=.`�_�E��(.ɿ����z?��z�y��7+�U�IP!������|���g�X�j��7�iv���wJ^Q�5�ؓ����Ui0Dv��c}�c3w�}����?���%qAV[�V!�n�$��Yi��>��ϛ����3��ۿ]Q�pLĚ����B�ƅJ���ַ�����7�q��H%��B���5a��~{�����^'�V_�]��A2_T���`@j�|B!��+q�apla�~��/\{.���-�&�B����eǜjAk�*�\�*'�%�B��Z���%QZ(3�U���qq�%*�B�x�ծ�8��Ǐ���,w�2��C!�B��s9ǘ��r���B!�S��<��6O	!�B4��/�8��H�WB!�;a.+k����S����=k����$��B�he���ZE_�Y%�L�>�}�٩��
!�(&/��Rh=�F'�w�+`��U|-,,x��]E텄B�b��r9��_���L�����0�C!�B�)�{���g��IR�>/��`���BQ|fggS��<�sr_@ `�5::j6nܘj��eqคBQ|8|�\]�n�K��$�����T|�Fɼ+x��غukU�B�Ʊfa���Q!�hH6�����#G�x�crr2��h�瘢�<�رcfxx8���/����믯j?q݈��B!�cϚ5kb�m����s��gz<x��ebf.��2qJ�A����*�B�d`��ƞzg>�j���(��\
qq����܍�z	!��	����@ݎ��RU���"����H�Qx�����B!D�������޺���Ö�"C��ѣfhh(W� 0���(�B4<��z$�//02a�[�=W3~P�0	�Q�	R5�NfӦM��+�4��v����2B!�#%��z�)��Ϛ���1)�Q��Ȭc�8q-^��}��I >��\����f�⬳ΪY'����&�UNyS������W_m�B��|�#f߾}�����?~��.���̋�R�3�b�����p�`D|�dA��G#O�:_�i[��������<܌�{�����_��_��=����?�yg�>	!�(���7��M�o}�������9��Ӎkl۶�<���u�?s!7tq`I
��QG2aں�u_�@�G�yK��f`\�\^���`��B�������gq���*ۆ���*��Z�Q����*�,��`l���O��ߔ����.�<[�C.3�w�l��F���9�����?��?9Ixq!�ڵ�l^!������SO5k׮=����<�����Ñ��|�^�v ����瘙�ƎF<��+`lVo�;+�ZVk��F�bȝ_~0�jm����{�ns�}�i��� �u���k���-��p���?l��կ�9V���ė�����='d�\w�u'�#~�F�
!D#��/xq�]t�[�{���m^}�U388hDq��j@����s�	���%����Pj�/�Ȓg�]m���/Y\j33skLG��ii�>� �bK�!����"��:��F|_j5�fi)�R�?��r���^o3f����6�����})�*�'�Ņg�_|����d�4��F��|cٻ�ė�4�əo�0|�l9h�B�j a�}����{u*W_a��zӻf�����	!����Jx�����X�K!D5�NQ_$�
��bm�H
!�X�,,f��P�G�@��)�X!Du��-�����8��*�B!���d��F�����a����VF!�ձn𰙚�6�S�F��/���*	��%�5a�B�j�,ؙ�v�G���fv�ӈ|��r
�n9`:��MK�
�
!��5+f����-�e��������#�� m-���s�!�Y��z��ZZ��Y4"$��B!rD�K!�"G$��B!rD��A�N��X�]^i6B!D��z���X�]^�$������4�%�B!�dy��鮡�
^{�5���S��ZYY1���:�sL{��B
!D#��/����g����n�ښL6=��,aH|U��w�Y��:~��ٹs�ɂ��������!�h<������۷g��Kj���e�����lii1��ͦ���,//{���%O�,..z?�B!����Z���~�6����7����[����tvv��������ϛ��op�B!�@_�Y����$�5������l�B��� n*� X��1�l�ө�)o��B! ���#OZ:::�������H+��&�0��]a`=��ױc�<��B!V'�1�,��k�3>����'ĒR�� �k5AP�###^� ���زeK��#B1iI\��(��˹瞛K��M�<���#G����1S�S3�[a�������C�X�c39����_\kY˪��o��oz�p�"�B�t|��\`.�m�6����_�	�����)"3��U|�%��`e���B!�K�<��������4��� �0��2��}�l9���3c��F!��~��g|ص��[�0EoW���BP�`�\���/��ņ��~�r�&�1��EȄlmY2k:�𵶨��B�p��c�'���c�\�p�8�kݺu�P�\���b�	+U��\|�����D3X_��S>m��?��́ʾ�"-IP�B!܇9>����g>�%����_7o���y����/��ܞxܦ��#?'s���c�#Hm߾}�?�������w�mn�喊�ᤐ��/!��q@����={�$��_��_�[o���|���>�@kPm!�ؓ����w0��q�=�$�GR7�U�.� [Qz!�9���dj�='w;II�9���c����2�d*�l��kp\.[��N��~�پ`�{��uG<��BQ+f�:���fb��,,�$��Y�"�aU�3_���&�� �2j@ܡ��:�;��ts��-�����cF!������̾#�sM�IZ�5/�B�{�L|�B���!	EiĽ��� w��b�:�B���Ɂ��ʀ+�j���r_��\��+�����f�����F!�H����2�\C
W��B����z)ՊZ6�΋�y��B��[p�R�׵J�$�U+��-�V(�*�BTs��r���0�0��*�\6���h��Q��B���hף�Z�m�T����0����!�Ql>`&�{��|�ݏE4�@f�2.JQZ�47�6�K�W�B�jhi^2�n~ռyx��*͇��Օ(�\�k�/��.�}�|�h�:�?f:��LO�LIĺ{�B!����Mk����n3��a]k�+m� e���Ff�^�.�/��U�J�k��#�Bd	"��{ncF''�\��-aǘ�:���˅ϊT�K!�'��\�����H�����د�J�y����I�f��!�B!��,M��4�#i�(���勸����L7�pC���v�m��c�M!�ņ�=i�W�q��&z��\xK�L�������������|��_N��g�y��933c���c�gzzڸ��L�ye^K�m!�"�Cc#f|j �k�:��5�ŭ��裏z������x�׼�f�ڵe_��gaa!�o�����)ϢU��������y�������d,��+̀�	�EzB���[0��$���������(����(�L��
+S��/O~�c�j_q�V+���c���/|z���'�S!�(0G���!�������]@���hUe**%b��r9B� _d9,�¾�����ZZ�����"p�u�yH!���=��c�{�9�����q���?��+�DU�����\|qcccfdd��-}p7;�ވB!D#��CO��ăU�?�KT�lhh�.-�� \^V�x!��QA�P��^�6x���ȭ=�m��r`��G�UB!;��*?Q�.�_r��C��288����+B�!�BT�lD������e7ɽ�"0�2���G�W���M�6宬��r�M!�ձ~�zg�W�S�xk�� �/+�F�]�2èˬl-R(R�P�mV."��A���Fu�,�:�B�*�'���ɶm���?\���
D�1��
fKi1�iJV��$B��"B��j,4�t1|^5�;�B�8`��
�F@kP�*�%�te��Ma��Q%�Ep�1(d)��r���P�l�F����6#c�^{tb�L��+0+�bu1�7fz��sI�=�,,�J��4�0�F�[%��ESk�U����c���ac��Cu�6�1vg�����ڙ�N�/!���tMǞO�7�����>�����O��ְz#o�S�+H��,!�B��U�娜_B!���ėB!D�H|9��ԀyqO��h�3=��ijR�B�ڱ��b�N����p����ק%�jD��A�����l����H �֍�MWǬB!���t�y}�i���d@=Ш�����[�[^6m��Q)�"=�s��on1++��Y'"�UX�6��0B!DZ��%�U_$�
���#�BT!-��H|����&�B�F	\�G�@�v��8U!Dq�]3�%s��!�U�:����#F!����#��t�9��bD}��* ��:}�^�ܴl�B�j�h[0�n~�+5�X�� �� ���{ʫ��_^�B!jEg��9��W���39�k�;��d�WxUd�ė���?}�F!�Ȓ��o���13sʄ��/!�B�������f�����\\\4Ǐ7B!D^H|���������Ao����DWK��1����Y355e�;f&''�ѣG��!��D��Af�ט7o��Zzt��q�q�Fsꩧ����D�c�����+++�ȑ#���f���f~^�B�b1>�o�c�v�x�� �� ���&����k�>�l�a�ϝX����ڵk��mo{�ٷo���/~a&&&�B���^on!�UXC�����\p��Q���6�{�g�B,e�k��Ç���?/&�p,�����E�'��������m���-���fii��^XX�zL�q��\u�U����҇�&�n�j�;�LEWX®��:�{�n��/*`_QW��.��s�������oi;�v����N����8!���X0:;;C���086[�

�`陙o�DcC��%�\�����3�8ì[��<��fll�!�pt«�0k ��Ex���yz��ຊ/��:�ZeP�|�1��5��Ƅ�.܌y[��`�p�5ט�;w��{�!��f�O#T2�yǊ7�a��`KC�������(���20
�T4�0X�l&�K`���K��7d���B!��%���>oxx��荤���	�Q%�_502�샚M����+�������9묳���g�1B!��.�e�)�.̤u!s_X/����
�"$F�O^ߥ�p�Q �H��T�l��݀X��"���� �B��.Ƽ�>����q/&,���\��˂i��]�8������,l�S���j@xO�+�H�Fȫ��j�"kn��ƺ�8l۶�<��ù��ƀ���5��\�U�e!���YP�Y�������#�"�x�������V�����Z�`����儸�:���>oz����l��[h�j�XI/����
/`�q�e�����'���BQkz��KsJ�g���/7L�Qoo���Q��\�S棌�!��0ER���f�ݝ�������9����ׅ^hFFFL���'C�g?��B�z0�7f�ī~?�{M�ŗ+IYķct"�/��G�(*�K_�R����W���ޫL���A��r�)�́K�x�0�*]3E�j��~��#�Y��Jo��	!�HsL\۟��z�P���|�<���e���y��'S�e���dˤ������3?���G>�X����F�X�~�9�s��e"�$n�ͻY)���+^�P!��H�g%�w�_�����̇>��ZFST��L�Ww#+�4��v�[��c�Z��W�p�]|��U�.V�Է���u�U���
!Dy0���\���������k��P_�^�m��>	���b�X���WK ��j��ə���^�}τ�h���Tް���+
]_�� Z���Z�c�s��A#�Y0=��4�����vo+"Qa,��C ��2���`_-/�a��1�b�x�9<>����C�`�1���7Lk˒q܌d*V2��Z&j L+YjyV0�ܐB�Z2��a^�ZI|7���ވ2B�J����+��d�w�������q�a8�F��Axa&F�`u������Y�� �`V�S�ݤ�o����皯�$A��{�>�7�N�����6V|ı��J�N��,Kv�X���
�Ū�/)7F����`|�+�Jߟ��<����5��[���>�s�����f���2�����.��]��%���,�q
�sv�0V�3ap�qNw�����\�bt�$��c�������p���r������m�/�o2�
<s�lT-\�a���ė�.�j:�׃��N�v��a�"<��X�zn���7���e9�s#��l�,�?zCnݺ�$�ʵ���Z �{���SOM��={���;w��{������Z*��L�Lh$������c�c��_��+`[K��ic������I�Elp��9t�پ}�I���������oz�LK��τNF,1'�İ2�9Gd�FMPƔ-�X���7m�y�V����]���\?$�׏~�����yˎ&��?��I���ęg�Y�9�����FKs�,�h)S���z��q-�����Bx��Z����@p�i̗˴����5�7��駟^袨� �A�����/��Yڈ���[�x׮]�x���1Ľ���n�T�g��B�a����/{[�sQ��~�ZD]prN+�Z"�7o�l��c��BͼJ�h&/+ʩIWI( 8�F+	�˱r��IK�p\�k\�mҲ4q~s>���wzǍ�����9\���Gy�&��ZA\q�P��<W����[^vsL���ڤ�Uj�5���8<�裡��_��_I�N�J9��**�>��z衇��? ��C�U;°�S��|׫.��VC�r�����ڜ�0b������j�v6��?�q���s�E%�\>�]�,U/,�I��/��N*�N;�H��߲�댌mzV��H#���-��++ś��(�\��ܶ׉��t�tm�N[T�	�QpBbR�O0>����?b(�����H"Rp����i��ā�p�"�2V����"~�1%�֭�UL8k�8㌓~G|�Ɲ���M�ӕsm�'�um�Nc,j%FE~���3q��Y�*�/�[����5�sl�z��f	%���qA��9?�c�"��$��s��Oa��9��m��w����Kr�{S0����L���gb�x��#��D�F\�|ng�e��f���wq����i31�8Ŭ�Hf����/W�LD��rܬt�I3�(�h�x�~������<��Ox0�7��V��pu�`饗N��f0�')���w�.�F�I�8�Z�/\XAa�'�Z�uL�!6
���[�{�I���{��ֲ�B �R�"�p�Yx~���_�L�Q�K�6x,A��W�����o,'� ��0�(
$����;!����,h�fLYPK�`�&%pm<��'}o�Q0��{��H�.�q����'���KZ�/��5�+������#�&��,�+(�w�j`�������++���q)�\v���/&N������@Gۂٺq�iku�'%+�(X��Bb��,��c-]��AX�P�g�� f�&)�����ݓ���DE�����
��up|�c�M��V�+,�:(��b�8w���⠒�+���G��	�(ga����z���=F�!�Q���_� AH��
8��~�K%���������g�_���=�8
Zu�&N�Q���x���U�t͔�����x�T��<�"���e��rs��e��6o�:�M���/=X�T���B�ꔇ�_<���3)GA���l����ܸm{*�/���������q_a"�k����6ޅ�3(�jY������,&�(�U�x���G�5��
�DW�B��[�"����	�5�P��Q�7,]�y��q����y~`���Z<-�'_-<-a.ް�������Yhz&L����31�c�;J[{���\��-��/�.)� .����q�eC�wi�s�y0�'���2����|je��s��獵�]a�$XO��M`2�:�l���j9�1�L���r�
!�S��e'�0���a.���6l���H����J��ᳬ�/,��k��Ձ�q��r1T\w~���ъ�`y^[��.����F0���Փ��_��ؐ�v�cf�L�`.w9̉�a�nG����cm�w��q���o�߮
�i�=�x����J��3kD0N⸹�A�.�8�?;,a *���6⫖rbs�M�����Z��z���c"W犉���	�VB1̝V����/�l��}^�WPL��(�'�>���la�*��B�}򚠋˲_�|nP|űXs��]�|�s�=�-H�.G�*L
׫Z%�k��Ms�Rz&���DF�	��OW�G=�2����p���D�J��j �*e�����tX9'���!&FpyT"���q�_~X����+-��+��j�1^a�&��R*���4B�ϳ����/i�J ��%��0q"N�.`^k��1Dp�d���4�s�}� x�����"L̇=o�Xvò����>�X�l�&���}�w�"����pMQ�&
�!�li�X�\�Q[E�p��*���LKMp�D�e�a������q�w&~�kՆ&�`$�B��,L2X<��&����p=XӅ�^a'Ľ]��DV�<�)4�C��o��:� i�z��8cUl�|�����ZQ�k�Akl\�⋌�(8����6q�w�}����r!���r �����⠥7w����cLc�B�%_t#�$����<���8�r�-��̌/�=�02_(>̹���pc�z�����j6ˊ�k�����K�x���'Z	�,X-��+N�s^����������5����-3���B��ld�U��#TE����kfu�n(�����[�Da�S~������K7�EÊ/^k㥂Ԣ%�;J%D]�<���8�J�k��F�9K��q�?�i�=I ~��9�3��e0�����y��	)�q`�y�5ל`��<q���"�+�|�T��G�J}R-܋n�h�?�X��V.�%�"�<���9A�8?��ϙ���j?ܤ�`ɨ�qZ?4R����a���|x������e�]���A|Qj��C"*9������ܰ�{X(�Qn%&'&�j�0y�w/�,U>�g�_<���w�*D�m���v=�/���XX�^_�OiTs��{O�0�T�x[�=�ҿO�i��q�ۺ�6Q�Z0�/ƁJ.C���W��§�]�k{96�m���`h@_���׾���b��6��W�x�%�e.�P�X ��-ܠ\����W�,G�2E�w��lE6���5h���V�����-�uZ	�,2l��Ewc�
�pN+�pq�t�Ғ�H�-V�G����`�9�Z���&w�>�L"|�	��( &)"+��ŊSi�&b��-,n%X�5����$���W��Ú֐;�q���"��`r�?�2ƛ�+8�C�Q�p|�Ɣ�i�㾌���i5sc��>��=�K{!N<H�|����!K
7p���r|��0E��r�7�����7l��C����k��Z���q�"8Wv"��H��Ͻ�����&J�N�a*�M�k����_�!L|����Ik�<����W0��J9+!�+̚����$�"(l"L"8爬`r������R�⫝̸�乊�1�|%.(MbNZ�����sïvl}�9�\\e5�g`��U.��7k=:�sB�6h�M�(7	0)[q^n�����T��Ek�t��K��z>7��ʾh\E�wX	u���<���R����EA�;<G� 6�G��
VH^5�=�\f��ԅ=?��8Dݫ6h�c��Y�{1��l"�յ�^{��)���5��,!Q~��+��cJ�BI��9��8��Z��ͽ�y�[cm.ji�V�^�Un��+�>J|�o�r⫞�^�����*���ײ��b=Q�
����Z�j�`g��(	�@����a�u��^L���!�G�`�M�p�?5�l˸�X�-� �.
1��.hɢ\u��V�(o�(� b�8'օ���qTQ��BP �-�Q�=_®+>�W�]�y��?�˕� �«R|�%?d�S�a̣&797���Wf$��(��ǆ�+�X�x/&]b��I��u�*����$?�#����LجT[ۏ��m�:����¾C��U��f|������?��c�t�L��D �� �(�Ũk7ZP|a�z�;��]֢Ÿ��0�O�vD� ��~^�@�(2��;~1<����0Kh��B�2��[ll���ĞE`��\�I��\�؃���A�ŠX���mc��*�	�����dQ���Ju���j-K��8ɘǡ\�(pE���r!�9N�3¢T�&L"J|�M��.X���5V��$QК���/� ��[~�d��]cX��W�-���0E�Z��2a����3��96�	�6V:�FX���~W.��+�/V���Ϊ�;�P��NK����� �U08���@��Q���}�6�&�8;;�q�!ZX�E%�^��.�g�'�rE�\���B1�z��T���f3F�ᩅ�������{�Gų�RW]uUb�­\����Qs+	dԺ�X�T�+�X*�#�����`��gas����<S�9��Ek��D�M|,���&`p҈>�Iγm�'>�Bd���VX3(��(����:��,�\lv�'89��
�56�&nAC�jV�U�ė���0�U+W�͂<��3O�=n�`;�ß�����'N�C�)�∍Jǰ}�v�=VJ$��gX��n+B4n|g���?��Om^l۶���z�=�����͕Q�-�j�u_[���
�����c��=|y�Z���A�_a1[���q'<й9��s�\C.g�r�cl�-��B'��&����������q��`��#��Un����u��:���*��w���3ߠR�$����?g�����[��-�e�|D4�V�"
���`q^qA�f�`����{�f�$
��$��/��
++��r,��,��{8n[K+c���x���(���ظ^�,�5�=��ι&�Z��V1�N�/?���"g[^%Ͱ[[�L{[<S��b�9�T�����_�Lظ��2�Z�����⽘��V1�V6�ƨ�<�>�ݐ���y��j�<��)�
��jU�.�����.1�@���4��=�X��#�ӈ�$ߟ�,�xq�{�V���T�hE�h���<�=��	ƭ%%ι��#�Yƃ�%������Ҝ/�un���lv?��0Yk�+��N�sN|���P#��}�l��a���&sx<^E߬�"&��\o=j�T",S.
���\J8B���rDJ�ϣ���B./@�Ћ��Z���u����aؐ�Ff��!�v`4�k_�}��r5���(���Cj\���F�
�!.�������H�P��B!�C�K�VdX]����p��Y[�B��+-����իB��@�K��0���� 	ľ������+���4Ģ0��L�BQ[ܜ!W9���ȱ!��>o�;gLSSq,�R��n��Cum��]^�R2�b�6���Êz
!D-X^i1S3k��b�Y<.I�i��[cv�eJ8Y*�6�2E�'m��/��������im*=�T��|@�&u�'�X%�.�ҸBT��r��wd���_-�.!��8��x��3=�e�ܴ�DÎ;�B�d�Q['�J�AH'V���͛7{�K��lw�E�R#-BUm!D1Ax���l3;�iD}��*�S�(�~��5)�N�b��c�A��1j�Ԣ�*�&�^^I��h0X���ǿ��D�1�{M
!�����^uF�@�M�N|Y�����K.���E�83܇B�
��[��l��*Ǘ�s���@P/,iS`� ��V�BWX-s��H|���Ƴ+u����T��] w+1o��%�p���93=W������@���-"2&�z�)�eQSQ�<�����%�p�S�����I|����ܼb���c�:�Y�-`�"�(P��Um�b!�Ȋ��q�q���;r��A��a:��Mτ9e��י~5B}.�2P3�u(��T�K�:����	sh|�LL����nd��$�d�o�lY��ijr�{= cAC�CW]��w�6�>��q�m�BY�9�yU�B�/�9��λә����r�&�,�`Ϟ=^��/�ܳ���dgb�B���ܼl
^[h$�Da8r�׶�����z��ǒ����i#�B�E�K
��#�<�"��5�K�,�_|Ѽ���*%!�"1_B�y:��aiy��C�cE�s�9ǫ��G=0\��v��b��)��CAո�����y!�� �S���м�駟6/���ٲe��eF�Eb�hο��(�;��ۄ[H|U�4��vj�<�W^1k׮�x�uv�o����޽{���bB8���7��dq2N����ς�Obz�������� ��_���M�DC5B�(pm �ظf����������]Olmm��i���눟SSS�lll�{�Ip	!����뿚�{Έd0O�5����X�a�sD��7:#���L��!.��쬧�U�RX�H"�ب�/�(L��z׻N��$Ȣ��egX,ٍ���I�T�S���ި��Uw�� tww����������l8��!D19��3O��[KuL���a#L@s�b��+M�n�����mX�� ���������_� i;0�R3��%)�"���O?=���P�zfz����[�Eoo�g�U��g�5k�xZ񟔺�/���Z�Xsb�AB��M�6y������X��L��zjU5�X��J-�}��y�8rM�>�vV�����u``��I�r_��������� �d�����(�(.<c;��/�,���^g���]H�.�#�n��Y,҂�� 3bΊ���z����E0������������\���<����c�5��������(�Y����o�W�%
�LNl@���d,]�r$O�A����g�]�s�cD�!����/4T��G?�QgE�mۼ�py��]S��*�����#� �M|�T�z�ʉ�}�W<B�V}6������C'�F�~_�&wj�&�u��y�(.q�W������?�|O�!������7+���כs�=�*�w$��Ϣ4�2�\�y/��M�G%d.⋇r5��Z�����`�H�u�c���-�UX<q>� ���<L��DW��El]|��mo�D�,��`���+���&IƘ�c8p���MA��#�`�w�yU�.$1��.�>��'�T����Wc=��������{��>nPW�^H���5[6��{n2��G�Y�� �P=���	p,@�
!2��,*X��8��ߗ\r��j/gB�`�b��%��ƍ�����V~��K%)�:묪�癚bO<�D�ɲ�l>e�Y;0�/�>�����CU�.ܯ���%yd������>��W�����Í�J�4d!Dyx�!@���m���|W�!��#��s{饗����0&2�X���҅��Z�#��VT��~1����_�,t^xab����5�\c��y�k�.#�	q^qC�~����g���۽�@hb��=��=��+=ĸ���~-�>n��V�s����5N�_�&D8�.�Od���C��%�ѭzAx�"���T�������'�B���$����A �l����c�yYDX������؇(V�r�׾����;�����?��n���ڥ�J��AI�%7�#�<�x����̽��kn��X~^^Ê.j@�X�`A`ʣL���L��&�,|�0�!���ܩ$%D*��H~���Bw�Ey�˴ ��O?��Qo����!M�v�CR~�����67�|�;X4PT�̞8��$��d��4,V7.��ťV33�i:;Ls� "{x� ���Y`)���Q*&+��cǎ^�"���"W$1avbc!x�СC�K[X��F���A���������Q�O�Y2m%�4n�$I{V�{�L|�0�g�A9���1]��21��m_Oפ�0|���qW,�bC0=n��U�D�6�c��(jXp2�K��p�(QA�D��
Fl����/O��"��X#3zl�_[� {p��U��2Ȣ�E�XtM��z�Ƒ%���q��qu�TKp-b�Z-ֽr���y!���EqE�"5�(�ja�#���B6�3)�k��)A�[v��b�&�M��nq8#9����ʪ�R�h)X���#�MO״�]�N�(.���T���&ᖸ��+3){C�C��rĺ�ʹ��s�x(W,�VTS'����g�}��n�ZOs�Xװ��n	Lʡ���^�z�&�[0�0��v]ܴ0��ȱ!�/Q5ܛ�d�I�D��9Ӿ��R,��ɐ<p��WW�D�8!ӎ��Q�o�5d#���R�=�G�~����{?m�KZ���ɖ�@c!�>I��a���I���#�p3Ԙ{tb�4
E��9���4��nv<���n�����B��dJ�f��"���J�t=#��r�Wڀ\�V\Z��g�!>�y���\�".8+b�lvR�3���!P̴��?�y7���_R�T�M�w����;!,��č�� ��n{��P��<�w_2fDs�m���r�bak:�^L:T��%q0E��δ��)��dC-6Pfb��!!j�uq-�q-@\3V6��˵���IY=�m�ԟ������u� �H�~F�1vEo!eio[4��n{��R�v���/nd���+���l!���4�����%U���`R��s���+�4���n� �w�Υ����D��ړǌ�m��S���±W]uU�LH,�;.��3�?f��`�"��aǘ��bg.�}-L|m>d��UnB��
�LtI���X���>�DIkx��dt�5
��`|���_��Xh���e�F�-�ĶI�ߥJ���~�3O�'�#�h��裏���nఙ��6�Sn�]����b�U|q��,�8�"@�������.�jK�\,��'Kn�"Y�,�S�)	XG���v�Vr��*	l�"�9眚�00����g��O[",`I��X�bW��Ǧ��u�./����3��n��Ja.;���7�˵�v)`��0|�tu,��f�/,�.��X�'Ya���r]���(D���r����id6m�tR!J&�I����|\�jq� ��x����m�;���D�O2��|OT�H���-o3�����z?�Ģ���g��"՗�_Wq�.O[ˢ��j��fQ?p�$��!����U����1n 7�'nF*�7:a.g�u�zl�ܕl�-��%B6������Xa	�E�M6���o����I�~�,H�'�l��Т�ֺ�m--��鶖9	�AΣ��E��Ff⋛���Eף}p��PL�W\�L�y�STp���bC@`�+Z<[��r���@!N�� 6�e�&5&>V�L0��?�ӊx>�I�)���M��#V`����dX�����5����WVI�Gס�����+�LKM��ǜˍ��O:U�4���T,O�0�H���Z��v��i�
!�����?�*�`�	���O
���I]}j����,�m<[��A2KXp���(8N��Qr�o�c�6�c9ū�{���?�/��$V�?��?Ju����*��#s�Ū����C�����,^aM.�h$���
��S�����w�K�55�Va�+�2#��V1V��Mly�aX�(X����%�J�uX���9����<�f��/�0���!��XJ�ވ�wܑyfs����/��N9����W�b>��T�/��q�x �>������R�b�"[X�+\F���/nb����,[-PU>{˳�a��S�2a0�++�7��'��:>��'��uC��x�g�W_}������k���a��:�x_Ͻ�7�7���]^)n�u�ς8֯[o��|򓟬*f�R��(�#d>�H�����Iji�����r���� �:�:�"�"���E�3VS�'�*�[�3��$p��EAEA[+�r����Tþ[���J���� L�|2F�J}9�E+g5p_���U"�R!�
g�x౺a�Qϊ�<ljmb����M�8�i�q�dτ�}TDX�Ѯ&XZ�:y��'DzV�(h��F�c���`KD���c��f�bM�+�
�c�s��V�X�\_����W�E7
\�����r�<g*yr1�p�Zd���Mq���mܚEd6��;[�����;�bjtX���X!�+��ڬ��ŵK,IT���\�$�X\��45��,?�ٖ�j�1�Ep=�&8w<��� ��\����'+��^�֧M�0�Z���ˣ�_�ĉ́F��X	b���~�:���X�(�@w2o��� |�!���T	������RJ5�Jn,D�j�W�.FGG��?o��7�s5׀%�� ˪��nJߢ��X��V��S�-���,N�F��F*��0w"�=asL=��h�d��(0���ʲ<��'X��7Y��_}���I^��-� ���Wȍ�q�ܣ�m�VY����S�F�Z�u'��L7W�s��eF\[��9��~�[w��uL@<�'����e>I�F��n>?L��B�[.��j����4��ds����U.�1����a�¤���A����,K��8�<,x�R�c�w��(}Â�����	Z�x6��������T�߾}{�8����OR��Y�X���!V���(c�չ��;i�w�`p�����1�5jm��ZAo�1�ԵN�"ʔ���<X�<���S�����7q�m����-L%���������?ʊ4Me���*?(����I�I�Dͯ)�Z.[�	���0�\�5E�=�H� p�㚌���[.#>���9k�޶m��Q���0��	���Kk	â��`�Ƣ^�"U|�l�P�7O����]m!3�u��;΄Cq˕�G7n4�z>.�b68>A�R��T����N2�&�<��Șв�9��*��<B�%�\�j?X����c�������,�PO�%�^`�ްZ��ҳ�*�Lv��3����7;�Z�'[���/�y���犚�
���(�P�~�`�j!�巌��'�T\o������E�a���I�[ŧ�̫���`SGAr.�4e4�gp?�_���T��U��Ƕ#��2�k�F�7Xxd�5�_A�ҫ1P�����8�5t��:36Y���hl���� )7i�8Yz,Ҳ���*a�(H+���>����&�3V6�30yY�C�m-���+���sc�s�Q��hQD�VkXQ�gص��Z?t���+.�k�f3��]"���l̫��i�ZimY2k:�Ů����*����Ji��:q&;bJ��wd5�j��0��͈D��>2j����͛�>��J��҆�aƢ�`�*�@o�0�����A\n3�޶{>inVu��p��B�&N;�F�ű|����q���ظH��{��R�1a���E����W^i~�ӟF
Fb�pA���O��f�S��������US�H��!
��8��)�/� �"S���|�I\�����:*nL[X�R�n�d��X�u��y�z��q<�Ϥ��96�1X��u�m�$�DRt�8Ȋ�_rQ<*e�Y�,Ò%��
&6
�,_Q R5Xm��8��+�ċ�3*@����O{�K/��jW$	�&��i�_p��>��k8����6��R[~4��`�4c����}��wO�u�GL[�b�Du�P���2TM��.*���ֱ�q�^�>,]Q1Yd�>��C� �[,7��/����*��k�.OH%m��0�kD0AG�=����.f�;͡�39�k�eM�=��7��9�ظ�����=q�+�u5�N�|�,	�r1n�=�e�5D���EG��0��(A��4qY�8u�}��п�]9�4��N?����Ͻ{�� ������l���NH|��f�k����/���d��D�7C�QDK�dlfI��-�y�!�a,a�� v
KX��0"+��kӂ�1�~$�Wa��?t��,�.?�:�Ic�\��DoN߈\T��WAX^n2�Ǉ��S�4B��;�u��k�%%l���+(&����x�ю;B݃T��jq]�y� �8��;���`P>�;^|�ES$��3��H|���d�6�: ��B�����~Wa�cS��h*�/�6y�!Y���@�a9
��s�y�(ىi�g�u�I��Ф͕9����T�]êV�n+�󫯐�kH|��f������ǒQ)s,nVd@p֪hg#�\<�\3yrJ�P����M��:F�Q���4gF�}���"F" -	��AAk�����%���aEE�@��YM[��HT#��.����e�"ˠ�j	++<����a��F�;��80?$�41���e��+���x`�Ԥ}���94�ֈ�!�U��8�_�U��&�J�)`��U��{�*�.���`|�����3�Y�q]t�E�5)h�p+1`��H���0�+�}�رĖ5�I|m9h&�{�܂���B��q0�2tج��v�'M��[�4���~�I��}�d���'������r��.��@$�!�jӦM�j��O�X�h%_��Y��r��0{�7��%���ɼ��r�������y��9e��%�Dy�
��4���ۧrxxxU�/���_�-g�m%�zťGa�|�8-�q?�9�J�GI>�J�Z�*b�O_�ל�n����1s�m���:�x�1��]G��A��缪�B�1g"�bwX�V�@P���d�Q`s5B	���388�e���w�O�`����c���{	\��� ���a�� �G"I��(e�h`#���ۘ��C_9!�%D@|�8܊�@|��E��Gp2!�����7� }-��+/X7��_@ :���^K��
+�JoEji�)���2���L*��F_�>H|	� 0�T_/�!�0�P+���*�����f���ܰA`��E %~�Jv$�F,Ul��jIX�T�I1�4�|x���?�p� �,E��5!�!�%D��$�e˖����p#�/bw�9眊�cL��YZem�p�����zf��6�%��k�LĨ���6x��M�� >m�֭����.��"�5h��,�$���ǄC��A&fz�+{���T�X�,_��������D��H�f%�����I��W\~������@D� �T�<�L���c�f]��N���-n��^{���{�s�F�a�_�'�}ű�ZȢ,b����3>�j7��$7$����e=��ȩ�A����Ê�֯
X�c��Q��	b.Z?�0�̐�V	,d�v�Y�p�b���j@�PA�W^~x�O��.�̋+LB!,�jc'%��j�3!���]T�\4?O2E��d���b�Y���
�����!�8�<D�-*��կ�"p��W�@ŁI���,���l���+!�*UC�"S��_��ZC��e�At%^~ �?��y�����b1(�vi��**��lRH�p�t�7���4�H��0�����,h�v�X�9%�X��@�J��j�b��d��	����c���?�8�����8Z&��5�Ʌ����LV�,y����b�p1���M��Iݚ��~�\��m�AnGp'W*��u�b�z�j�5��⋛���E�tb�����Y9+r��U�M���(�~��4 � V	kI�(\�b=�ЪzF�YC��j��s��Vi@�3T�ȥtG��Jk���e�&mb��3ت1��U|1�ij���ʍ��Q�����B�W.�J�8����G)�a%�)���
1bE��%��/V��	��$�q�^�����`�xX�x?�^���OS�k��6�1��j�<�V|����H����C�F0ҠjU��5�U6�[�.��5S�ZÄ�g��E6�j����x.b�*A*>�9��� ��fg"���`[-ُ�H���Vg�}vE�E|إ�^ꅄ��ٍ��q|�SO=u�g��mI�Uȳ����y��(�ł7R%�������j��ϖEt��fR�O�⋛�+�v����S���]��(j���A�Y����6���Di#7(�����
���^�È��hz���^�3�5�+�0;v��P�F|YO���g�.�\�I�Q[] �F����
���7���0�b�a?XF�zr_��<�3�<\`Ydu}�ӟ.D�c\}��#��Ϋ�Z�&ٟ��'��)*|_�ĉ��;_y��'�0��e�r�e&� �~��^�DB|\ܐ& zD"��א}�-gq�"�_|N�:vA��Ń�-�p�С��.��O|��D�m۶�^cYb��,�kQ��a���n%r_���!Tx(�~y(,,4NGz!*�a������x��W{�_E-?���5�\K4�,6O>���������F~Gƨ�dIE�͠�<@�k��!���+i?�9��D����}�Y#�盘���o-@�`��/����l�W����ŀ���~��Uq\ψ�����<�装]�`i����ȸ`��a��[��	��"��T~!��L���s�F|���H[�HZ�Em��g�&?�^,�dAV�f2?B+|�wd�ɘq���i32���щA39/`T�>��	,�[���u�]g�o�n�Z��/�1�q!>�L>J$L5p0�Y���1"�B�6Ԗ�I�@���ZR�&д��(Kh����V� ���1ӻ&�x�?z�YX��UWkp�U���e[�E�⋛��
M�]>��nr�89i7�}ތ���3s�_�,/���'F*�@�p�P" �.E����q�3#�w�˳�5j#nV�|�`&,�9�x�Pƅ�_i���j,_i��)�5��k:�|rx|����&iā�V��9�b�LD���\BO���F�4^^���~6�>x�bJg�L<�	>]YQ!V�:`��>����c�㙬��wx�*��?���c�y,I�7�#\�<���a5\n0W$�8/�� K%%|���??8^���hI�܎:Jd��ⓤ�ħ>��D�q?X�y6p-�_<k�{2_����y.M��?��?7��s���[b��Vԗ_�&�ޱd`�$�I�q/�"-Zx���g?�bޒ�r&��@��O!Ѵu�\a�E���L�"	�t��u����vCc����(���n3��on���;4P��|���u���'�O��`�$��j11?��$p�P	�� \V���%G�9�$�X ��c#��:qtą���,B���``=�j���[��@L4A7c�"�A®��V4���&mۧx �{�t9����tJf����\Kx�F����T�yqw���7��f��XI���!���aFo{����="���mc��b�`�Q�
`�K16�K��E�����u��~ܿ*�V�*�i��M�
ȏ�W8K������k����|�zl.�B�}�_��/��A�j���r���[�m��� ��_7]�-�)���^�FL�i`5g�A����C�`	mňKn:,݈��/�<�����ϻ08O��J�`KZ�!ʵ凱!�!a�ZҖHc�dL{E�w�˱�^������R][<Wϲ<��&%�ِ٨�<�����[�0/�q��`�K���1"_e�%+�5l6?����ϸ0%4����Im�<*q/��h�W�E��8^��Z��L�	fNS)҈/��d�7�h���/��Q:�ſ\��Y0�	Z_3_�,r׏/��Cc#f��F�Z���A�i'����`s���i�Y5�/ܱ�����ˤ�[�k��A\�A�֗#[��K�^�;$O���?І
Ѿ��8�G���o�E���A�cfG�j������Պ������r��;�u�ޔU��#+�/K. l���vՎ���f��l 1�MD,٠a�8(�V�"���*�;/)���������e�� k�ر��.�(a.;�L�]����KA�"�\�Z����[[�V0Jܜ}��^ }�� QA�q�b����4Ȏ���?3#�F�h�ѾX������$���?!@�ˎ���J�E��U�RοB(	TI���8l��x���fK#i4�ьf������g������ݷ���SՖg��^N��{��9��FV܊?�p�s��\�fEK�  ��"�����k�����k�U�a��1�^��Z�B�bC��n�mOD�!�(���"A[[��5@|�&i4����K�V3�w#ؘ8V��BQ�b��I2Y/�,�1?0	a�&�&�d�f=������$�]�|Pe��{4X��
Ta,k/�V|U-kuW�Y�jȈ�Б�� ��s`ͱ��eR�MyB>�Xɂ� ��U�:�#��f�eؗ�H��e�r��'\r�+Y�jDm��$M����.�?6�N
�Xo?_ܭ�'��>MDy��í`���l���U_a��[�3ȕy�u�V���1�6�5�m��+�2��#���EQ�2kxx8�9�����bb֏;��b�X�w�������㠎w��b�I	nhI��	��VUO>�d�I}`X̒�s���a-�q�;rё����y�� o�N&�q�@+�l�9o�.��3�x�c��0��-�X���V��%S��g�tu�0�=�����"7'�b�8V��ψ�%3��i'�mU��E\n�AQS�E��O��n0�A�1�"e�j���$1�U�@�~���?�v! �X1>�������b����?����w�~i�aIZ-L�^��ןj�.���V��1�\��ys�D�{-���+�<�Ub���n�⋊�6��ٖ�(��ھ�5g\��U�Nѕ��O�L�0�O̚�l־p�A�X?�4��!¿�!P�����$[�T�� 9��&9�믿>�J�^�B�+"!WO�!�k��B>�NX�p�rN�z�&��,��C��c�%�Z���c���>׌OTk%$}G#�
�$�.��["n��ŋ�V�Oe`p������Eݣ�9~��t�X��Ǻ������?e1C�R~��m�a�u�`+���w��7�!tB�;'>!� C��+���W&.\��`e�r9�p��;wײm�Vt!��r�q$n�����b�:,O
_T`
$N����b�J�apLJY���Dta��%��76n�N��<��ӧ^���� �AT>"�뮻.pe�]f�i�a@Ԥ�5�}�s�=������M���6�Qn_K_́��n�m���4§���v��"��`�b���b>+�,����w����It��Aa��'`�#�����M0Ñ�*?tʸ)�\׼G\��"{�]� ����ޮp��B��-i�UaM2VD��_���@�1i�@�a�"�m��?.�<��\��P�l���X�d�>v{�8�n�)w����#W�EcE����#���7��е�I����U��6>�m����zl���ִ`��ƍf�љ�iF�(�`�x�'!��{�gR4lVna-�
6�[,B�^�;�����u�ƊB�G�T��R`�Ɗf��q҃� ��bXX3|��LM�%�'�����;n.8����?�ӆ<��&���=�G�2�aЊ���y��-Gx�,��c ;�9$I(�"�+���0�ؘ\y��x�ħ`Q#F7����	8衇2�BT�#����f�M�ZC���hG�0}1��`�!��_+�l�>��X�5��w%�b��c��Ct�Z��=��ў��O��IQ�T���8�ǟ����@oDw�� k={�����4��8��Yζ�_��_L�җ�*h��*���a�.
�	�����s�r�Ă�Ti)�"�b�I"�Vl�B
kGY�`�!
X�����W�X�;���f��fR^+	1r��H\E��PK���W_}�i1$w�1�؛u���Ħ���g���k�/��D��	�j��UV	oE�U#�^^�c�&F-*�h-�Jl,��ʴ�.N,Ya����i� C+Ⱦ�0���/+zҬf�:qԕW^�` ��5�H�	a^�0� ��$2��UD&��>��\�l�-��D���Թ�S�pmƬ8��Pۜ�>jY^�Ԭ����z�M|1�"f����,�G�������Ϩ�	�xp�s��	=�q_L��H��آ�'4��&@�>!��`\�[����`��$A�i� �T,�L�U�X*\.�6�-k ���{�6f&���?�{�J ��Uq:n�^�C�M%@��qѥ�r"
�����.�u���Ҕ�4,4��
���[i�mm���n���`��+�f��+X��0\�X�x�;��c�M�*���Q3�B�j��"|�.#Ώ�H3f5mI�-���,6� XW�l���p�꼲Q�{$���K/]�;�Ã>X��<��w���7�.���??،Z!����E�Oi�4��G�"����nd�j�N�X;801�z��9�2Q��kW�\_���n��6�$����#)'ܝ��ܘ��B4<a6�:��O\!f�
��"������@F�p��l}��u#ڍ�9Z1���Cf�ƽ�>���fsh8IB��B ��3�\Z�&�"4D,`��pc/��2s�]w%��H!�f��}f��#�>���s��D�-�nP�56q�6֐>���p�5��Ⱥ//��r����.h�q!�Mm����~z��1������B�rb9ESJ�%Z�.��Q@v�VX��rz��۶m<j��B�/Qg�uւ�q1#N�	*��Y��y�'���_*fK߅^�,B!,_%���sbr�Y�t´��F�,��{�I�ː�����)������L�ܬ|a{V;ZlRI�!���l����4���f�_�H|��cc+���m��u7��.8�8��5�j�f�
-�?�lǻv�2[�n]�ѹ�+�%�(C#����5fl�ۈb��*1ssmfd�/86�=0/��*��ٸq��#��JU���%�,+�\T<���?o.��S�[�zup?l=!�ͧͼ���y�U���	��������5VIA�n�6\����k蜤"��L{�qoH�������5L�KQ�vIx5��
qdd���˷z��A�$u�[���l�UF�?V=����m��SO)���>6`Ds���DV�n.$U�V2�:��Z$�Ki,�Å�����ݿ�;�c�k���X�n]gτ�j2Y!D�05��?�!�U!:�V/bď�:rda�e��tc��9��[l��Bl!�HgᮨL+�\x&����ݹe��/!D�Y�d��L�#Lc�"�U!�v�j��%ت������+�
"\x,Ė=Ș�+V�܉�w\q��<x08��Q!�����f���F4���@��=��j�傕�ꫯNu.\�,�FĪ��ޞ��Db�Bp%Y9���4.��\fq@��
��N��(�ב���m�.D�Y��9>��4�A���q��A��w�T����vzD��'�n���Vf"�]�
�Z �Y�-D⫌ ��;�<�cǎҋ.�O>�|iBd 9$����9|lM��qbj��"�UB�pm�\]�fIG�W��_+7V���Uˇ�6�}\QB ?nD����`�����x�UW����*`A��{�1��~#�h"'֮<Sӝfr��}���_�?_%diǴ�]^N�IR�\W,En��+��}�B�Y�>�Z����a��dU��a|饗nH,aB�l�\:3�3K#
@�K䊿�Z.� \�H���U��.��ZX�@�1����{G�??���F!��ė�?n�HwbX��;�
�$�`�
��u�>����W^1U����_��\{�V�����Ζ_�!D_"7�z�)ʘ�u�m!���d�e�'o��g���l����^��f��BT��24����xv�Z���.D������G�-�E��mY$�b1��Ц`o�8��I�J���͵��h���]�W�7��~�䞶B!���,tM��F�GxQj;��%n NH�+�LP��Q�X�Nj�p!��I%ėƊR&��g?���{���� yh3` .���!]�SփE
�߹g�m�$D|��_5O?��)#UZ�xn����F�FBfם��ALu����
q �hU�T����b#jIW����.��4��o~�#��oڴ)8`O<�b��U���1Q�}a�:��}c
�z�>�YV�~)�B�|>�q2�SH���JG���I�\�����-I�Ht�0�7\�_�!�	i���k�
}	�m��&�k�����ե�M|�����͂ըj<?[n���#}��j�>�}�����R���,�v�[�UDC��^R��,���|�~���?��?��릊/� \�Hh�XT8�xi;N�=�>�n�Q}^~���іi7n<m�� +������[�.�V'�ݲ����?h��b��3�8#�I�0(rV�FA�]r�%��Qw�=�����s�1+V,\��@��r�c9`7ʓ���'9�v�����������잇{`��3�<S3e	;*��qx饗̳�>�7p��c�����u�� H`�y�{��q�����w����j�F���}sP�h��b�)⋂�Q�1�js�����_�LT:xW��Y��\s�5>�2͆��+���:h���лv��,�I`�����7����_�0�;.e��D� >à��N���/k
���:+La�{�"�x����L!h	U]���w�/�%��/���D��/u�V�p��P�Q�D���/�3���/��z�,v(W�`�m���h�A'5�ނ����,��c��3;P�I��]p#0�H� �^0ͦ\y���_d��L��З0�1�a)�����;�;}ǎ�,�j �����+��������a9���A�N�c�r�1Q�˅z����r�/�z���,&7XH�i<ן������.Vk���0�1��BY'��P�E���ZT�'[(���pC�z뭧�n��h��1/�k�BR�Eg�B�`({
��M�K�D��s��燊/U��������.΃�������7]�[��
�.w�M��P۽{���0>\t�E���:�X��w�Ł�>�䓧}�u�{�i�A,\���.��"W$~�z�Y�Z�w(�3��\<�G>����L�]w���,��'qM��~���
_E/��,}�zu�]�Yv����߼y�錉���:�}R+֩�;�U��0�N��ז����X���g���s�*�1V\���r���V���2#~(�2Ŵ���1�>���C�{�9s���/�|�>����K���Zܻ��ݾ}{�w���H�'�܋݌�{��0�0I�;��އ�� ET��i���Λ���N����ϔ[��	�+�(s�{�9j��2)JxY�W6�&Ny��)*v���[�K�
��3���8Zg��6ϲW|щ�)ȅW}l�m���Ѐ�V�T3�c���0AÒ������=[�]��V-�㮨��VO|q�*�W�~@:.Zw�v��r@tZ�	n�������,;�l�-�P���\تh���y�ٯ�|���Bx�y/�NB�>��@�����+���u�\�/���LL-3U��7ʟ~��u����4�BD'�vg�eeIǌ�X`IG�&qf�V|�`�$�/[�lhP�<�H�Ϝy���͠�[9�V�Ur|5+_�X:N>�
���8le$�s8�<c����ݏ�+߰�Q~��lP��"��v��n_��.L����ܼg�*���D��0K�_'�kܾ���b�'����]u�(k�]^�ۖ�"bƗĴ�'�a�1�6�:�X��p J�E�6�+�8�d��(&�5,)�%`1�`�բ��Ma���R
[��I;��SO|��׿����N�-�
��L�7�-��߹�dXPt�w���:�� �|�%��O�����+�l�Z&�F�հ�"��EX)�VC�
)i�03s�MG[�c/�.�+�#�eX��.��P
����Χ>����P9>wQ,�yr �3ͨ%�UW�;C��>��I��-۴3RNgS֘�(l0�����a����^�4;L4��.^΅˲,y�#�y����n��(*,�߻���fES���:��M�T�;B��q|�8�<=+a�q��k�Bw���1KZ��P\�'>�`�W#���gM/�Z�|s_6�q-l�3��7)�}�{����}�}(��1K2 N��j�*�Ȣcr�8A��&�x&���\U�W��U`��M1a��0 �����RY�9����[D��>*>��IrG��Q��[�X���{^~��s�/,�P�x���
�O��u��A1mx������X�
q�1�Ɯ)�°F�:".6�}/�G?����s�M7�M��-*Is�o$Ia0H}��L|��4�$�v)�2��##fht���0+{G�ڕ���%�q5���ź�5,�K.m�	���ȹjM�����v�,�</hO�� Z\'�3��*[2���<Szvŝ%��W,@�1�$!��Uk�]�=G����H��]�6I��Q��[��'KQlaL6��$t�_]˸�$���v�_'&�̡�5fd��LN#$��2>-q�&�!mR�� �;�P���Zn⋊�HE���ʼ1��\�|�X�Gט�w���/����]Q� B�Ro�<=m�U\	��Be�AR��Eڋm�\b��!�$�]�ݯ\W_}��{�^�Z�:�C�D��H�i�� &�(R������:]o������B}mt�]5��~?�\�G�0�Z��V}�4}qay�xbA���N��␺;�̝>�<���?�!k�NY�������^ 7�e�,XC��
��m7/���\���VU�(�ɱcapA��%J�����/�>v���'�
�2�c�1j��wG�ZX�lت�(kVh�g�a ��O~rZ��`� ��A ��V�6��`�Y+(9i<l�>f9�ef͊
Y��ZLbe��^�4<��c�='���
l�+�%�6�m�%�!��}�s�7�7�V�6��9��*T|���e������63xt�ٺ�ږ��L��$�� ^����wP� ��V��Y���������Y���f��2��IĂoT�*H�0��n,�ˬ��{؆�M��e�[�\��$��VyfuK-�.uw�/��Lu��&���xG��e�@��R���a6�NO�RU��V����V|-YR� ĉ��V���-oy˂N�X�{ｷr��S�.���B�N��Vs�tOQ�5X�ĺ�"�l[D1Pb��;H�_=�L]u� �����u�a3�ZP�������lXx�=���n�=Oعx����'�����9�n{�.$o+�F��Mk���:K9 �O���3K����r{��P��<�_��˾�n���7BG{y�i:���
&|6��R�{D�?���S+��b ��+��Z���~�Xb�
^qr�����0��֒0KH��a}VR��[�� NZoÞ#,h����n��P��hr���5������arA�$��{'E�Pom�ţ`'�~�O�91?1XxO�f�E""�0�s�_�G�͔Q��k�ʦ,ap#6��T1SW^ye���L�$�`@������Z��_~�47\������J�� ��k/�bU���s�6��>�;�_~�vā+(,Z��.v���n\�U�b����a���U�@���D��"���������W�#��}9����'J�I�k	2_|C3�PON_�����	r�U���Pn�+��6���f�oȴ�ڍa-tf���˼�p��p�=�P��3�&�YV�nԹ7��M�RX,ȣR��~]��o��1&v��JE�|�d]������`#mұ��7��_|�X@�5��P���Ah� ֊��M�]�o?���/�R���u]�P�|υ`w��J�7݉������C�G\WX�7ޫ����:ee�&��&r��NϾ�i�A32�W�}�
:#�B�h�WUH���V2W4m�c�`�z����;�Raf�$,|���`�u�Ug�j>���2�j1k�~�jlVd�J��J]7���&�e@����\����C�B ެ�E�`�!�;L&ٞ+Op%�����Y���!V�f+L��}0�UĎkEC�09�@��₸<���D��;P�XFX��M�)�-��ɖ]u�;��܏/�y����jZ�*L���w�s����b��p����
�3l�&�wUwȢ���漭ϛ}�����UN7Q��<�s_T�2���º�N����f��Iӻ�$z��Mǂ��L�[QF�MY�Ed !�����Θ%�E��w��^�p�(�A�,�XY��$���??���Z
����'�qݣy����Z�a�%���(B�x47���X�4��O� ��>ŭ7�%�t��zjc������
����G�d�.a~ǳ�Vϰ �NX���C��t̘���-�^1�O�IVY9}���.Y��˃B�V��%^�X昢�'���Cf�@g��if�� F�!c4���t�0Sf�6�Q�I ��w�SS��\ޏw*�&anL�H�6��L�퓶�[�|p�bю��"��E	7�7牊�b"��!W��}���`X�v��i� ��q&)�����������:Y��ਭs+e:�2g����ގe��a��oXL�(:ufŸ�Z-�4�y�~�rB��6���˾q4�;�1�P�M��*�
��yy�e��u���v8`�o��^Y������f����,�]X�fJ6ۧM�H=���E|ba����� ����V�,�vX���)+�*�%,P�kp���/��)��Uu,��1�&�in��V�g.s�S�kӡ�l�xQU��/� �l�債�����х�F��N�Y<��~���71^U�4���N�p��6�e�5��r����h�u',.���Xkʝ���@�B��1��S�]ToTV�7ܰ��(���C��ْ�A���:��>��$�83�O��2`����z�<����Ħ��c�+�D�~�{���i�'�7�pj3q�<���Iӓ��iԤ��D��\c��|+�`(*_�ennq&�,;�� �̙���k:t�̊���e%�(�<0��ߨ�b�{����s�C�}&��X�������� )X-��p��5���(�'�h�I#�wx���%�-u?���	��@y�K��j˹:w���_���-�l+�|F������2qh���a`�`���/:V0q �C̌�J�z0�ff�,�Aε�%#�p�Tq� #�� \�t�`��_���ζf*!�|^��W�8LVt<�o�ӾԃX⼓a���]|�e$vA2�^v�e]˚`�Aa�}�0}rip,v�P�����މa	��@sEu�����	@\!ܘ%ŝ)Q��5D��t�g�Z�0�S�[T&({�]�U(�%D2&�������jm�ׄ0���|��1,���"�et���|
�ӟ�t�i�8��5�ja�Z�#� ű��������̬�Y�U�ՙ`�h��^Į!D|p�����[�_��_�	}� �j������`Ѩ��E�
�2����|%\8T�"ݺyaE��,�h��N��E�XO�,�6GiI�AQ>�����n�zK�}�5�4{�#�\ϪVȴk�Ǽw{�.��c��p�j��B��  ���A�k�Y��g��4Z�߈�)��BT��2�_i��¶Y*
Ɣ8+��9,K�N3��%ʢ��ԌkЦ��5Q�O��d➶"A�8"!�h�ۙP7#�����8���7U� ���)�Ģ�zV�%�B!��z��`6�J\�I�Ѷ��Ӱ"����XEp'	!�b�`S�7���:y�ķ����CI�@����K�	Y!��.H\��r�+�#���޵��3'�qd�s�a�.
�UE���/�2r��27��B���|�����s�y���v}�Rx��kȮY��A��A!��&���9�%RQP8i
��G�q<�E.�"h+醣B!��Ee�ʒK+eed%��#O�izJQ*<
��f '(��砀8�-�,�U���DOטY�2޾hC#���x�s�	!�(+����xi�^=��LM���*X�8����0Vã5����j�Z��_.��VNl���I���H�ώOtI|	!��w�X������_D�b͠t�K!�����B!�(�/!�B���*!���������e���w���3Z�(�"Kf�:��H��3�S�fbj�� �UBN�t�=fl��>60/�&̎M�MW�6NB�8#c}��g�铋#��lH|U��]湽g��?k�t,B!c|�ۼ��L37'�J�����'����k̦5�B��W���j2_���n#�B4�؄ƒf#�U!���߯R!Dk�\�G�B��"B!������YiD���l9�v�a#�B4��ǎ����#���W��5���1�F!�h�eK'�y[w��l��#�UB:�N����k��Z��B!��q�mϙ��32�k&�������̶�?_%�o�q�}�^#�B��\����>׌O,7"$�D&����;v����]���\���իW�M�6���^�l�2s��I3::j8`k~V�Z|Ŋ����qs������wᶵ��3�8�lذ!�����9z��y�����d�w�G>�233\�c||<���k&��^�n]p�|K�.=�|���J�|a�������/�ߡL�\�g�X�|ypm[F���7ǎ[�y>�y���矘�0���[𻎎��׮]<��&��5:y��+W�5k�ĺvTY�:�=tw��D�ĉA}
�cXݠ����P?�Α#GN�.ף-��ߒ4�͋/�x�9����}���,�u�{�P�#@�P>aP�x<��Ԕ����:;;�󌍍��=�k�޹[�������sֺ��aϞ=��w˛{�=sM�}ɒ%�����9j�\��b�(s��:���G�Kd��\��:5�K.�$t��Sݺuk0H>��cAG��`��}�a��@DG��O�Ç.`�ýꪫh��O���_�:t������<+��3�<t�i�>�;�`P�a ݲeKp��~������:���Cx'_|����9�o��~�-%��$��wꊯs�=78o����ɀ�裏���W��s�,����:�;v�?S�^ޭ��Ԃ���}��'O�/~w�g�Ѳw��@p��}����Y�������߽{�)�Žq�ZP�������P76��{���j	'��K/���zF�3�8�s��~���C�9�����_�;ʔw&$�ޅ^X�h[<���C���7<?�Ň�FDR���_�]�/Ql���7-t�`f�q�������ZЩӑ���x��WG~���o|����{+VR�>:a�#ZLÄ��#�<r��}��G����oxC`�������S�Q�</�ʠ�����d	��3��+�^�U������(��w�P.�$��9�wI�.e��q/<�@��ƶ�U-����^��(��sժg�Q�=і�@9S7�>�պ�'���w߽�,�7���+��2x���ࢺH|����n����X�e��V��N�����Ε��������]:G@ĉu0ȼ�u�3���/MZxNf�X�܃Y��ĵk݀�������_�K�i�2۶m�����u=A�XV���=�\�3"ɵ�" ]�e]�.a���i&�5	�Vgiqˉzh'1����%�g�������DV��
��ׂr�*�z�>�NG�@�`�x�����Ym�]_%���9��%j0����B�j-\t\t�an��۷��B\�'��4���A
�f�G�|0p1buy��|�������M.6F�A�ٰ?H�{\�w�u�i����L��e@���� �A{���_��׿������pSFX,([�Y�g�n�0xgn\��
��.�u�AW�g��3eR�;J���w���B�z�g�D�B�^�:��]p5�NC��")���r�1JQ��%�����5�����<�_�(c\�v��=ߡ��Bw���X�/��RЖq�vw�"����Q�yo����� ����빗0�E{�����
V�6'�<u�H�52��\H|����/~�S�Ǎt�}�-����1��Yw��c�;G�����}��+��]����b C�0����&������E]���&�y�Ν&	��wಿcPs-����G�vC8��a����uDbW�A��W_�65{�Ϣx�[ߺ�g_�q����w�K�mo{��拙0x�����-?���Oѳ�>�m�+�V�K\��b���?~�/��{c"cw>g'+���{Ԣ@0�e��%�}�aψ0q���ow�;&0�І�:�h�E�
d�%�vw�W��e��C�������.\����O��073�ߏC�w�Q��⸱E�#�� _�җ�]v>��O�^��0�����\atl�,��#|w%�?���}`��-:Ḣ��1�a�` r��bo�
x�5�,xW?��O��08�3w, n��Z܁ú<mp4e�p	[����µÂ�����w��=�۷� *Þ�z����ǽn\���Սa j������Zr���
d�v�bخ�s���;���.p�{gW��ж���Xf1.E��3��yܾ����Ox�7~���Z⋺j�ݷ޹��~·2�ې�Z��_�u/n����/)#Y���_̢��h�k$��Aŧ��٧u�dA� �P��NY8�%��{��%�=,�#��~g�w��
��n&�@�3��0�ET�8���[����4����˖�^g�M2h���'k=��V�5
�Ǒ�@³!�\���i��(�Ȣ/t��1��_�F���z�|���<�����rWmu4����"ތq#*āɏ�kL��g��Yk)��;*�����mI�.���6��A_����8�֒KὺZ#˱�4⋁��@%o���k�0��Ē��û��1H����$���$�����o���N���	����(�S��^��b��qp>�ϜyN�Ք�"��F��ւ6*Ƈ~�Dy����u�]�|11�*]��>�Ν��w�s����6W��e��/ߚ�?�o����E���BP���n���U�M�uזG��q.�)m��ƽ���V>3>�NTx�z�C��f�(D$��L�樷�ڇ:B;�h4g[�ŗ]Ꞵ,(U��a/��Y�x3Ww����2� ��V<V~����X�4�N�{s�PT�4��+�����b�a ��G ������fה�;�"����ػ��XL��������.7��A�t���q؄��q�L���w�.�P^L,x/v�@�Qv�E��U_�$)_��_��_���w���~�o��-�Սs�ߏ�7��ߺ�����]��E�<qy��wh���[x�\�,�Ac��ia��A]�����T�c��}�,�48�'�\�n���8��=�(���d�&�<i|�����JV��f�B��!a�n[h�y� �A���_�6!JZ�Q�q9ւE����т��݇Y��ĉ7#p��8�6|�e-5�.V�[���]���9f���)�@�e�� F8��x���]�b��m=σ_w��巧Z�BL�w�Ro�p����;s]��{_|��P��, �Z��t�f��z!"[ho���d#��᜴�4���/��7����K[(�8�~��3	������Η{"Y+��o�q�;����w�;��y��]�	O=�TP�/w`���|�7��]���^V1��*��Bd�Y۹/���Z�⬀��:A�^���6�'���}��W�`�q-�a�/�_{��_W�!�\q��kd]1>����&��~�?W�{��I��@[�:����;q�	�{�e��J���a N��t�7V?�3S�,�i=k�����a�â�$�c��� �e��Z
��W ��7��P�^e^�lt��J�̳ޠV����4Z�:�T�Y�N�c6�f\�O�˺VV~Y+E��������0��PnT�5�r�I:�w̻�^v�k��V�E��oic�(k_�q]+�r��x��fQ~��B���(mrU�Cz�0��׏z^�����ݿ�;���z푿�&����IbL����sO�w�{B���G�[��ix����e��;X�����e���D�~(�ǭP�EA�݆#-�4(t�+*������a���?�����b��s��i�]1�;+�n��֥�[Y��{E`��7�
loa�p�l<�T��m4�<���>�[�<OR��`K*�(�.+�C������1�v!��J`�P�-�Ą��	"�we����W�G_�����\�_~y�~����������W�s��]�#ޡ_�<O.;�받(�k㎮�nˬ������hP/ʺ�=���(RxYl�i<
qƇ�������V̴�����4�ˏ�8?�c&�ʙ�'N�� p�F�T��Z��q!�����?�C&mwYz�@�[JIW�5ƵlQ޸D�*krwA\����9!�lL�]��~��mT|�u9�_���}�l5�#�A�B��\kH������ql*	,�ĖE�D�[g�+�����]qf����w���}��>��X������^�^k՟��:��m�:�x���R4��9���D\���7��<��f�{��͏)��VD'g���!{~�^Q��Y��zb��R��ZaМf/�b����o��3�6���=7�V|����ǌ1�2Q���qs�$��i@��ua�a��e":|wIZ�,+��.n�~������v���eŗ)��H���%�ˑ�̽w��D� �=���()��.c��$Τ_c5�����b�me�	#u��MWP٘.�����8el߷=�򖷜�ϊ�p��NDQ�&��C@t��s�}@����[܉5�b׵ǭ�X�\�5���r&uqb��b`�Q�v����ݕ_�u�.�F�1	�����O��{)33�e��q�cK}��<(|���F`Yͳ�*���c�������a�,��t� �w\���p���Ӭ�c���_|�iW������w����x�8X�f�Iٺ��u��$�V٦q9�~��\�ȝw�X1��X�S�DL�k�A�y�+��q]Y��c�U���bݗI��O]+%�d_|��x�G�E(lW�Pw�I8+J���.І�N�x&W|%�)h�?�'x2��\�y�l�b@kĉ����[S���%��N���0�Va��]���w��Y��я~����?4��rK���c���	K>��` �;_�1*�Z��׭�����P6u���������$X��ٽ��2�ݿ&�]k{!,l���u���<s�)`lἮ0�c#��oABt��#t�D(�ˑ�^,HISS���ϩ���V��;3d��������͵�����I�J�/���>'b���Z$i�X�{�^��ޫ���..�}ӆz���I�+@��Ņ��{��0K�XS7�>�_�m��Fx��RV�&���Ơ��#����|�|�s�37�xcM�8}}wT��U|ёǍ��&h����c D�6�z�A�J#p������v�X.��"�:A~v;x:|2� �e���=��w��{�
3;[AW�v��S��4
��n3)�����3����s�<�	�b��[�DE��x>WH ���"A����������PV\K�P�-Jq?�<Ζ(��%�����Y�x7n��0��&�x`��X�x�J����$�yL�l�d���/�(+]�XW&5���GQn�Ū�/ʆ4-�Ѣ<��X���������Z�(c6���������:�����c�o���.�X`��n���BB �xN��!���I��[�w����\�W�6ͤ^������wps$��3j:����It�tr�>w~"�(��������uIFa����R�s=�]+	>&�4��/��8.R�8$_|���B��� �	+W�d��b�?/���q\kv�0�\�v%cԾ`S�}�oe��U]�DVھ�n^���]�8ǂ�o]+7����]��u�&��?�Vɤ�^,�%J8�_w�&X��ׇϗE|��\nF�z��t����vs����e��=+�tDe��M|�a��+�e_S˂�5����a�u�~��޺�:*'V�k��6U������~�[�D]��(i���4֙������Ɗ��`�����F&�Ѭ�eA��`J��m>7���UވW|!\�X8V�8��\�>a�[����Uϰx�7���$�β���}�3:�k�N#[�	�cƓ�����W��Jā�m��(?mfhdU���3�����6�,3�%��=�0���]ѱ�ЏX�0��T�Γ��#��~ě0��jS�$�_��3Xo�K���qK���|'�����u$�˱�R���g��)�"L<����̏}��l\�l��2�:�&��n3q���JL̹�uU+���^=�aq�tJ���"���F7Un6X�v�>�T=�����@*���X-	�_�1>��>�Ƭ[��k�Q�2t����cf�c������t��X�l��0|���|�~��w��4���1ۍ��[-W�݆�v�ρ�b ��a3໢�_5�l�޲u\<�]Yo &0�Ga�I�k]p�6m 610ڨ����;q��V°�LY�����?3��,�X}lό�䙣�VR��4P�g��f����(J�p^�ZuN&��6,Ζ�`%�$��n�NhC�9?OX���~	���Ӷ)kʼ�����7�V7�����#I��Q�gK��5���ʑ-#��hV"�8D�r+�2�_]���)OF��J+��T�b��`Z��7In7�fR�z�z���\uV�փ��/�����Ө{�A��mW�I�%�w�x�[���ǭ����lYmpN=C��Y��ⶁ0�֑f12�<8���},���qXr��4��ɒ
�����JBњ�͕�R��*�兊�2����F��q#�B4Bw�x�X��0���c�%cN��f,�1�V�w�	!��q���3s��~���&��y�F��"�׎�/��[��0B!�K����̍���[��l�C��Q���a����Bܔ9��⫽}�t.�~-�j��;��)&�B˪�a��}�96`F�{���23ur�P(��$��
R
M�ʲ�2��Z�*7�U��f���|�B��,�8i�<��� �Q�(�Xn	�����QʜhuzZ.<!��ʠ5���*��H"�$]�\tǎ���ֺ�tCn!�B��'Mn�4���L���=cs_X��kW����xG��|�3�I��r���B!�(�"�F|��?��}�p�l�R���j��;�m�ݖ�vO5�@۽���W��:�i���ߤ&����B�\��;��̔7N��/�F\���w�n��kw]`{�Z{��b.�\ŗݐ�V4��w����C5t-wc�Z`��R�e�]�[a�y!�������ʰ����|-~��{ 7��3�I�_�� �U|!��8�ׂ�`o�ᆆ�7�?��B!��h6�������C׫��$����'��X�W���5?G��&�,�^_��WL����O~�f��֞�!�b�����y��L)*����ȈY�2��]�x��Z�����Y�fMS�`"��^a$��Z\ ��cۑ#G�b���u?��^��B���ѣG���@Srq�����VhK!!�B$�C�f�����W����!�V�ZU� �«
Yp�B���S/�)k^ĕǡ0��a�P�pA"�^r�	!��b���OX܈q�K���yq��!��ߟk��_�phe�B�� .�Ev荼>w�NҴ��/��Y�E�,W"�P�����1x�e'�6OB!��{��󶷽͔�_����n��_��Av��
;X�p5�1�4E|Y(̂�NH�=��&Q䞍�O�.km&UH�!�"1��M�E��j��O�M��=��=�	]9W#���*�,�9X��5F�\���C�f9p�׵�c�t.�'"��;�əR�F!�%�s����o���T���ZN�ā#������(�Ęݸ��q'+O�Fm�MǏ��P��lA�r,W�1�}��X��sp�94��!�>�ڕ�r�=���`/�V�`�>�?����`��˰S*��Ã+7Wk�*T22󯝅?�y�fs��g�ք.���(:U�ŗh-�I����~�3�gϞH�%�_q����*S'�B$A�K�޽{�W���@t����w�mx���w�Ӽ�]�j��B!DH|����e�ȱ��y�tw�0U�O>������xSs�������o.<[�B�:��mfl��LN/��QI����3v്A�.�6�u���T�EO<����>���G}48Ǉ?�ał	!D��u�W�7��W��Y��E#�Ur�O.5{7��'�͎M�M�8x�����LV�>��3�����y�{�k�B���잳��Ʋ"�U���4C#����aS����-X��(?����_nv��a�B�����$����W�8:�_�E��$��;�0�7c�B��ɼh._�J��?��Or9/�n߾}f˖-F!DrN�h˹fS��\������l\��?�|n����%��"%�%�p�C�"�����"���ܹ3�l�O=����?�C#�"9���խF4��
��ھao��
9��H���B���8jNL.3���$�JL��i��3b�2˖V����'�ɞ���%��ؼ����1�Gך��>Ł��W	Y�7l�m�k:ګ��x^��[�n�_B�������k�#gf�����2S]F��W	io��������\����K���
!DVt�����Vo���Ld�ʕ�����B!D�H|��9��L[[[&�
E�_!��*_%�}�&�;c}vf�|A�X��8��gϞ\��%�!��!�>�x2;�fD1H|���2oy�[���f�ƍ���6B!�����!�Ee�+�X�&����^l�}���L�����Z�(�"�����(�����<uttt����8"R�A}jj�LOO�6������Ī��n�ͬ^���kR�������~���U�׽�u��K/5B!~���纥[#����2��X�lY�5�9�UvAkpX����xV
��Cwww��˗׵jP8����^�GB�LLL�����sL�>|�T�"����/,Uw�qG��B<�|�ͧ5!�X��Q�tCOO�Y�ti��#�8h|&''�����T����;%��B�P0���Җ������~PI���^�H��_��_���B!D?��h�
�2�o춒V�5M|Q��-X�sʉ������b�Z�~���7�������n
ޫB�,\���:D���-��z�
_��U�Vf�<�Aa#��s�7%�s��W��.��|���7���C��֭[͟�ɟ�K!�")yV�X��5���Y�&�I�`��/܃���o ���p�!���|��=�y�yꩧ�Ν;�ѣG+%bQ�i�&s�e��2!�"���BU0�`C����&��^L�J��|y�c���2�L���/!����w��\w�u��<�����G-��E
/<nx�X X�B�q?�����U���L�lV�!����<Cy�hD|p3g�5�9R7V!��P��aQ1Y�P֜#B!�H���c�� ;t�PMo[���� js`�`�f�zŐپqo���9��^c�B������+����3��5������OTrA�$,���W=JA��?�C��!���}��^���$(�B�� wc\�����6���׿�u��c�E��yG�܏���8�a�*�	���?�3����p��>o�.j֖DB!��tD�8/�0�C���������g>c>����7�:kF��+.� 	gRx0�%�-������B!��Mi��ۿ�[���߿?_B��_���D^n⋛��wR3�HFڲ&_=9�aNLv��ΩyA��dB!�cf��LM/3���m��,�W�v����~���*�W�4N.�fpl�?8���̊��f��Aӻ|�!�Y14��]c�&�R5?P=x���
�V��*sa Ⱜ��27�f����k_�a�F!�h�6�ҫg̋�U���a+�
�(�Q���L���g����w���q�!�i<��%�Ta,�O�<��wy]��Y�;*�����/!��X�*�S��7
_e6B��/�ɩr��	!�(?Sӭ3�Ta,��׉St.-wf~!��g�i33U=�OU_a�r_\�̅�&�k��2B!D#��?��U�_q�5�ي������W��!�h�����'z���U�
cy�IV	.+�����J��A����ǌB�(�<k�K���j3xt���pX��r�^�����I���e�J����>n6�>h�:'��%�XB!�lݪ������Zf��R9!�X���������u;�Y�P�òҹd*`B!D�,[:3�j�T�FY�=Q��su;R I�*J�Re��Q!��9q�D*�&�g�����-�\�����c��+V�}�C�����~7�w��ń/4�ڪ��L!�k��Ws���E\UR1�������O��,�����/_ooo��{��޽{ͷ���T�x�������S=xIev��e����W�.B��/���-f����f�ʕ�>��!�}-�����K����:lCmK��GFF��@�V�'>�	�կ~���9r�lذ��g��Sv�FW���+b}vv�����s��s�9�<��SF!D�8��s��ŧ���wh�����h��+o��z`eB�1�|�ӟ6_��2��۷Ϝ�����Vk%f�%��illl���Ca���on�:�-�
=Y�ssmf&�Fp��1�f͚S?�[�μ�o8���B��w�`P��<;���ݔ����p0��	����kCS@�e���$��z��Bd.�@̤Q�?�\��= k� Ӏ�4��n6�|��_`��������ͳ�>��F*�B�����6[�l	�I7�	��/|��ٳǔQQ z06�q?��+�-�+D|qG�܏�H��)��ǵLU��g?k����nA�ݼysp!��?������o�o!̆q�Y��h�81x�)!,+CCCfժU�Z���r�ŞZ�7������?on��V��B��C�ȗ��%#N/�G���x��!Z��
0L��V	d
�rz��G?2��B!��;��|��0Uۣ�H����ߟ{z%�M\���p ��� �<
�k ��2�.fy�@|]w�u檫�
��e��E\`��wq��
�_kɒ�,�Q���<�5�`�U�IB��{f�6P�y�б�uvԡ$ɝ��3F�l�/_n�"*14�(/KvY�L3����!app�<��c殻�
�_ԇr�3���'�5�4m])�0��0"Ĳ��ge%&GY���2��g?�2q�7�;v�r��}�{�����k������r�g�y��~���~�ڵ� ���m������뿎�*8�����G�G�+�����{oh&(�}�{_.�|�W�����~����>f����C�C�t�Mf۶m�\��O<q��Y�����=�kr=��g�@�n�h]פ�brDXVB���Z�tMM�A��y RQP8i
�0
TfX!�B���6Dh�4�Y�z��d�Ȩ�`B�q0������fu��f]XϪ��K$��ŗ-m|���st4^�c��Ն�GGW��\{������O��w�\P+{�͒���-S';��X�UE=�O��Yl��f0qX����9f���X|��~�i�������Dm�������3�g_a���W�?c[&��5��=&}ݣ�Ѝ��_��]�+�W:�����Z͑�W��˅��Xl�/��0x�h<=��Բ؝lo��ٶa�ɂ��x���m&�k�9�Ō�wݍ�����;1�_�=���m<Ven�=��BPgU���=+�g�X���6n�?0����B�d�����[|���U�������К���~��QS]_���b͠t�K!�����B!�(�/!�B������L�Ye&���Ću.i<�lv>|��?�m���L��]>f�X���>3;�nz��ͪ�c��-�4*����2�'��D�/A�y����̉#�9�/�?���>3z�,�m�o���{�����73�K��DÔE|X�䍌��3v���6�ͷ٘*�*��g�7���~a:�f���i���b|b�ya��ya�۪���f������3���};�Մ�C�̺U�������7��<�p'�����3^�$�9�cc����[1dy��:s������|~�`q�����e����� 1��+[��o�����*����&p��1�m6��{��3
\�W�-,?8�6X�y��ݹ=���f��栌-<�9g��d�b����^�����qO�N�(_�2�΋�]�l_�����6��m����L�S����^R,���f��V��>�e^ ���5��;�����Ybv��n.:s����B���m� �n
�kM� �]�e�w��2�ּ��5�C<���]�ep��L��C�CW�!�����F,�{�5�$u�3��[�5Yo�@}��^zu��p��\�!A�KT�  �ev�m��L��(���5����֊������e�{a�%�5��Or���5f��l�5!wVt*���|��wezM,�X��88/����l�d>�),7�EV9�$���o=tl�ٰz0�\o.<cT���u������@dz���!E�KT�zI.�ط�l;�cǹf�T�N��ӕ�u�� �!��Y�_XDjqtdE��kx��;�	by�	��+N��`a%,�|R_��o�oV�kq�(%���������9���Xo���!����/�(_�2LN�$�X�:3�+�'��}��kr���\3K��%�<1���.�˷-��e�� LL�O"�5��̮95���cgY��1�q�g�N|���y�A�f�ԫCy�B4�ė(%'&��6��:Y@96ַ �cz&�N����k�9c'�O�)�eYqa��';>�i�3�9���'g~{��1�6������C���zM�����sq;:޻@���]�Fƿ�؉���&�����=��4>Y_X��N+������12�cam�{�`�Q����t����������BQ�f"�%J	��I!8>-t���&a�40p>�/��5���śݧ-���iҒ��^��J^ ��j���X�VM�,Eiʉ�i�4�RP��*a$%m}�4�_"$��B!
D�K!��@$��B!
D�K!��@$��B!
D�K!��@$��B!
D�K!��@$��B!
D�K!��@J)��,Yb:;;MGGGp������6377gfgg��̌9y򤙞��B!�H���t��Z�Vkp̹��6Hi����m�-[@\(���	3>>�B!D����.�|��@t��555�'N4,Ě.�(����D���PC�q �FGG���B!� <j�����H1�C+V�0ccc��(���&�����O-���900�����$�B�E�	�ő�91�`��󖔦�/,](Ǽ@��Y�&`i
E!��kתU��� �F$ܘ��É�`����+W�6�%eJ�P�0!�B,0� �l }��Z�z�
ơP�EA��+���1#�B�֦H�e�Ѓ��ȑ#�B�
_X��^�����Ǐ!�B�&dN(ZxYpCw~���.�B��Wc-����ՐZ	)�B��=�^RYp� k����F��Or�С�KC�BQN��Fs4ܞ�<��"����QK������_����*MT10�	!���'nhӻ���@4����o^~��ȿs~��F{r_�^)�Z ���ַ���'?�I��#��6��<.Pb��HB!D�I"���� 8>_�������}�u�֚�C�`�"X��/.�q�}�݉�������?6��rKl?/���B!D���3&�?�A���u�]�[���������{¶"�M|��K�����{��M|�4,��Q�Yn�)�B��I��o߾}�����q� ���蓛����	�����BQ>���*��/̀e����*����՛�oX@��~�@��0Hy��59w�������E0y=+�y�AC^�d�tX��&DY�i3y��Z�ł���5l�e�W�Pk5��$7ŠRV��nn�+������a�j�<���Q$����3Es��~�_���Q$�w�.�|	�h�;M��(O<�Dpŝw�i����c9	�?��M|�!�F-�~B!��M��^�s����H33�
!��q�+ ���F�k��*�0!�BDSUCJn� �2��B!�MRF���&~β"�%�BT�*�V�7����$_!�凕�e'�sSG��2'Z��B!D4e��B��I����k�JTRH!�BT\z��������/���z,c>-{oB!��6l�SV�511��\���棯������妛n���Z<��S��K!����H�a�n��.��?�|��b���/�U|�oVOOOݜZ����SX��6�B!D�����H����?rج��Sr_�q�+VD~�B���g�|��k!�⤏�kca!�B4�Wwww���ԧo[#9��/��Z޼�sAP ˗/��=x�)
"�kS!���ƕ�+W���#Gr�Dݱc�j~��D\G�5k֬i�>(�z�!�B�jBHQggg`k&h�z)0
_���@S�B)��B��`�"�;"���W^X
z���a,R�a�Cx�TRU!����c>ƞ���ƕ���V�Z)�"\�.,n^B����!�a��&���O?]����B�\|�ť��e1aXs^�.�^q)|�Er^�[X�����\�B�f@_G'���<�<Ղw{��gKx��6���Ve�����|mc�P�$F�2>�M��B4�!�}֯~�+	���u��`A�('�i�h�,�`�;,]i�<M_�ҰPQ �Nhd{ f��S*	!D��OB��Z�괿1k~��sO�(�a˖-^�Z�l�����Ԗ0��.��4U|��`�B� 9�X���{��8qګQQV裈s%�B�����sH�æM����덨ia�E��h�Gh��h,hYy՚.�\x@��;��rP� �%��̔��qЏ=�装%�ٲn�:�q�F#�	��	�M	��@�Y�a���ׂ�R�/\-!D����}׮]�W^1�z�^�ڜq�F�L��6�΋R�/!�o!fhÆ�U`���Ϛ��$d�&��߶m��Q$����s�y׻�eZb(n��6����%�UMHW�cǎ���"Z�/!�(���A�ꫯQ=��;묳$�DfH|	!%�p��?d�/��� V4�ݻ׈�Aj�W���ŃėbQ�5�Ukya�l���FTR��>�D�B�ėB��m���Kگ����8�Z9��H�j�B�]���3q`���%����Ȯ+B�B�K!r��lrBŅ�~�ڵF4�o�x=!�@�K!��@$��B!
D�K!��@$��B!
D�K!��@$��B!
D�K��r�s��s��I�*���6˖,|�ٹ63=c�������l�1����~�cc�ش_�q�Ϗ�]j���!�he$��(!�m���n���i3B��H|	QB�����C+�b��cz���Q��H|	!�B�ėB�(l��>�SSS�b��d�e˖��9�V|�����wtt?����	����L�B��LOO�C�������]]]f�ʕf͚5A�*�b}��@o�����<V��F|�����f�����F=(ftfrr�!�b�cpp0^�&���0G�1�6m2���F�� B���Kp=hWht�A��=�&��������/
���R���fll,((!�XL �v��mFGG}+�[�n�ٰa��U�����x��qȺ�W�X0��,-M_<LoooP���������|Ǐ
F!L8_|��`�,f &Z��)��+�8D��4nɦ�/
 wV���B�`�w��<(�ef���	/�Ƃ	Qu0�X�L�V��;v,Xؒ��ŗm�YX�j��%���ѣ������ev>�^	B:��*bV�Z��Ř����'.��.܊�QQ��W�:&�!Z��fz>����QT;�9�@�pݸ���h����&&�h%FFF����A|���j4CxY�~Y�Q�B���x5kdIu�:�� �򀕓+������t�ZE�Y�Uǹߡ>y�x�5�}0�B�V iZ����U���2��@�$��Z�湋�8��^xa��a�u=�;8r�e�*H�<99;?q�\|V��YV'������ʋ<ܙB�M7�s�9��@�}���]�`₱'*�h��kS�%�|�#�H�k�w�}��2:��,x9,	U"VQf�L͚�����;��~&^���;�"Oa'D�0�����t�MA6�4<��f�Ν�����Y���=��/�^q�ܮ]�_�����͝w�in��X�B�a�RV!D��;��r$���������~:�w���/������o�������0�Z�{ｉ��&��ė���1���B��4��%%I�%�/ܛa:%7�",�2e�'�V>
�xa9x�}@ޱ�y'�T�UQҊ�"��
_yw���I|	�x!6���I�I
�)��܃eX5&D=he�(Di���8�}��ѪG!D�a�8	Ӟ[��Sv��0�H����eF�B���
�<���X0%D٩�X�=&��K�-E���BTr	��z봁���/Q�0���cn������.�%��8�����w����)D(�րB�IL�\(J�*�h�ȗ=k%|L��͛KG#��
cy�=.Z���_���lٲ%X]�&�B��U�
cy�=�&�H�P�tJ3!�h�=���K/��:����U�
;1�������Y|i�2!D+A���;̫������A��_�>�^wB4��R��Z�0��T��4j�B������z�js���`+�(�X[�re\����� �8�Z���Fnw����}�De�B�*li�}��`�}���` �`���]]]��mm�_)&D=�e_�[F������A��~��f��݉�388��;yo�!�e ��L���a�����o|��4G��.L~�r��*���b�/L��r�)D!�%�B�����d?�[o���<AkD���0�"�%���������on�Za����?�4B!Dˀ'�����;�>���b�q��
_"����'w')�MFe�G|��g?k�_GP!e�B!Z�P=c���{��md_�zq�$>���8w�("�2���&�9e�B�C,T��:-�|B��W��'�<*��R�rX����L�@ j���Bn�M�6�v~B$��(�+�#�J��oƕg����!˚{{{M� �0G
!�y�5���Jq��!�hhh(ر�hƵ�&8.�6g�e�Z\Sq^B!�䢋.�č����
��\0��J�-	m�+�w�R�P������RV`��ʱ!�B��v���`�$)(Ҁ��Г��D��_�JȬ�l[o��B!Z�PX��H�q�����Ct�1�4mI ��o��	d��B��� ��Bd0� ����0����X�o�d��/K�`d�8`٢(T��F!�����56)�v�2�>��BQN�>��&�=�
1�.�F�LM_��")�[8 ��@�ɵ(�b��mf͚5�����/��c�N�(���?0�0�7�%�""�����h��4�UWbV��I̚�lL6�&��Uc65����X�/�S@�T�a`�c������2��GUwW�S՟�k{C�tO�]����<�@4�}��=��L7}f�OyC����cM�jH�4� @����0Y�   ���  "�
Fs���Ҙ[2.�C����q�&  �_(�֭[�o}��Ps�ԩ���g5���^�ܿ�U�� o�/  ��   BD�  �   D�/  ��   BD�  �   D�/  ��   BD�B��l^bv���cV�9h  ��
Fk���1K��  ��  "�  @�_   !"|  ����Iܺ5m��<x�:tȹ�v��Q�C����o�K  ޔ3tss�2GP�
_
Y-[�tn͛77%%%�ј^�������z�w�^���PI+SҲ����lj?:n�ر#���c ;)c(k�h��4k����)�8p�����s��s!X��˷i�ƴj��	`�(��{tk۶�����cv����'�W�vnA����
�̔�5Z�n��l�Gt?��=�����ݻ�z.��/%ϲ�2'D��}AuS���-X:  ��BM�v�<x2q?�Y���z�I��/_ZZ����J�;w�tn  �8)(u��!�b>���sU�����]�	=|�	w��ѩz�w
a۶mt��cժU·ȯ���@q۸qcA�k�Ba�:�,$��N�:9���yj�����<�$� �E���0���C"�W^y� @.֬Yc`U��yZAS�GE��۷{�Z�҄�0�W��U ۲e0  .���P��� ��ل���^.u��n�J�0  JÌQ/���B�X��/��BOv�KC��G�JH  �,�*Ĩ��ѶLӝ_Z}����R�� @rh�O�h�OŞL�_*�e��w��]�?_�g�.���z���D
  �A�/�S�[n1���9=�2�n�=���;wn��i�S���{_��m�Q�KC����K��/}�K楗^2&L��<��R�-�`��}M̂u��c�Պ-�NO ?nU�ܮ��t���h��N3~�x'Kd�!Pu[H�L���R�����c����_�٦M��'۟ �@S�rY�7q�D���g�L�L!/ն���/U��l��������#F��P���g�1 �?���)o��m'���~�A���Ӎ����<�$_ �˝�d+�W#�/  �M�+�Ͳ��aG=��=F_^WD���  2��\���i����f�U�M_ @~l���9m���L	  ��ù<�s,|i|�	  $�9�h�l oqh�*o����C��6�  ��C�
�ɪ����W (.}��1]�t	��/X��l۶� ���rU�R{_ھGKڊ�@q�š �iS�Waq��ꗭ���7ֶ9�(��#| {:�y!��t�����K�{�!m�������	�  �_]]���}���r���z��gT^^��~[�n5={�4aٵk�  񧀣y�~��k�gMM�	�Ba���/���V�R�\�~�9��S�z,u����A�H�L�D����Mס�>����b�y�f3g���V @.T��С����\�Ҝ|��ybTi�V9�4���H������2��������7�w\^��%x��|���4o�9��ܻ�):`� 8��Lmڴ�4��O��S��G��`�i�2��*�i�v�LԔB�� @�h��=Q7xWU?�<�P�דв�-[��(3� �dR��<��;F�4
��~�*c��/ѓ�������) ��Ҽn��۷o�c+p)�x��Z�ғ���v��1�BѤ/)  ���ݻ����܊�����/ѓS �F�{�5˵  �'0���
Ƞ�߫����
5|�*P�UiP!,�E/��.�  '�|UUU9,�9��3�K�B��ѵ�×K�K�m۶έ�TY��Ì  7w�M᫴��`�Εa4��k����EѓWjTE���(�i5�n�.  А�`�)�)k�~G�4��Х!�|�DG�\n�N7u�ׄ|�0m�?�*�V����W���K�U  P���L��j�5�@�\���+U�(��8V����U,ċ�&N��c�B ���>n'
օ/ė�֬Yk  @z�/  ��   BD�  �   D�/  ��   BD�  �   D�/  ��   BD�  �   D�/  �� ���כ����~�Ν;ͪU�́<ݿiӦf����ӿ����M�^�LIII��7kƩ���P�v���܂����y�⩾��}�ѦI�&i�ӲeKӡC�A�������l߾�,_�� ~jkkͺu��T������ t�1�8C��7o6��M�6�V�Z����þޢEӱcǌU1 �`]I��G|���Ӫ���C���_bj�9��w�1���3(<��O<�D���o;!�x�r���:V𪨨 x!g�/�2;v0�F�r���6-2�vl��g�(�4�;9��g�&|H�G�e�L���C�2+V�0�6m۶u.�^�� Bкuks�I'��ӧ��ċ&�/[�̌;�Y�
�ú𥫉�͛;e]]-�M�������X�"ą*&Æ3���A��޽�Y�:r�H*_	���f7o�T�T�p��޽{z�dM�҄F]j\�ϛZ/О={>����~B��XO7n4K�,1�2���6m�8��K��T�Q�P�7�E�4~�������Ц�ҩ��� [i��UZI��Q�j׮��ѣ�A<hDM&T���g����:g��&ʍE�T�k߾}A;�g�g*ժ��R* �F�#F�0S�N5;v�0�����)�`�n��)�@Sȟ����� ��*�Hҧ�cP�LՓE���;X@.t�x��';-(��?�xh��1c�!,�GY@��rY�F!̭�m۶��Pd��KOT/D>e??��ʜ�B���Mt��
�̙39FŐ��̚5ˌ=:�<r�@��d#4��������^ �a/�nZ�PSS���u:u�dN;�4Ř*���B~�o���0W�*|���֭[=���WT�Y=��`� �a@�0���Q�qG���M�%|i~W��5`���C�?�G:����D+  @����e�;}�:���aÆ��e�� �i�-��9W�&�kH��o���k�������m�Z�a�\��  ;��e��k��戍ҽZ�p���㏝�n����
>������4F�������ͤI�̄	�>��2A�  @2ht���>�����}��殻�2�Ǐ��x��Ǚ��h��ثn^h8��7���~�h�}9Ԑ�Q}�����2����S:���})~6{��\�W���[��G��P�G}���?�������a+�_�뮻  ;U���=�ؓ��6��qװ�Jx��� ����ɭ�_zn��<,|�m��]�K�0��H  `�V�0��j���ؐ��  �/uT��1*�F �6|rCo  >۳�F����������\��  ��sy����2����  @fq8��z���  �(��=�l]�(��\  ��ù<�s,|i|��I�t�  ��Ws�MVm_�K  �W�
L�KG�s������a���Js�	Ï�zi�zӪY~Wyu�����G~�Ly��w b��s�
=�;�@�]��R����~�\��r���ڷ/3#G�<��u��};6���;w�0�;9��ӧ��3 v4��b���5h� ��3{�l_�Ow\,|)�)�zz�~��ƍ��8��~���ы�qb ��}���n9��+������9��ԓO���:������Ǝ��{��y_�߳gOʯ:)K/H���qO<���[sz�U�V9����^+m��Y $Cǎ�M�6)����0����L��M�K���FYY���������r
��6���öm�L׮]3�WE�t��_�v�2m۶���Q�z����~,/�KոtI  ċr����ɓ͂���\���d_;v�H�w��/�Q"�D%׫��:���:�Y[[k  @rx)�4t�W��x��kzS�y������2o�Ro�c��Ȥb  �EŞ�۷��;z��������M�$***"� SÍ�^ @�-^�Pg��gcGt�Uzw�̌��4�ȭ�EIY#ۢ�P���G���#y�񫫫�!���[�fu�Q�0FY��yqٲ���<+zҭv��L���&�) �$��7x�Z �dS�E�e��W�j��n^���O� ���xj9(� �� �s�V?�5��F?m�B�|Q�����Y��K!�E��F� (.:�+��Ӿ}��F�4�\�6��EG��@���
��@/�^p6���4��ѦE��CNSޜll�s⹟9?��?��O�F9C�@U0�S�y��7��.zr)�D�\��*�&Ʃ4��� �_\/�V9�J �[YY�@GV
M�0-HC0���
>������k%L�.M�W��gd-���R2�M��4AN!L�L��4�K�K7}�^\ 	��7[�V������%�M ����؝�g���t����?���ѷt1�ܦ��U�"|��¨��NZӋ� ��*��EP����˅�Z�f����h  �h܁^��n�P���Ԫ�՘^ %N  ��(d�9`u�  H��0t�P3r�H�ߧ��ĉ��Ͼ32�b���C�n/�w�^�g�c��f%i��hx,�s��[�����`�v�ښnݺ��>Z� �I�k�ڵ������k����L�h���7������]g�w�f?�/ @,����Y�X���&���x"| b�	`M�����i������:H���"| bM��JK��ɶ�y�	 �_�BISc�{ߔ�u�  f_�Be�CfǪ���I���UTT��n�鰯͛7�<��)�?l�0s�UW��_|Ѽ��)��y�s�9簯���%KR�	fРA�}�'?��3���N{���ޚ��o��?��a_[�h�y��R�����k�9�k������_�j  ���4Ǥax�L{�5o����k+�t��Z��k�?��4�Z�mx�LC6�p����>� ��   D�/  ��   BD�  �   D�/  ��   BD�  �   Dև/u�vo�*�]�\���i����������/������}�ߏ��?q�D_?����	����M�^��`4�%CyC��X��������%%%έ�8ۃ���;���۷� �_�i�$��u����e�����:v6���f}�7
U �"|)li�4�0�򩸡L/Z�v����ι�W0���ކb�UUUf���@~�/�5t˴wl��+��E5��ٓ�s�4|�/++˸�:ٴm�ֹ)��ر�  ��|�b��O&��馊��F�!,��UZZ�����z֪U+�E	j�  ���V;vL9�)*��VSS��z�R�JOX�1(
tnEm۶m�N�  �Q�GY H�2�:ur���yj�RR,///xMG᫲��lݺ�U������9a���S�ט�  W���?��4|�m�o�nv����{B_
\�-���� f���>y��P=X�ak @���?�x	`��/7��\��luu5C�  $�&�G�\���&��աCO�:��qY��h">  H�絘/J*6�أ1�F�ODZy����,T�  @2(���~Q�(�*`Z�N��+[
�v�w��8�k֬�z?��lٲ��.�6m2s����}�� ���Ʃ���Y��wۡGy�s�ܴ�S�+��J7�h���b�g���R�������^z�L�0�S�0���*H?KB�+V:7  �й_#[^�#r�䀛n���y�f���Y��9i�y*��/�4������h� �A'_-�/�)%:5�h���rY���C��?#g
g����k`�K/U�l�D�P�� �xӱ�n�n�r�
SL�w��>�h��Vzn;w�<�끅/[&٧��$�\�f  ;��KsF�������!CL���<�s�,j����D6���  �����aV�n��7iO����v�b��О��7uN���Gt!�,!�:��= �SEa���?n��G�=�=����� <amW��_�w+�_���Z>0�`�-t�P�<M�U��j�)�~D(�r=G�����L	�B�RjkkS��3���m۶5 �8��S=���v5!� ���5���L��zK �)�9�h�l#.4�7n�8O��>}�3<X���o�V�hr����ߙg��y����VYI��Q��c`�KsClzl<�
�J���K/�t_m��m۶�S?��u�'|�K.���h��ń� 賑�i&���P��*�ؼ��  -u��S��e:)5m�|$���=���a�hOR�^H�q4�𥃱�]g�mv	 �����)|�<�)�m�;Q�P{��H+��@��󹭻�����R����?�-4!�	���_��nO����wʀ��+x��w��FZ�
�O�%|�2O�υ�rF�����yߵk��@UVVf���~���~����޽� q����{��}5��ϭ��Վ���X�`�A�:����x�Z�� |�@��ߝkƏ����ϟ���z^�Vc���:xg��֛x�ҥ�G��1�,Y����� ��^�N�̠A���O��Y��KD[�f?��G�U��c�J{��?DC+{;t����֭sFr�~��;�8��90[�,�j��78TƊ����������<���y=�N]�v�x=����֭�9�쳳�OUM�W���ձcGSSS��J_<:�1� J�S��h�]w�e|���
1
p�N��:GfZ�x��/�'���X��:+���x�B����L�(T�gGW��*H]��@�[�&,�=�y����tL;vl^-�:w���3Ԥ:��×�ڤ��.�j��G�s�(���l߾���
��mzT�W�>��}��t�T��l��B	_�'��G��
AW���B ��Т��欆M�K��������4�_����C�|�aO/) �l��?�4���:I�LGY��<�P�Pn �F����qW�W�)��R�ٿ���MY�z���Y��׿��s��)��ڰ�7�����4�x˖-(F:�kN��]�W�K��Ϝ��� �4�tXZZ�*)���xG����o|=�{S�L1�3�������s��N�<�̘1��J��x�oX��͍�z��F�(v����r
>A}�7TÜ~�<�O��?z�zaڵkW�S��v5��j  �M������F��=����5����,|��b��t5�[./��h
r
t�.  А2�n��)k(��-�(��gd���E��˥_H��nZ�nm���e�z�tS��MIViS7�|zu  �⠊�n�n��MY�ݣ���&�>�n�(+�WCJ�4B�F%�]w���j~��n�|_F����p�X�_�_vo�䊤����n����&s�������b���� H�b�@�J����jiiK+m�U/��������I C�  �   D�/  ���Ć���٬]��٢&-�]�r���лw�P��J�����+=�w���l/�`zx����3�8[� ��H����}6m��s�[n����O�t�\�YB|�9��̤I�_��_   !"|  ���  "�`9m�M7y��֭[��[n���6 �A�,�-e���=�W�"��@$�   D�/  ��   BD�  �   D�/�_I+Ӵ��*�����شykc���v  \�/�^�.�r��p˪)��ߪ�	�y���g�d���mۚ_���;n�8gst$ӯ~�+ӦMO��{fÆ�}
�z���,�F'��;w�F-[��t?�8O����^hڴ���]�v�gϞ&n���̪U�
��;�X� ���*� ��ر�9�3L�lڴ)��/u让�qn�v�r�V9p��s+))1͚5s��J�z���ʸ� |j�����Y��ۚի�s�Mt^;����ҏ�������Pڒmǎ�{������YSLTe�H^��흼ѢE��=�5�k�ƍfݺuf��;�dz��v��T�*++�4� �:��t��}кukO�ݷo�)Vg�}Nڹq���ӟ�hW��$���K���$0��.��5k֘����
�*�t���t������H×��[�z�Y�lY�W"J�z!uSl���[�nTÊ��/�lJJ���7o����/��RN�htA�]���g?�t_��K��n�� 𯶶�,Y�$�E(�+:����G9���s�,|��?���~֜9s�����Ý�I$�G-	�q>��C �MYZ�x�3�J�T�\�b�S�4h��ׯ��z��/���;	�P/Dc
vo���9��cM�>}  (.۷ow
2A��S[�h�3���O�U5|)����{�Xk�4Of���D��C�2	 E��n�9t�C�(�b�}Ai��y�B�+�e�3e�3j�(�#n��/�!%P%�0�\��	}� $��S�4{��M�w�4J�撾��si���?��5w�\'w�Ess�M�fN=�TSZZ�����/%а��K�ZM2d�  �I�#�^.��3g�1c�dm�J�Z�|y(C��hE�zuh�('j-�����}u�Ö2ɥ���V�����^i�ɞ={���9�����N;-c�2��n6���~������=`I���͚YӺ���k��qx��7�����):���?�}?R+�h�U:J��Ǐ��q^x��ܘ�z�}������ܥk�	��7�WT��g�^i�~�E�����饗z����:*(`��^`=z�p�cM%��0�U �(|i�Z�~��Y�f��}�z��:D�k7� d7|����m4�������3�v�	'�#����o�}�Y��j&*:-]��鶐J��KMȼ���o���1�|�M��k��	&�W��  F�IDATxZ��G��T0 ���ڧ�`̖�ß�;wz�7潀b�B�zz���������S��_|���6�I���r:H`�K�~V7*%�2Q8���_Z���V1@ش�����mO��6�x���7�p
9�P/0�4}�+��bã�:ꈿ,|UUUY{�g�_�� @<id �6V^蹅�������� ���P�
*��h�b�iQ��/m�c3۟  ���s��)��q�������� HO�,u�m���͌'O~ݴh�z�㕫V���5�&�v�2���״��jsʹF�STY�۪��j��B�s-|���e>�L� �E�86n4ݺv="�͞5�ĉ�G����PV��ڢ_�gI�	_zS�f��,���K��n��}Vts�Z�婞c �KW$j㐩�}�؆q�ϓ׆��OI6���3mqb�1��6n��0�'^��Ki��8����K-�m�eGą:u�z뭞�F��gL.����O�S�n�:S,4�r�HF4��%�ù<�C���v��Y����	  DKY�v��3,|u�����g:t0H��]��t��J��o۵��?p�5�*M�b W���㻭�����LII�_,|u����F�a�?�����SG9�i5t��AS��ͼv��'��V����0}��'  \͛7w�)ڵ�F�;wN���ҨJm6=�����l�e�ӦM�t_5�Cr͘1���]���B�=�_zn��T]�~F|�A����֚�.�,��*.��=�{�6@\h9�C=��;ع!��q�p={�tF��������l��F:�RENÎ��F�o߾fٲeYC����W^1a�\��ݻ  z�ӧ�Y�t������`w:8p`ڿ4|i��<SuJK�o��6s�����X�x�p7d��}r  �����oV�^�i�׿��?~|^���8�Z��'_�.]��}���T�R��L�a�ժ⥕p   9Z�ha�;�83gΜ���T� ��4lذ��	�5�ȑ#�[o�i�aM���b  �xR�E�V�\��PL�۫�PV�|���J�(6��� =�ƅ�8��6%^�M�X{�}�Q\�=�X����͛#y|M��իW����)����t�If��١0�"O9�Xt�R��w��龧�v�Y�f�A2i~,��i[e��3g�-[���ؚw6h� O�uGJM@=z��5kV(��*p�╭�  �ALE����r1�j�СC��^���z^�;�yQ�ܒE}?4�+U[�bԭ[7'�f3`� s�9�d��ʺ^{O��^� ���Ç;�7���y�6mژN8�i��G��K4��Ot��.Z����!�Y_c��yw^��덪�i6����  �i��ђ%K�V������ti�W.E�HK�+�
�
�����rBU�~��9�>^H�x�'5����^+�l5�/4���|�rg.d�s����t�g!T��K����n��lܸ�Y*� ��D�@���Ի���T:���7��t��۷$�=��c �F���4:VUU�ܔ7�=�5LUUK#j����S�Q���WC��!/w�Kc�����������XU�R�4����_?��m[�߮�n߇��/[G�> �*mܦ���<fe�TR��:]'V'-��/�T�inj �!����"X�   ����KB���/��% @~t�V#ոٹs��߂�/�$   �B���o�aG  ��   BD�  �   D�/ @��h��,^��`���N}����'�  �Z�li�~�q�/�:��:�(�x"| b)��u�cMӒ��7wλ�6��4���4��~�/F��C���� @P��^Yi�1bD�����8��¿���U�V��\�~/�_8��M� 6S �޽��Iee����g�l_   !"|  ���  "�  @�_@�h���u��a����X��}S\���047n4 
o�ҏ́��mxA�d���N��С�����ڒ%K�K/����4\p�a_�:u��={v���~��椓N:�k�<�Y�jU���_0}��9�k���V������6m�|��;v�{�7�}۶mk����þ�|�r��sϥ�߾}��?��þ6c�3}�tSH���@2��)//��v��Ɍ3氯�n��̚5+�����w������ʕ+S���c�9��s��M��X��c�=�k
G
U��v�i���m۶�S�۷?��kӦMKy����߾}�Y�t��T�_j�WRR�ܚ6m�|MsY4���:�q�  ��6)W��MYC7k(g(oz+k~�V�Z9{u���L���۷���f�޽E��* DA����4m���+W:�X�?�h��ǌ���O�;N~�u�i[&U�5�mՐ���\9���� ���×>��ڵs^�Z}��O7%�]�v9��l s����ѣ����U������}m�y�iQv��Aƽ뮻�����6��x�7����{[�h��4}A!LyC��Ud� �2z4�5�+%ѕ�^�<�(;w�4  ����UVVV����)|����T��$|���SA\=�!L	���ƚR5  �
;
]W:��*�Z裢���/j�P!�]�(��EQ Ӝ0  PT���oe� �OC��^瞇��>�¢E6��$9  �1c���Ń;j����)�E�m;vt��x	`������K=�&��39 �wg�2��[�
3x�4���X6��/��^.0%�-[�0 ��ҹ>�ը��iR�3	������C�
`   Y�AAŞ���F�2�����0[
=��~��>�(�V$.M�s[Q �N�y~��þ��BF�5����D[	m޼����_�>��_�u3gΜþ�ia͓O>y���LE�m�ܷnݚ��k׮=���W�6 £���其&�a>V�X�qxQE��Ǵ�_sͶ�S��]w]Ώ��k�9:����D�8:�҈�N��w��|�?����6�NeѢEƏt{P��]3�<w���@�����_�tC��̙3͂���L���?�rI��K������?����~��4i��0a���R�SP�� @�����5�|������{�ǌ?>k�L�0�� 䧱���g̘��q����"| �6Q�%s��=G����X`�K�޼l�wsV> oZah+=�P�W��ق�pH�  �T]�y��tY(�g���]���L� ���l\YZbJ��u\��y�n��þ�o_�R�=k(j��"��_�?? �KH��-)ij��~�o����e�k�Z�6m��܀��wc!��x~z`	���^��7��p�駛Q�NI�w{�W������e}ǘ&%G�4��;~c  *q8��z���v����  d�$�+U�,|iH���ˮ�   �H�7�6|�� �x�ù<�s,|���[�n�6  �[�婞c`�����f
�   �l?�+�Z���\[��!�m�  �=ntS?-����/=�Ҟ��
U��� @����9�X�(]/�@'��i۶m����i��k��~��7��=/  ������,Y���c�X���}U�J�����]��h�1۪G���o}˄A��m�  H�f���g��o����Ԙ �ڵ+m[�@×^%�Ls����򗿘k��6���x��I�
zi3 @b�ر�������?o��⊼VJ*sd�~���t�శ��yA�M�S��:ujޏ�%x���b  ��q��^�gΜY���D�'S3��×|�����DI�C%F:�@~�=�<䈯�5�6MM~m�v*5����G:�j��D#[*�D�ٶ�6��h�
<|�&�)�����( �� ���>��;VM3�3�t�iߥ�iQ������d��ʶm�Leeed������5��%�rы�rP?V8 �l���u�V�!��_*�(�yZ�M��Ӿ}�P��$x P4�`͚�s4§��ujS��K4�� S�C/C�  ���N�[��q�4�����/QBܲeK`/�&����z$����i��<x�4iZ����}�>��G�g�6� ���RZh�cfiii�>�ߥiM�y"	_�(��P��9�q;�+tپ�7���ߞ���5� @\)�bQ;��h�!LaKY#���˝��C�iukѢ���U�R����S @c�
L*�(ch�ME��"5�L4�BLg�<|��n����>
d�,�?�OK�eslo�9�s���G��o��ٴi����ի�9��"{�ٳg��˗x���N�ps�n
b�����7�5
]ܱ&|5�V���޽{�q��E�����#|H�.]����:+��_�~=�+O
W���K+�  @R�   BD�  �   D�/ �/���RN�n{��ij�k�][���o9�Ү]��$�/ �/.tn rC�  �   D�/  ��   BD�  �   D�/  ��   BD��Pee�ٹs�a_;v������3����/�`,X`�������-[�#F��\�,Yb�nݚ�������q8`�{�þֶmی� ~u������N�%%%��/���/���Y�f����{S��)��b
e�������G|}����M�6��/��1�Ν����!k�u���3`� �?c�����H��(ȝs�9&_����M�n���?�>}� (���j�aÆO�ܢE3h� ���=�8��y������?�4i�����޽{S�����Ng�ʕ�!|  ���  "�  @�_	�I�w�ygڿoڴiA�ꫯ6W]uUڿoժ�����/~�r��P��W���9t�P����X��Eo.���ӛ=�Ӻu��C�T�؄q|u�b�RA�aQ���Bo��
_���A't���՘^����;+�D��^   �,�n�h֬Y�� �?R�p���w!X��˫���!*��͛;7](x�_ˮ]��@  А
:�X*7�{���D�K-Ft˧�i�R�*++sBT>���dZ[[[�t
  �K����	]�ΑS�L��]�vfǎ���.�I�r_U�
M���߸K<  (��۷�\��JÔ��
t555�>��/� ���Nz����o۶�	�  U��(�4��;|�o��T��
5|�I*x��A6�ԋ�m$�4��l��b��w�� H��V�#��:t����4�܋�*]a/�[i���Z�����7�a���'�3��e˖��' (�뮻�t����?7�_Vb��R�M��PW�˥ �0ZR  ���<�reso0zԁ!�P�q���旆<��h\  $��ykbԔy���2������폑N!�>�T��*A����g  @2(Gh����S�ȴ哊=Z�N���]u��^���;��P��)��5k�d���q�H @2hU������g�b�\h>��>���f޼yi李O-�KW�	4|�����P;�\�r]~��楗^2&L�TAӄn�(��c ��t��e�1�iH?��O�o�[3~����z*>i�y*��/?��*x=����O_��� ��S�'��KO<���I�Rq��L��*����h#�Uw�| �xS������G5X��V����_.U3  `U�l-�F����C��_  ė��6�ks�_㕑��� �n,۟_X��*�?�Ь_��lܸ����VjWϒ�ݻ���:�{�YW� �F���,Yb�/_n֭[���1V K�VQQaz��i���c�9�#�=�����}��uS�ll~AR�Z�x��<y��5k��#�WJ�}��5g�q�;v�s�  ����9��8;�|_��t�{�qǙq�ƙQ�F9�H-{����X�mC�"�VBW_o���yꩧ��ի�����#ѕ��$��eR��}��`�w�^�b�
�
��6cƌ1�^z��ݻ��b����=��s���������n�8���c����qV��t��	Z�Y��z��w���W]|��梋.��{;�K�7�k�E�9V�Z��y#(p�`�i,�O7$T��}5����:ȼ��[fʔ)泟���ꪫ88 (J:.���k桇r&X븩�F�e�1ֽ�mX�R�qV��{�	s:ƞw�y��� ��ވ6�A�e�m}�x��JL����O�W]����t��4i��6m���̉'�h �Xh���n.\�i�O#�9��t��<\�t�a��~���s��񐪭U`�K%T��W��gI����s����o|�	K*,d�Ꙛ�*����?5�]v���+�rh@qY�`���㏝�����+�b7��X���}���ַ���#F�b�sy��_��ؼ
a�×V����?6=z�0o���ׯ���q�ĉo.���I�����O:�O���6 H6M�8����W��g@Ã�<�Bӱ���ܩ��1�?���_o�<�LS�l?���,|i ��n��$زe��я~dN=�Ts�w:����7��_�hW�W�f�������_w>�l�� 	�v�Zs�:�H�^����p�
۶ms��:��u�Y�X��c�4'-RK%���m�7kR×��~����|�3����ߝ��n�ə} �~BP��ƴ) $�*�������m�ݖӾ��Ѕnǎ� �����9�6�+��l�b(]�t½^/�龛6mJY��F��/�I�{�N��<x��կ~唧�������&C*�i��g�q�W ĝ�S��r�s��ܫ3fD�<�4�LA�?��?�o�[�
W��f�~��x.��OaI��t;��jB'/�K�T4a��J��_~�)�k5������Ѓ�KW�ꌯ �����Ԑ,^Ux���� t\�ի�3���� ����b'M��D�;�ÙV���4���*~����x.40�T�@×^��2u�Ձg�ʕyO�dD/�B�'p���Ϗ<�3�K���ATw�(i^�Zy�����|�;ɡPYYY��iL��B��׼l}��z��s�;�w����.j�^^���AG�W�k�E��7�,�	�:�x��ת��O?=�ϝ�o�'�]��]�7Y�S����	��O2��q�/�'Ӌg
^*��٩�]a�AHG�������!Q ��9��a��?���Ta����>���f���E���3^�:�u�~���V�օb�a��×�di���s���͛��F7p���F�TE���O<a~� �S5¢y��-��p��h��W_u.t���ȝ:u�<+�d+􄲽������$Ҡ�;�'��H��t�i�9��{�=c�����ܹΞ�Gu���P�2d��+QC{6���s�>��9���M1��QqE4ʅ
�zل�����DQU)2��+QЛM=f��Q���F:0hr���!! ą;wYMTmUhHU9]�j$DSO�j����:�h�W����e�-���Q=��T�R)2�+�T����s�u���N�jl���J�
��/ q�ڼ����f�~��c[��K�Q�0���2���W��/Q R�M�����`������K�.N��y��Y����ЭI�j�ѳgO ��E��i����m���V
�:��\P������U��Z�r��\�D)�zR�ZI��KָY�p�3A4��f:0�$��L�rTO��j�Z�_��G5.ׅy1�������jQh*(iUc.E�H�/�VA�
V�d�ԩjW���Q�ו�9���Y��l�n�n����GmF�a�@N�i&��tEX���I�^�,���ą~M�N�|�|�r�,����M��ĝ�����/Ĵ'�.��7r�Y��	�~]Y���7�J�I]͘�«x�{�v�� f3�D�n�:S�4�ѭTIb�~��p'دY��ā;���'�t���RSӞNU�Q%�o�GA���^0E�\
a���͝���D����{��àA/�n��t{wk�;��+:�o�G/�p��3����������t�VY��q/#u�N�0Y�L'^=�Lϭ��;�$�����u�Ҹ���}�����tr�4���sJ��s����.���?k1��Gq�/	������oI�@M}��R�Ye�J�0��s�f7orw+�WC�eU�����>w�8�� _lJ�6���L6��$5?���D-K�ո��/>�w�uWl���袋̅^�韵cE�}Y���g��ꪬ?K�[�詨��:��4�n��˞�n�Hj%�P�Ģ�n]��wn
w'��æ�P!R)��@\��˶���g{	_V#|Ř{u�}�a%��k�N�aU @<�"?H��@s�a/�W��.�
���T�92a�x�ͨQ���\�����ƽ���r���b<��I<�MH�k׮���C4aW�]l�������ۜ��$��l^T�Jf!�3/�6l���ދ�s��}�خ&Ν;؋�c��h��;�Y-'>��c+w�Z���M����>gN>�䜾W+sl��{�7-�6�IW=z�0I�;����;�۹�YYۍ�s��bƌ��VO�I�&[�m5�w�n�⣡��L</wn�����6��4F����_17l�0�裏:=K�:�,s��[�rB��9ûCE����˼�B��O�N9�g(O[��Jjv�E9s��V|���9r�y����?n���Z��|��������j1���L8���l����}s5�>w��{����c*,���~����ի�s�s����6����/�Fn5��3�4�'	��!�0�д���[ou�m�(�8�хq��؍� �{��e|�ĉNwkۨr���Zc�3���a�b�|ia�ܹs��/z��A �������φ�1@�J���>�<��c�^�ҳ� �� ��$���[�i��[9s�L�c�+×��䗾�%��@C����p&�kd[h�LmT���K�q{�6(�	���:sl�}�]�Ҧ�G헫M�w�s������0��y��W���˝�-[K�L� ����iRh�lR��K���������eC%P�z>z._���⡸?I	������7�w��]���jX�J��u5�=�_�'�+�{2���ˏ��T��q����駟~��4d索���"v5���+���4�C��D���.�t�������ߛ��:� _	ҿs��W�?��Of۶m���"�m>��Y�Ksо��o'r��0�̈́��?�����lT������t��5k�|����ܡC��/���A�J��.���nH���+�����*T��?�{��aGؤ�+_�J׿�˿��n��i���VC�M�K�iU����W.pc��@�]w�3�8m�4'�i�"���&��˱�矮Ȑ;��&��R�(��U�o��f'�mܸ�y=�j����]�Z�n�r�-V�Bf�������=s�=�8�-[�8��G뀠+1=����}s�'������ݼ��)���׿vB؊+�[A_�jn�F4S��؝:u2��WB)���?���֭�y�ᇝ
�&[�<^���v逬�S��۷�A�_���o�~��_�����tFt�����Pr"��]�ti��	�>�n`��#|%�>����upX�v�3K���7�)t�+�X�s���kL6t-�lü���x�Η_~ٹ�u���m��Х�KQPeM�
W^y���d��,�?�W<x�����SO=�&wx�m=����+^�-\ܫ_�-�����NK	��a�cj��cԨQ桇2o���3<�I�Z�rn^W+p�ت~�
^j��Y[�i5{ee�A�Y�T�ч��S�N�t�d�7�ޜ�P��+²��x饗:]����5�6mr>�z}��Z7���juk�z�a@?|�p�k=s���{���V�k8Pm�}�Y3e��BW7W�c�^���Ycݛ{�Յ�6��=�
O��^c7o�������7����90_V�/���2P���ՁK/��*1��p��L��B����O{�̟?�錯7V&��i��aÜ��p�`Q��m�5c�$���׿�L��1vΜ9�qVs�7/nLN�c��V�4[v+I���)od�i\�U�B7U&��H����s��&W�T�ѐ�^BXfzݎ=�X�&
^�֭s�M�*Mo.]��e�:�hU��U��@�_�鼤�B�DÐ:�*���eu����l�=h ����q��KKK�C~r٧Ho8��
Y���������l����}�>}���G 6a�1w:ak.¥
��-�7��?[E���×*'z�	EWf��PGW@�`#��Dy#Ȗn�P�O�5|)x�/J��>������`@�0�6b�#�@@�.�AyCALy�˅sh�+��Ր�,鱵�4'T�`#*_�]��˥�S�Q��v�-|E�\zA46�qY .�l1���"x�����F�B���)xb��K�:+��ѪJM��wy(�a#�l���-xi�y�[�����>H�wqӂ?�;O'�O��h�[:Z���o~3矯&v�6G-2�/Ѿ�
`T;�F��(]x�\���������Κ7�{�
R	<|)�x�P��_��tҤIf	Y{P頡�	��*_�������E,l�����fmذ���|��_u�{��n:z~���N����/5z�X��8u�Tߏ᷷�ʁ�&��Z�`�y������_o���g�N�8�x㍇}�W�^��`+�h�=|=�������?�w���m����?����}M{�ƙ���y��b/��ᕛ�R�@×�Y�����j�禹�X'�����~vR�`�$�xTw��sr�nmg:�4����M��C���7o,��!��Vd��fh̩���`)&��&6�=/w�����B���t��+�V�/؊���\�T�J�7�����K�����V%4Z�E��!ꕞ_h���+�f\��rT�`+�l�,�y#�gl����SՋ�[��#lǼ�{�����!Gج��,ǼA��U/،���P×��m�.%���>.���i5�Q��~�ŋ�͛7����Ç;����lF�2�w���h��3Έ�cő��6WcS���b�4�'75u{����}EEEA���o�m�Ν���v�J���!�a���SO=�l1�Θ1c
V�x�'Ү��c�_�R����U,�O�7kF�����E �v�	����Ѫ�[�h�`���o�nV�^��gd�q]I\���+�6M[�l���:���6b_�m1t�aGXLU�T]��D�7����v�Z�ߟ�3ZSSS��W������z��i�B�!�\c�P×J�����ﯦ��s�����
���
,����˾~F��4�{�ɗv��d����_��1
��Î���K�Gjkk���	��w����vA��Y��W��|:V�y��:��E��sM��%w����Z��3��*�駟��qr餯"�}�;v��Lx9r�_���%�\bN;�?}�t�R���tl�_��7t��ӧ�9��3S�}!�]��)�"h"�G}d��އ�~�5'Y� )����t�^��UF��y�s�-���6lp�����=V��t��ۯ_�@'c2Ĺ�3g�������/]�j�nܸq�?�&梨�F?�:�L�u%{�i�&s��7��'��X�v����R	<|i�N�U
_����Y�lYޏ�%|)!g�D�aGخ�����7�\TWW��˗�;�T63�@×N ;w�̚Fuq�ך04�lİ#l׌���F�4���
�;�|�]H��QU��a�q=�'��~z�í�j~�>X���J��
�*������=���~~4�\su���ȇ�?���i�}.�r�Ueee�ej}��z����w�n���kz���L�l׮]���{l�ƍf�ʕfŊ���Î����y�N��
�>C]�tqFA2�h.������4�Y�jˤ`e��p�rO&��/����x�� S����|����1�6�s	����6p�@��Z�=�|_U�O�|�v���Z�~�y�����������bF��Q�-g�����ӥ]\l��ګ�'��Y�/�^�C�z�轩���w\���T�=묳|m�D�Bd_٪�^�BF!N�l�3PۙŹ¡ʓ��a|ܼ�K�3&5f�֭�I.�ɚ
|z!8�!�G���z_���C�q氎N��D:�̞=ۼ��E�����_A],�����BO��U���芦M�6�=��0��hץ�^ꔨm��� �Վ
a��r�4h�����u����PyC]t�s��Za=AM����s^�Bn���!���l��,4����Ϸn�<�q��F��_��W�+��bfΜi�tܼ�6a-t�P�'�ǩDz��W*ղc�R�7�-��j���g./����9�c#�QLfn���Яi,��_�� #wR[jaG��(ܼ�ѵ|������/��>LzA��(�����/�r�~q���xu��f܏2j,A���^Ðz./����qs��7�5�9����*Dз"|��Tt�BRL/����~a�� r�����K��@4<.Gm�ȑ�yc������)ć�7�
_���	�3f̈��mZ���[g�}v^?�]0�U-����^��Q�d��5?����������N8�����ο����|�����^w� L�����V�k�F,�^���.�e����M��͛͢E�LX�{D9�L�/
'̼au�B�ԠP�b���?����ja�z頮0�p1����x���z�Ν;;��A������Q��AE��jXT�q�c����.p�Hd���/͋��Y!A7M|nx��﫹����ѣ�9�c�^{~ޯ��/���UB/ڜY7�/��^hZ�n��{te>e���劣X�j���ޥ��Ɓ����Î��L�^����ơR�q×��k֬qn��u�':�,?�[U�.����&��f�/$����>�h_߳t�R��s�}zbS�+U �����t;��O>�\q���[RV����c.���ߧ��T��ԊGej�Ă�E]����W�^���7���lE�B���Ս~L�6ͼ��k�r��N��DU���sU�s�|1�2\骬�z��(*=A��Ұ�O<aƌcƍ�yڀ�vj� �a+�MsG�쫨�Rj,4�h>�;".����P�Ϥ.�nԭ*��-i�
[��hj-�՜9s	^~1Wqf�/)-h9��S=�ԨQf֬Y|�`%��{�D�F�'M�d���$�.��p�QGy�"��ݷo_V#�J�/$�&�z�+�^x���!9"N��r��ǋ/�h���ZO�4����X����t��?�ج]��؀!�I[���VA6,�}`M~�!�����������Ӎ-�|!N���Qm(��/��Po���*؄��D򺲰��ƬZ��؂��8	{ΗkÆN��2�S��lC�B"yݞeٲeVI�'A���D����/��n�0��H^��W�M_���*_�u�fyy�lC�B"y�����؄��8�jΗx�<�@_H��-[z������!Ve!F��|���y���c&���I����T�'Q���ڗ/���û����ܢEc�t�G��"'�>Z^?��6*�D�B"�ٳ����LMm��#�F,�����6�lC�B"���z����/Y��؂aG�MT��k	�� L�/$��U��{�6�󎱁�^T�7�SU__����Ŗ-[`�iӦM��׷o_ӪU+�ÔA"x!��X���}���=lD�B"�y�&�g[餿�q�f�2Qc�qE��c�9�S	]Ь^�� �!|!����O�>Y�{ꩧ�9s�D��� +CaW������O�t_��&�k��Ş�W�� 6u�T%�Ga��:餓<O����`#�k�泟���a��c�:�F�v�aG�Q��/��z��g{��.f�ϟo ��XnЕ�СC��WW�_�җ�}��gv��e�@�B�5�K{4~��_��\US����_H���~�{��<�l:v�h���J3q�Ă0/'(��(�ʗ���_�y�Q�L�b [��h�7o6~��2d���w���|��_5O<�󽅢�l_����|鳣����l�2g�`+��W^1����<\Q^^n&L�`&O�lf̘Q�PD�IT�K��#G�s�9���Z5<i�$،��ī��1o���9��s=���u�#F8�5y?�.ެvDzΗ>{��v~�].}^�j��P�O�n����T��А��_l�;�<gȕ+W:��m��lث����i�R�-�>��#NHꢟ�/�Q��WϞ=M�=���j���Ϗ��ڷo�ӏ�m۶�&�]�tq>?��yIe͚5΅`;����J�>��3���_�ЪI/+'sE�U�Q�9_6t�(�<عE�d�z�).b�/�y�s��W;W۶a�q�ގ��
�裏�Z�A�BQٺu����촔��u[(x�GQ��ؐ��c�=�l%��Eg�������7W\q����*A\EY�ڹs�s1E�B��P����{�5_��M߾}�~:T�[
_��}��.O?�4C��%���;l����ގao���ga�/}V�N��t��b��"|������E��vZ�N"�3��Rۈ�i�F5P��M �_�'ԷK�v�w��4wԒx/�Az�`�F��&��gA����B�*]l�� |h2��O>i��ʜ�^ڔ�[�n���~�:���w�w��I�9_��TC��/vZ�����w8��A�X�3,X�\� IB�R�$�iӦ97U�z���t�W�{��lٲ��xU'	u��rwU�4��ƍfժU�׽��8K�4!~�̙��䨣����SYY�|M7}�>;��(`��Х���ݻ�T�/ ���:��:���g�z})Xi�P7 ���X ��Ъ.�J홧�#G�q>s�ܽ�X�u�U n_��_��>ݳgO^s�
n��Vg�v�&�(W��V��C[�vڔZs�l~J��!|(t�R������ôp@!��30�ߒ%K�=�����+�l��
V^^Z̆��8!|(�jG�B/��s�뮻�w��ӳgO��i�Q���R���^��4�=���/��`�B��۷�1_�����?���G�y����2��^.���V�����X!�5�+���^���ɓ�g>���x�P6������(���O�B9jX0,����9��r�Ia[�+,zO��|�����򥡬��zi}���*Hx�U�Z��'�nAA �!|+T���R�_�i˜�i(:��E����D�P�+̪�K�����cj��Y
s� �� +�c�6o�l����E���U�|�����9|i�S�۵kg�ݎ;BY��X����&M�t��d�/ bq?a)����"xI��1/����X!*_Q����kWQT']z�( E�4�@v�/ b����I5�֭[x��׊y_�w�/ b��Z��W���Q�c��;�8���ɝ�$z}�����DܢE��{}��у6>h/��ݻ;�j�I� �8j�s�:����kF����X��[�li�v�I'�3r�H��o���A��(���#|RիP�K��p���K�.������չs�К�*��Q���xG�"T�ץ��f�֭&����"]eWz�.������xa-� |����?�*_�t�̳gϞ�SN1ȍ^�W_}5�_z/�1�K_�w�/ BA�h߾����
��V�]}��T����k�1��zk`�W5K0����D(��
D�̶m�L���/;�/�[�n�k�裏���¬FQ��S��oa@$�j���m:�����v��1c��g�ajjj�K/�T����ZYYY(+��x��1���'�o�'�@��tަM焨�{�LU��.�̜y��u��;a��'��{�)/U=�^B�]��O>�;�i��ɍ�D �mft���4۷oϹE���޽�6U�q�he���:_cB�QLtΈH|�h� c�����1��Qc�%5�M�F�^�(x!��`�$N�!�vX�m��:�tk�z�|?I�<��s����yN]�Z�|yz7{�ܹsU}}�jiiQ����g��z��\!��/ o�t���Q J�X��Gҍ���m��K��E�*>�o<cƌq�/�\��'�|y۫���u�Pr�~�2P,�/ ?����f�7
@YLt�0Y����I�{;s�@y�b�(�؟�߀��{�-��v���c�PRL;�L��&����t�uvv�����w�PR�|�L_@N��`p0}k�a�� |%���fB��&y�-]��Woo��n����� ���a6�F'��X,����×�z��|k%�=� ��`6�|��K�-]ޑ��p��H$�j�Pt��r���J?n(_�W��<6�t�.]�-Z��g:��]�G3�4$|��]��7f��U��`���=,�F��J9�u�� HgL��t�+`MvL;�z(���Хmhhx���{�|I��=PdL;�l%����o�|�+e͚5C~��F��V���f�G�8����}�䚸IWG�R7E�YO �M���rX�E�I�H�l_�$G�����_����cġP(������P4R0=�800� �=�F7g�����p�I	`Ӥz�Ppl�
�a�=0�H$��h?su��|>_�0�GS�@A1��a�	@��S�H�s�0�)�����P�.!�L� ��fC���I����h4�n������� v��lCӎ0��J�ϷI����������7e���}ss������YB�t`�_0�|������F"���I��v����I�~��ů'�R�C^�
�)��_0F�`����t6^���]��ٙ8�??�툃��?R</����ϟm�uR�Fʋ��^0#=�Ź��s{���|/�|2�Ϛ� R�ht����|>�Y�P.���P��}ơay���~)�;'���F���Y�iE����藜���ܥ��Ӑ�Ͻ�:(��?���o[[[��� .I��cAl�0����5"|e�f���O�b1LVuuu9О	_����+W�U N�SP�2`�fŢ{ 7�Pl�
�b�=��(�̊��F�J@1r:���b�ȍ�YGG�����镕����`V6�
�W	Pd�d�T*u�����/}��nW��,3�%�<��(_@���yR,��g#��v����TUUU
���K7���ȑ#��N8	�(���V��t]�=�㛾����a��m��k�$���9G3�K������6��/�H�z\
�������x�̙o�ڵ�i��(���T7^ݼy�.�YF�� 
5Jqg��n�'u)���T*ծ �J&��'�����|���l�����x�ޤ�F�
l�֭�x<�^�����S�~��x�+�zS&&A�~	^��f�i߾}OIy��F�
,����%�.eMM�KR]]�M$�J K?�4�J��D"��|�� �PH���+��̱���\�U
��J��3�O188x�^�%���>vK �IG�
H�����)S���p8�
������kkk�>x���>wӆ���noo�=o޼�
�0�P �p�z)|�cix�JԤ ���L�ǳ�СC�;|��<#ջ`a�/� �l�rf"�x6s�t:���'��l6ۇ
� 	W���?O�7K�:C̩�����3�.�����o(��_@H�ҽ��u]/�w��5�Tꯊ��Z`MMM�I�����	u���.���d2��ѣG/>�k�B�Pw �ND�&Hz�WJ�Z���[��~�P\��
	^(���^�^)�ٹs�3r-���x�=p������:ul]�;�%K��� �!|���\!��A�����I ;\YY�Bcc#��b֬Y�Jqώ;���ɲÇ�(Ǻ�R�p8VI��,�_�&[�A{�    IEND�B`�PK
     uK\���@  �@  /   images/c19b89aa-68d9-4a98-b509-123aa1ab0169.png�PNG

   IHDR   d   �   ��6o   	pHYs  \F  \F�CA  @hIDATx��y�dU���{VfmY��U�������J#��m��x�x��q�̙��?���s��c�>}�uԱ�pCYD�Ud�������ʬ�3#22�~�o��ŖQY�����w߽�����{o��W_m�t���^���w���η����r9����d,|�k׮����L��oTp8�m۶�����$����f��~&����^��}�B���M�u�{m�®�.[�|�9�x����ȈMOO'�{x�$��mi�-[��z{{�����;���رcgMNN~����{m�-8�A�s�=�֮]kccc���۪U�lpp�ϔ��8@�����7��Ͷu�V����1�v���A./ff@ 7�̉"s��իW3�lvv��LX$tvv���|���zf�HnB\Azt1�I�ѥ���4<	����<���o=E9Ǘ�
�S��SSS~f�����'g�� ��StȎ;���@t�D�@=��G|� �����3�I ���l ��2K ��\���3�y .�	 	�mi7iF�$F�!�%��D��]|��
�Hy�� Yw��m.�c�%^��1�˔:��+�
���s^�I�4	�9���� ���5[B(ƅ�w����{B<��#�r��"OB� ��{��g�u�.��?����ѣG�i����鱉�	�:"��,Y<H�c|L`f��R���EK������E�V��x�����������y%Ozꋇ�S��=�!��`<�YY�"����g.qN��Y��BW�O D��^D�.8��h.�9��A��'�?	̓4�f��n>	́�<u�_�B�''z���SǘR4��SG��pq�D��$Js �<�8��@��9��d\p��Y��[>��o *r�I�4*"��ַ�նo���׿��Ǳϑ�7�SǛ�C�W__��M٭4PB������!
���@���"�L�^Bp5OS���Ѽz�xϞ=�!C&H�B�_��3e��>��>t��>M�;�5�b����^��z#Aĸ ���paC��>}��h׮]EO�,�0}�A�:�8�V^w�u^)Q�7����mbz��{�sv啗۩���9� �����Ͽ`�om����l���˞z�)�U:"���Sgf��ˬ,�pf0=O9�o����[G��m��MNw٩�.���v��w�ůw@�\v�e�	O���=kS3ݶo`�gV���/�\&�D^��=�$@��ʻ��L�F�;�4����x#)wDMk[��y�t�#�S�)�4�4�� >���e����:�i.��Ύ�4����YG���6����#]6�o+ƭ� ǉ��4��n��w���B1��޽����8��N=e������7�����|�+�{�^�1k�7o��V��G��|a��D��>�Ӽ��,8t萷"d���_^T�6?b�zld��Z�6{b����A8���?�����ّ����m��O<�w�C��ۍ7z���Ç���Odb]�����H����1�z>?�f�z۶�ۦ�60z�k�a]	��y�mݶݶ���L�����q�i����/��Moz��#V-�$z�P��z����%�A )���9�y��f�坒�[�GZ���ӫ0��T��,���?��
-����1x� *��e!aW����o�N��x��5�<��*���8�7D��dm`�9�]�N�wz�.�'/����KR�RN ��Cqf0��������������;�;N��Y7���o�7Z<D��G?���t����O�U�_�P�$�'�ԙB�H�䩳.wǰ�c��Wڱq�9���#��G�����N�g���:7;Z�y�����+Q�I�%�*\2�h�����ӍX��[[gm����ɵ��X��=��~�B�|�����ML����{ɡtF��H�(O=��&r���?��VT�>���0��l[d�"$����և�ʈ��sx�n6M;��ҲscN.���(g�۰a�����#G��uv�:�Z)ut��g�v:b��+uD��Dbƚև��T���,y�7�|s�R�wJ}�S�7���2�jF G�>�l�7	Gl�W^yŞy晢1��4cP�?��O�RoqJ�-P�0o�?����c.:�a�4��P��j%.��AB� �����^�3C�;�m}߀�:��ʕ:�G���|���8:v�g�{_}�U���䘒7�H&�	��T������b2N��M]����>d(���_k]�{��)��G7�:����sO����	�n�:��L�(�O]�əg���+l����=ԍ2��H�9?i�z�G��(uڤʛ�4:��ut��$u��{�{��� >9~� +�r\�"���]&;����B<08������{� �He�<$��kY�O;���/f�P�=��-}s66�g=�+����h/[Ɍu�az~���$t"n��
99�II��%˔(t�5A<���K�-��;�������Ђ8 ���mo��TY�v���@�8�P[�l�dp������hj]8ϧ<�v�K��}������w����Oz~���~f/3�6��ݻ���c"�j܄✶`�0eQ����)@bC\-D3X:����9mG[mȋ�!'�V�c�Z��@��8K9hKt d�0��=����:��p�kA83c�Ν~�;���Ċ��l�|ӦM~Y23b�F��=���h���!:3��Ѷ�d WS�9�����S�Ȋ/���8h��-/�,����Z�_:���M��-��R���R߸�~S����L]�G�0(�ϋ���:C�Uì�M��� �gh93�l��z��;�h���-���������1iO��34����m��j���Rw��%�S�ԅ+1=��}�1�͌/)r�Zz����̍7��o�Nۆ��n��N�o.r5�� ��������O?�����r�9����h|���E���<�6���zd�)�LF`8�B�ILr=��|r`�c�0�Z�7aeL�gv�-k{ɺ���`cq�<��Cv�w�)ˋq�;𭱔���!
��k�DQ�o�ŉ��Q��u�z�Eޡ��]!���F�^�(��;~�Pp#���p$bF� d�]����"��G��	�"D��������L�ߵ�)��P0��>'�&VY[�2��"�IɩJ8NͷVr��Xd:ˈ�VD��.À�%m0($G��~Q����p.�w��8���Ԓ�r��U��6�%�"�J8ikC:DƎ�^$��Xl��xN��(��Y4gw;*g�C��\�Ag���=T�źb
3+0-��+܊�b&T��p�0}����͒9o&wJ}��)��p�@�/rgH�E�,M-U��뮘R����o����g`� �;��6hO��j޹:��$����Y�T
F���HC�`�����>K�׽���<�Ce�z���,��5^�GB�)u.@~#J�`d)\�NnDw|��J]f例΄]eӳ�A[+"A��TA�(y�\�������[��,/~��I�a,�)0�������2fƊ�a����{��u���I}���'��s�3r����~��RH}�w8�������H�3�x� ��Er�<u��Rr\��x�s�67�e+{�-;Js��BjK��������(~D\�(w�S
:�Zh�	�с��c���������� q�?�|��¶���+����j7�C��]8�c��3�� @�z# �$�N�/�/�ři��!�s6�k���R��X���1���%����2
Ƭ�j���1��1`>���q<�����w��]ރע�R��tn�wW�Z�[�(׾�qS�
�eˢ���b���	��I��Q��G}��Z;�X��4������">�\��@b�`~K�u�d8�g��4q��b�ţ�>��
���X�p6&y��Թo��C>�~xh��U����x���)Lq=��y��\���5�EK��K)S��<�믿�iV1
�-��4;�/p3/�K��TmK�S����3[��A�N���_�/q�=����ّRom�C�X9$�V�q�BK|�=u�iQ�04�겨:��-�mpd�M�Lٌ���<\��M?����)��u$¡k�K�D@U�C$2W ������n4�V3���{����y��Wt��9�Wo)*����n��O�Y�����%�%�SWy�>'qY��y���I���w2eϚ�9H�Vy�p����͐C�1znt�!���;܃q@>D�M�N�Q��2��Wo����ybI�)�%�U=�j�V�3{�[s�|Y���0��T.j�23��@C���E�$�A���UL��Hȟ�!VV3��,Aġ���!7��Xޓ����^ͷ�6�S�� �!Q^�|Б�CN��Xk{މ�ӛ�C4�1]�W(��d� �x�� 3�$�]��A��0��A�+tt���Y���ĐR����A_�;pl��U�>�E֣�
���<u�%��ee�,����@���ݠ�Z��ga�a�`��q�.E	'#jH|Q��9܃ށ�p?3Ŏx��,CW����8����o_��[Z^)���q��V���!%a�t�B�+8���4L���n��@�O٩�����j�C��sMQ������X�^�?��@�a'	 ����J�Ae$���K"]�f�]w��Z��+���N)V�P$w뭷k��xd6bR�68�<um5g(T͋��o������v�ζq����J [�-�&��F�1C3S)��P�q��'�*у����� 4ס�A�f�r� "��J�)
v��������ͬ���#
�ԙ��G@����'Q�k;��ġp�B��-g�Vdmb:Z��?��X��,\+q�H�yI
P��)�z
�Q�SDȅ�Ks� ���! $�eV�U��"��"2���Χp3�o�M̴��wp������5��2 $�+m�7SK��w��,�Y��{�F'�Y{ׄg%�X�!&$nS�˅�)^x��p�( ��^E{�6/�L[a!	�$C<��b�[�,p2Hc�IL�ټ=����ə=��q��辢RW���e����9M��u�Ћ��G�F2�*�GL����Y;���e���伬q
�Ɗ�X�=�\�� 	��uT=Ev����v��H���B�&�]�ݻ�e;|�c2���7�z�d!�(�	^U��'n5.�E�4�*D4�A��^��8����3��q��j�8݋�aٌ�Vޜ�r.t��Q����nHt,���A
}	�M�&���R�������:��]��y�����_��$=,GW�P�U8��|A%+~O�\��z�ω���l����b�03�*��8���5Ē����kyD(7�Xh�|5
���l��65M�s��M���q����Ƶ+���S��T�m�>s��lP%��������χ'@�2��Ua��$.��=q/���C�����17�F����d��7Cz��j�fo���q����'@3A7�	��%g��9K+��o�W�s�s>��P�x�
�1K d��U����ﱞ~��q~)�f�"��� �x�%s=>�W�+�W%�B����H��}h�OLes�����$O]��q\�ˋ�{��**�]Te� ĳ��Te�t�.�&f�t��-��N�,�ĿPԀ��f-�a�b5!�����9��8�(pz&N��L\�g�=����Ћ���7o�b�v>g��)��;<A�Cp��L
�~#!W��pB*X&/�C�@.�ꪫ�*���ؼ���04~�Y!Q��NўLV:��湹bT�� 3��X''E��M�0D�(r��ӵ�2Q�at�T�/��qH�B����N|&�ޞ�����%������}���RǺ�P0`tp��c=u8I����tT���h��ڶ�+��Sjq�NGH�+�����:�3��M��� Q���
���FE� ���;���f��|��W%%b�-oy�o��d\}}���N���N�3B��eJ]yma�>�Sזe"P�`X$r}�R�0l��"��ϕ�:�@i��/�,��д��Q�p]����<|�O��e	�h�>D#���Y�7�w0�*�r=�@_�� �k����?b
�!x6��:��Lfƶo����]����M+���B�C�V�S�GbGZ�����LC���c��l�\.c+W�u�Ӆe���aP��W�oVr=<���4_�$c�\u8˴n���]�1���� ���{� ]�]0w��:z�Y����Y�!-ŔrȜ�b�0X�`\��- �7Ɲ�b��S��}�����3L{%�B��(/nb��v��j:(���k�����&���t�@g��_Y��1����X�op����K˔���Uvt�/��8Y~�җ�bM��^�͸V��٦՘��k�6���u���Y�J:��>�D��9�~���s�J]3)\�'�ƴ��BO6����(�Yq�u�|����4��
�^`��K�u���=oIJ=�iM���^O} E��3P���p���3�$?Q�XQp�`�i�"�0�1 T/�=C0�1������E�`�`�q�Ƣl!�.�`������%�8��|Ͻ(q�����{Ď�����҃��S�O�Z�R���DO�FҎ��3��E�0�w�t��9���Ї>T� :���i���n�@ڗ	��iXB8c��!���O!B)��A<�GT�Dܧ�*�� <_�̄���6� �i_�N�]�����g������>�;��}�SoI�V�P��Y�����
��nd��j���5˷(t��:��}�Q"�V��N��Df
N�*P����j%-��>�'8k!;�iL�:HH�~�]Yj-�"�H���~�Rk�L�Md �gք�w67�'*�R�D�}��0���8�P0jd��\D�6�ޠS�I�S�~Ɩ�|��ѱ3J<u�y(5��jGg�RZe��� ]�����	$1�~�_�c6�;��]� y>�:�s���Jz$��!σp�,f1�1!.�2n��wz��.x��'12���KI婓��1�@+>��1pM�`\��q���G�-M��\��;��)��2O�6��i���ɫ���H���\��6��c���K�-/#� �N3�C-7`l������1c�r"r>E<�=�����3���CC��ӕ���r;^ZS�x(�ą��0p'PN��
JI���a��=�Js��l@��f����-��;�����BsQ�]Ԟ�����
�䆠E�Z?���X��R�)E8���H!A՞�S!i_�b{�m5�s,�KHq"x�<����~VL�f2��q֮]gW^ye�c��ǿ�_[K;a[ծ���9Dv�w��Y���;�^qJ�Չ��ǋ�^fm詫�1���Q�YY�"U��|E8xU~@���Y�G��"k���u�E Z��u�i{���c'�W�XG����Q2E�Q�g�������ɴ�琓x�yt�_�1�s��c+
J}�D��݃Xs�b�������g���S?�w��50c��tഢ��d�.Đ��q�С`aN}�)�+���^�SG��� Y�I��p��?D�\6�:5^ 8=��ḡ�ƕ�z�'m�Z���+_����L�B�.�a�n8���_uR��=ǉ�h��n�f2Ci�S3P�p?d�qfI"�_m�|�%���I�,(��;g�_g8o�|0�b^�<h�EYF�;��6F��zɆWA���S�=����e�J�<�S���/y�0���l�ַ�m�Os���z����rk
�>�!�__�t6����Ԩ�H^(m��O]'k��<��^�&��;�>�ޔX(G�*�|��I�e��7��B{��=u�:��U�:�)3��
bq0:!z,[����DT�J`6���E�Sꇎ��'��gY����۬(��B�t���tv�'풔z|�^��J`�Ҡ�b���j�nZ��&�[��)�u����p��tOR�j!a���%�f`$��l!�G�OR������ͤ<�R[i�������k����mz�W�I�,��ʞyVĻ��j1�D�2.����罷��j��O��.�袲�fu�|aﻹ<�Pp�]\&����4p{{W�\vڇ�	K��̤���2-�>x�Hh����[���=3�p{Gt��r���|7�X�P�퐝�NZR"<Phͦn,V����-�S��c������:�����qS��x�s��,� �o������;��fM�}�K�X��H=��~{��=��_�·����O��ᑼ��O��5G,�����~ж�v�]}%��l&�j_�wۇ����{g�q*Ñ��}���k���v��ӟ{�����O�g~�V�L���{��k��a�}�9$;��t�7���3�������}�l���Ϸ~cW\�v{���К�/O���?wϟ-�xƼ���B1dĸ��!Fx(X�.�)��䇤�"�!DU�n��R��e�]�����Cö���kz���1��a'.[mY�A�d����65��:�:�w��8�{��A�emx�׺���gY���l���ۭ-s�����MLt���Iw�!���������w�&;��Z���g����q3��9�����:20賡i1���Z@��q��V㕠4
Ad.g����K�Z"��~�^9�ř�]6>=g�3Lg���ՆG;l:����'�<�t��6owג�x�ӷ��V�ʶY~�!čdht�����':�#֞��R�Y��̉�N��l��egW�ﴩ�^��6�v�ML�t�������C���6<��Aü5o/��vR=�$e���?R����+��l��nb��Y���F��Sˬ�f�]�J$^��Ғ+\�����0 �
���6:g#eJ���6Z[2~Ov�ϻ�:9���Dm����{�v*�5���!t�1m4�EH�q�Ȓ��p;I��Ҟz �_�΂�m�_�m�d$�L�ް+�^�ni��uUx%��V��w�m��0L�SW4$�S'7��L�CnW5
J쫬_�W�H�K������
1�E�W�A���n�L���L}�3�������V�O΄��?�M*Q��`�1��B��ύ�/
�Zd��A�u�B�Q�m� ������FJ=�V�yO_�O��tZ���"Ֆ���7=�{��H��8�*4
Z����C�xVխ�U�"q�S9H� ��R���ַJ���Ǫ�'�~��!�������w�S��7��Ͳg� (�$���5T#��)��u(���ag��!������Ӣ�$���]-��jmUڜ��/����H�W�S/K�j1{�^B�`Ǘqo�6�P�W�C��/f
�R��Ht�`�a ��%�y���I��� '��\�G��@I~��a,�Io,��.ߪ¤�Z���c��ZJb p5Ղ�W�*
�%��XE?�����(z�܇�B�f�1��Юs�*g��*R��b�gն�sEO]�HhiaЅ���Ì�[[�EH����w�1�Ah����I��6
u{�i�C�7������Gl�3_��$�Q����1;����"��,�]���*F��()�Cj!JX4�H�q�`aN=<l���%c�yg:��[�������v��:t�V�J�/���P0:��B��k�sTS���;k���O��~���^%π���&�H��,���%8��_K1��5�P0��x��`:�d)�לCt��c��3g��++��=���i�(~%��%�*�y��g�W��^�(���V�ԵF�i��_�������
}�������Ml�0��فؠf)�z��A�X�g��+� ��#%[Y����"���y�F��H��|���߷n�Z��TROC%\/��\Lpbq
�h�|�`Z3��ұF�Ԭ�ȺI+��"��<����� }řT�����F���
�zg�E�k�$�j���	�Щ[�W:���-y��е�\����c��C?b-��uk'�pg�$hDLI/��J���@=�b���P7�cڡ`� ��+���|�0�Mvhh��pu�����cc��詐�~P�QW@z:<Pr�<���y[�� e�Z��Kt���h����Y�TT�x|�AR�R	z��?�Ŧ�������������;�WZg�JkimL��@�lq��phen����u
��`���\�/��x?0��23k���>m\���I�g�hA����)�l��.q�3������kP�7p�hH�`�	�)-ʍtb��8��ZT�y�w�a�Q<��h�M϶��)M�����kS�Y@ۄ�ò�z�1�S�@^E����J<l[a�r��`���fA�h�LFj�����~;ڨ&�X�Ke���O�-��i6���� Z�ɚD�R�[ӡ`Z��褎�x�fר����j�@��˴v٦-ۢ)���vv;��]�L���W�,|��Z RAۚ�A��C��tR�z[�����Bf��2l櫱o���#v�]w�r��4f��2q��9�@�̨	�j��Ϩj���ŝ2�r�o6~(X} A��{�֞s\�R z�r�"�T�T�$�o)��FA�G5
�Ӹ�` L{� Z�ӈ�Y?�p�� �?�+���0�1��!��^ӡ`IV5�pDa�dR��C���F�*%�e(T�q�j$S�JbG�ol>:��vtr�bY*F�!ȍD��J{�7q�L=L"+<a) D�t�����is��U��l��{~ǎ����C�J�i��� �Nokt�	dJd��l�`<X9)��I�loO���96�?痦-wV�l����9d�����d���ַ���@�6L[L9��j���M)��U��S��r��4奰X@��̴�zi��G���������U*5��܋���bKI1T ;yCXf/���Ne[�kOt�N22�h#��=K���s��wT\ti��:��e��FbZ�I
=����-��u��61�H���i����R���[O���e�#QK[���^�R�����W�LvƲ��B.�U'&j߿%����x(�3��*]R/��UnF^{��m���^���o�Gw؁_�b�	���}����lW!Ⱥ�ϼm۾�6n�d���n[X�[���¡`T��^�`*
��ӧ��k���V�+CV���;瑲����!��i�K��]9f�l��� ~��њ�!С`�(�� OH<,~|�b�^�g��,�~���n"�M�;88`��?t�Q�s�������Nm��N���F�����8�%D�D�!t+Xj���!�T3j+����+��vbͪ^��}g���o�������r����B�d>���[�RX@u%U��HPt�%��!µZ�O��^�@�Ç۷����hů￿�����B�m`V/�d�쌍����s�Ui3�I&��~[�El�q�]wy���q�ؽ�Fy�N��HZ������>�����+X��=u�5hW�E+�L�:�a}�8	+�Y��:��:߱�T[!a�c�����"1T�aPK��0s�e�ZNX�c�Ua]�%B��Z��g�;�z����W����S͒�G�thm��U��O�ď��i����P��њ��>&�_/^���; m
�O�;�����D�"�(,�Q|�npؾ��{}����w�*Ah��e�*�#���J� a-�(b0c�gXτa�s��g���.�H��*��HE���Sڴ�b6'�Ȋ��P�Z <���s�vFGU[bL���3SK��PҪ�m�Q� �aT�w�obB��a7�p����~�9�I'hV��
�"��������Փ[Wh ^*�0�/��Y��{�y���o�q�R����	q� 	�1 W�v�mU��&����}�e�tφY�J�Z�"<���e[�K��ˋ�Y�*vH`���o�{�)��E��e|q�r�-p���r�,d�OĀ�"��Ȋ'����~{]���$��֮�w�o(��Y�(%�N��y�B�Z�C\\�C! :_ )0��k��͛6�c�}�~u߯�C���Ϲ� ?��-�cT���{q�,�zA���}������z��֟�d%�3^�7�H
�&�! $B=������?�����A:^4�X�}�Uk��<�����[gv��.�8<��W����C(
���/Ln*]�I��Zg�JȣHR�O�_��g�8�i��X�s���<a�\Tq����{I��R�X7ZFp"���	$.iK*!SObF�ƫ�T�ձl�u-_m-�c>E�ֱ�}^k�Ǌ�`�@�fC}A�����439<٭V��F"B	�rEfc��b.ƾ&����;��"!1�~���ӽ��Zm�������\�p�Oe��#Vu����zm���ʺ�⋽X�������Y�@鱰�k۶�ַf�=��53��1��$D5�B~��bvE�B��
�	�5+r�/�4��E�<��S>���g(T��a�6+KIp;gUպ�s���D'��濮O��]� Z2�E	���	"$�!`G!0	����s)�Z��C�����g���ޯ��-�iÉZV�z�i>���:�x�S��'j�!<����������/��Y���L3�X� �F!�����tgi�#4km�fH��4! ���[��Gml�t��N �J�f8��"u�0��}:�Q�HI,��_BE.OD�ZLΰ2#��D��gW^v����J�sy����=��o��Jp2k1������DlT�ޢ�N�~G��g�c���RKY�W�>06���	B��0��^��i��N��N5�rj�Ӷ�a���7��ͦ���E��o���H	ḏN�?�Z�T����Q�`L�-�Z����-UII�G�t���l�2�%�iD>V�������}��"Xf:N�LNM�o�������q0o{O��(ž�-&i���\�b��Aǡ�08́����`I��F_d�B�H檶�����Ѧa{~�'Go��A��.��e�*߁A���ŀ��֪�x1�|aܡO�F��ހ�0��-� +��vx�tF�j�9 nX�@�;��T/z�
:���"���I����>N�T{X�}�b{�������X�]�Ү/�ԁ���U��V�� ��XZ1.�!�#V�W
�)e��-��	�i�L�p�i��r�ŋ���M�.���a��	�W�q"���=�N������9P� 9{�5�x/���.����>���xՄ�����!��2���Pׯ�`gl�`���j�k��=l�pF; ��Vh-f\�V��I	�[�cr���a;עԛ�<����='<`F���� �lS�f��?\�q�&����mt������i�S��!'rCq�3	�.&z�}:L��E��
F	Β��C����T����i�T���?�H��O~�}�s��K(��!���du���yN$<2hS#�N���S�%c-:��w5�)���v�F����,�P0 ��㇂o��kgz_ݵ�y�i�섷C;����\�O.I�3#�W�i��ٵk��yi���;�������b�6����`tR�|+}�L���ׯ�ٖC6;)�e�WY��j�{<�\�o%�&g̼=^���A�fm~9WH_��Թ@��<umCWK�*�p:v�����fm6���6g�Y���M�p�o�����(���f�=���޵�lF�u !H,V����X���-e+�`Cd�R���8eEUGȝ<=$ӳ����o�5����ky�f�Z��j��8�z�6j��s+����=Ņ��G�MȤ����z�����*����8�r�L�t(X�����/�9qBXI>	Ȉo��n|%T��Ç��>e���ur�է���01�O|�E�0&B�
j�D� ��zŋ��@|�*NW�P�|.G|�-<�q�P+�u��5���$�5CZ�|�5l5y��2�f�00�?����O?��1���=�$N�G?�Q�Ⱦ��������K�������g<Ls饗z�s���ӟ������^M���`���N�l�����4��=�):jx�7�tSIp�xZ0��u|[F2^����_���/�6T�0��]"��`$��"�
��J"�����?X��i��bG��|�u��c[�j�{3�1��mo�̦}���BGq3�ZH�{��I��k/<�
v�9�me)���3	+Q�;�Bt�"m�%a5}�/���U5��J:A��bm���A-~�j����#�I=�u�k�C���hs����>1��p�S��̭���o-���6@�?��?O��	x�E��
�3�P�l/#�
VII)B��r��`~�k_�m�k�j�lC��4�)�{��L���d��"����([�� ��կ~�?�V�C�`z鎲C�D}m���JV#S[�P&���/~�����vVΤ`�B紉rU�Q�%��ȡB�'էD���jǀE���j�x6����t-�� �a4|������qS�ư��*�� t-�+��P��
7(�A��nZC�=��Ң�T�Љ�E'��,��<������ʊ��k }��I��܃E��(�1�x���B�jSY��$OiW�j%A�\b���=;�i�£�kڦ ���g�ć�¤�}$���:���~ţ!!���ոL9(5t��Ppe���8@P��fgX��w������G�~L������{f_�50�\��
(�.��[P�&����íƫ�2�O}�S~�}�{�����xm�7A���!��E�@#��܏>KPK4��o߾�����܋6)c�H��W_]sͰ���㊇�I|U:L�G�p)�CĐ�RP�t=A���M��n�H.�l��	)"�a����k��E�&Nܕي�$�4fߴC�d�j+:��Jy%]�Q��Z�j�2�R)
�8�0%�1�Б~�(}TmKv���Y!&��c�S_�Sgfh�5��@?$
�l�� ,���ˏ��(ߦ,v��z�R�bfD��՞�Ic�X7�|s��"��	N!0��Q�!�����ߒ@6<���J��*OXB(�X��X��,����z�Hd��"�p�$��p�@�2�F�1�4����S9�rR�3+LBq4�� �"�5�s�e<`�)� b,A��C���G���^��/��ǰ����������$�U��K����C��%t�ڡ`��u�VU�����OZ&���%�,����L�ȤXs̐�qb+ 3!F��)�s������p`���h�u5�?"����pSSX�q�s�)"O�U����g|��@��(iGJ2l���XP�n�z��	�U��	���L�6 ����v���	�o,̩k=f-���z�!��v(�����.�-^�M�\O@��E��������/1��n��~`_���H�e�� ��Bq2��B���0\� ��=��z�����
&��('��ET����1��#+�QPuG��Bd1���x��-�(T:��^H��q��=	�͒B��ő"l1�t�<��b��ɛ����$Xr�H�bo�۬n��F>�(_J/]}� ������>ۇ�	hB��::���\f� �5x���Jӆ7K	2J00 4��vDo-e���$*p��t��G|q]X�ΐxV�\ᕀv�Ʒ�P�y�-���b�'� ��n�X+X? � !���/� \��G(�<v=b�oM�o_�6hH��"��l/��NA���`�Q��A:�	D�c�EװT��_�r�"� ���WYk�D�h���ND��	% SS����>�O��n�������)B]�'�T�$ahC���ϖ�E(�z�[�:uB�עc�
^S�ǚ��LP���F �Z�s�;<�%�v8�q��b�DaQD��g	��5�U�՛*��� (���j��E�!�5�����x4V��B�D#�+fɖ-[�n�Z�tC�'�A�޽�p�NpgJ�X!rT=O(���yi���2�IJE�H'�(�w��{2�p��Џ��K݋�/�0u}�s��q�ǜ����@aKܹ���[]7��,��b�$V�qc��I�9����a��^Kp&b��o�v���Q��Rq����o��o�!\��3�X~KB��}���� B'$��뮿�����N��5c�Z��}։³v���o���/��"�Dޙ��j����D������,���Gz{{��ݻ�? 뗒9
uR�ܬ��������o���?�w�^j���W����T�    IEND�B`�PK
     uK\}�?`X X /   images/f6e2a5fb-4294-42a3-957b-9521668fdddb.png�PNG

   IHDR    0   \;�   	pHYs  .#  .#x�?v  �eXIfII*         2       D   i�    O       NIKON CORPORATION NIKON D800  "�       '�    d    �    0230�       �        	�       ��    40  ��    40  �        �    <   �        	�        
�        ��    �  ��    �  �    �  �    �  �
    �  �    �  �
    �  �    �  
�    �  �    �  1�    �  4�    �         �         2016:09:27 09:37:50 2016:09:27 09:37:50 Тt @B O� @B            
   X  
         3064640 60.0 mm f/2.8 �/�  �iTXtXML:com.adobe.xmp     <?xpacket begin='﻿' id='W5M0MpCehiHzreSzNTczkc9d'?>
<x:xmpmeta xmlns:x="adobe:ns:meta/"><rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"><rdf:Description rdf:about="uuid:faf5bdd5-ba3d-11da-ad31-d33d75182f1b" xmlns:exifEX="http://cipa.jp/exif/1.0/"><exifEX:BodySerialNumber>3064640</exifEX:BodySerialNumber><exifEX:LensModel>60.0 mm f/2.8</exifEX:LensModel></rdf:Description><rdf:Description rdf:about="uuid:faf5bdd5-ba3d-11da-ad31-d33d75182f1b" xmlns:MicrosoftPhoto="http://ns.microsoft.com/photo/1.0/"><MicrosoftPhoto:CameraSerialNumber>3064640</MicrosoftPhoto:CameraSerialNumber><MicrosoftPhoto:LensModel>60.0 mm f/2.8</MicrosoftPhoto:LensModel></rdf:Description><rdf:Description rdf:about="uuid:faf5bdd5-ba3d-11da-ad31-d33d75182f1b" xmlns:exif="http://ns.adobe.com/exif/1.0/"><exif:DateTimeOriginal>2016-09-27T09:37:50.400</exif:DateTimeOriginal></rdf:Description></rdf:RDF></x:xmpmeta>
                                                                                                    
                                                                                                    
                                                      <?xpacket end='w'?>H��?  ��IDATx��גdWz.�����wUu�G��9��P� ��a�y�s���R輅�tAJ��3���L���6}no������6 ����Y;�^~��8UU�2/�Y�8�O�w��������`mm�,����<
k(�;�b�_���_����������׮]3�k�f����4����������_��O������o�Y�4��@ʼ�l�0��4z�F�l�q�lחF,�K�<˲�Fmcc�*K��*L˺��|)��=}����1/��߷8Ƽ��kTH������ ��$˲���<�,�1+��I���oxj�y�jv�.��EF�W�g|{k�`Gh���R|P����Y���)�yy5�m���V�N�~��'`4�{Eam Uynõ+�
#�۪P˱���D��SU��ڈ�:��[�]��\��HЬm��%9�/�D��E���rnf�Y�˫P�hc^^�rY|��` *-��|����v�m���� ����ׂ_�86��˯�ik1��lꙂ��EG�����|̆�'I�;��mDa�2/�=�m���X���0�-�4���0�V���u8f�Ӊ�3��eQ�Cq�� ���b(R)�23P��c�6�4%&S\a��0*�P�fe�Y��hØ�yy�m��kZ*SU`(� �l�Qei�����!�e�
�k�����5���\��3"�@Q�Po2etT�b]Ȳ𝂵y��W���Ƽ����� @�7�M|��%�*�*�"۲D%n�iV�eaؖ�9FRLuʠ�o�~r��}��kn0e$�U'S]X3�Hs�L2�>FY��F^��暎y�~�m��kU.S�UiВ
O�d d���x\$I��ph��킡�,�8��0L���b�q��6��m�9@jLu	O|^���L�1�l�e^^�2G��Z�)ΠU�e�i�!u��v���7�Z-����|e�=�I�Y�e9PGI����in��/����/�=|i8�u�ě@9�T7*��a<Җe��q���ܫ(G�0�� ��e����WD�>�ȝ�W���Ƽ����m O 4�|����(��B�-B*� \�b�.�Q�`*R�S���6�����
���(*������(ژ�f���W���Ƽ�V�9!	��@�Q�ꓡ�'@q�uɝ8���k����Is o[-�L�2�?N|d�)a;��D�>����2��ʊ�opN��ʋ:�2/�s���yy��s�9���LL���3Ė�L��W���$q\��S!�%}�wT9<;��ҬKT��.y��4��D�(
��:���*s�1/�Uy��Ϡ���j5J�� ��ip�� F��><+���k5E�'�*%ʢȣ8#�嵿���s�!��D����PR)�GYYf)��_������˼|/e�6��u,����wq�����LU��x���$��<D5��Qs<�uW9Ku��e$����K����j�L^M�`ћ��iD.���e^^�2G��:ڼ�F��u����CcR5�M �2/�6T�`Y6P�[��i�~Ey��?� �`5����T�e)��Р#�=e^.�R�*�R�s�"}^��*s�1/�U�j�q�'��¤*��V���7��2"ya�)�����3��Z��Tƅ1��4k�P�4�zj\X��8�y��W���Ƽ<[���h���mS��lǊ5.!p��4Il�
ꍪ(�*���"L�N�j�pnIm����شJ������uw�d�m�-�r/��o6s�Vі���u����̨<&�o��r\��;f��yj+�Q�0G�T_�P]t<�������Ƽ�VeJ�_ u�c�'i�[/A�Q���$�P}8y^h �8�����#����?&�%s)A�T�q�'M��\T�;��˫V�hc^�-����5�� ͚��P�=В�qETe�e��eV��k䖝TeTVqe����en��W�\#5����ʖ�z�UHuiU�јi��aKf-�_h����B�yy��m��kU�Ļ�d ������phf��Ғi[Ԑ�V�B͇Br�:p��؂ �?|�$��T���&U9�c"w�m�˫U�hc^�)?pՆ�Y�X�~��c��(	�,�	�0%�k�yV�F�
�o;iYeiU �8nR�A\:���f�aU|G=�9<E�Anc[D3y�߆����mH�Z|y�\>/�`���yyK%��hC|5l[��E�J��h���U�ap��W�6��[�">�� �3nc
w�yTײ/���0<c^���+s��C+���o_1	J�<���E\�/ɿ�_��aB��4��ziW�o�/.�	���[�]Di��4�XYD�*N�y��ߍ���$	b��� w;����լ�����^�>u��9/�2G��Z�ؙ��~s ��ՃA%�_�0���g��:b�+��`DE04��:l�)�g<��b��!��e^���m�Be&�0fy#^(SQ����J2�?����;�=��gZ��6-@]���'"&۶'�	j�ᘩb�	<۵,��ne�E���(O�sI^��{i�O��z�^Xe\$�CD]>��x!l�\��!y��i�ۖ�S�eX�QQ�"_4�_���Vqٴ��,O/]���/S.��_�������B^��_S�����㙗W�����\f�a��Y2��r�.Y�^ʇ�_��3���Ͼ>}����*�� �3��{Y�lG;��h00�-S3�y:+�$lUZ p��p]w4���zlL��\���T�m<��/����J��{:}NG�%Ui�3[/�+�7��(oMӘ�+ �}=����=+�r6$hY�}��F���8�U:���c�{��a���m|��2��&�/űx)
a���W}�|�O֥��w��_%��*����_�׺9�\���"�8 <#*h�}_�y;�V��)1-�]�k�8���,{i�e�$F�rZVNe�~=7�Fa��R�5��P]��Q���Y�Q�����Ų�ê��r���l��@�i~8~I\�K���7<B�M4�%��R�s���!�p/���*s��
��@�r���R�zl}��ٯ/>���_�����(�^.�� ��_U�J�����ECEY8���u��1���d">�B���_2��a=p����
OSs�i/�vy��7fi�L�.^���RM����fSe�l�2H&6W<n<k���l��$(�=�U�&{���WKϾr`�Ge��,���ϼ|_e�6��2j?��f���4�����j<����������3�M6�"��d��%�����AU�ϟ{8��e����^�6//Fe\"K�?��0L�i<fY�h�GGG ���f�Eea������׷]g����;�&�5I�,�j�S��3۬����Cui�_�³Sz�¿��eYMц0CUi��O�ARJ��ʼ@�vS�$_��5]1s�~)���8Ƴ ���Y�����_^D�y�=�%=��O^J����m��e�6����g���KqY`}�̼��$�2����% l3UJ�)61.eZ}�)����a6N�"��s¨��~N������ũ��%�b�>�uʦ.�W�w��p0�0���Lݾ�'I�v�Ѩl�����>���۷k��L�\I��yd�r\Eby����{��2��l�ϭ<��0��_uІhP��+Ҕ�Vr�8�����zY1�R��Xկi���w/�f��f�Y8�K���~��\���H�{1;cs!իP�h�O\�!�s����l�(B�eq��e��5c�ȌK2�kf�*��*J&
����Oװf��qC	������Lqm\F����~֠�,���^��HM[LI�i\|��~P��Z=�����u];+��^7������������?F�4�Ү[Yf2��s��l\��������uTjD	�\�(�-�,�y�K��`[-z+c4MQ�F4�����` F��Ĳ݊xF樌�!�<ɋ����3L?ӚL) �o\�<����m�����Zf�+5c�Y�	�Zs�e��r	�mN�˯�Ƞ[6g;^�2G�s!��}K.��EAj�9p,��|[�PɸD�G�K�s�u��������Іmڄ�3�0���rZ͚�.���r�ߪ.��T�_v1[�Y(YAx
q�\��x���5�D`;�ۤ�j��U"�@����ZZ<99)�Å��fM`Yޝ�>ïI��`�n��m��è�������`�rrB������jR-�l�1`wdR����l?X����������P�C�#΂�.(���Q<��d8�e�NH�:�8/Et�����m�9�?��b^���v�/��.Xy���m��~������]ƨ<-��/ՙ�����Ƌ��מ�r�
}��s~��r�O���V=���K#Ǘ�̵5������( ���N"MI��!��!n���a�a���$��`�s��K�/���V�LB1���B�F�����,���+-�� �E$2k��(J�UH=��/�v�>o2�P�$�ǱlF�`��O�T_�&�&��1qW~ZZZ�lz�GJ��D���R�� ���f�x�x<F5t�NE�]
2�����u�C��κ±e��8�rl,��d�e�R�T{UP��Ѭ�Gu��*��x�`��������&��j(4�1��*l��@���V�U�	'�5��i�����#�2�_�OFc��x#LM�
MS��,Ѝ�%4%�����L�#�+#(�w��\�0vW}�+�v\Λ+-K�� �yD�ĝ��U�#i����2Cy�&���a��'ҵd�GG��)A{u=�T�U��^�R����;̅V���H�� ysM���\���
��R��U��%0����35�3xwf����b_�0\����^�yc�/�}��ǉ�~|h�[��7���̨������v�'�H�@�P@���N������E\B�;b-�E�P%��$���|*���)~��D]��j�0�Iu�]Թq�FP�����lԚ����4ϗ������2DX��jc$�?lZ[[����*K<��c[Xh3�����|ɖ� ��*���R	�q���^!��w�:V���_'Q����O 1X��;;g�P���<}�����������h�ɓ'��p$��'�"��v�I(�
�#k�1`�x-�&���A/�Y��׮]C�VY�	�,+�I5������,���s�3�$=��K�ٖA����LE6���s�9��SDN�	Q/�7*+,K�D��	�p�F�-�3�1����+k�'�{!�Q0�Z#%��Q��{�{*�����!�a)2��[�],;��PM=�h�V���� �j���ml\y��q8��F�N�&{b�V����ٞ�g�ߠMl���K���x���N�#�������_��~���i��[�֧^o�,L���U���|F�v�/����7,s���K������y��@�QEID�NZ�L0Jn>.!~9Nby^���,�Uy;�^�Jb��%������m<9<<�O�f����� \�iȫ����`RUN���X>Fg{A�q6��V��(��x]��dҟD�ղ��������Dn�m8~oT6ͥ�UL�3�ze��Uk,,Y��x0���r�
�t��B���Ǹ�+��|x���fsq��f3�-@:�k��E�]E���w�Ν���l�l��N���F���4E��{���}��:�Q���5��60q �I�,�Z@��f ��bX����s��cs:�v4����:꟭�H�JFX����������j���Voy5gy�^�)ь_��>�G�ӾP�˞W��d<9*�q�3�EE��׶�`��z#,���:PF�������<����X�.��y�p8%��4��蟞lo?ʢ�{ｷ��zޛ�G���Pb�� �,e�ab�/X[�©�* ��7ߜLp��k�u��=������6�m��&C��ʪǙmDy�����a�u��^o��۷P���|���>��j�a�x���\Nk
���8;呯�,a��w������p6��P0rT��GS?���xB�>��WS�I������$���ڡ]\)G��p`^�9��w��L��e���dBĐh�#�
�(b
U(o�AǗ�HPE�&������� �W���h8���������_���T0�^徿(2�0�5���կ���}P O��, ��I�4��I���ZU����h�`��k�� ""aȄ7s�W������� x��� ؋d5��*� ��X����ˋx�S�@�"���}�k���Q�q]|�d���l����u�K!8�0�h��$y����IΣ���
�<�L����%�cF��D1`7b�������a�0/��r��/�ݥq�T��:Ɨ�9xr%��T��N�$)�(��s�>�4���N�ٻ,%���X��u&o���4��~��ð�I(|�d�Æ�V������0��ڍ�-�c �/Xy�c�)ڏ5�!O���I."��mm}S�ے-�~�ӟ�A#�|� �A��?`���.f����L?��3�qE������,��w)�!Hwa��q�)S²`��QQ��L�C�~�����=|bw�o��d�>ӵ��?ϩ�_g��W�7����� �ƳgSk���i��r��!����@�4��'@Ճp��PS�p���7���t� ���n9��؁m�텕��>?��U��x�X��'{縺����x�p����GQ��Faj��퍻Z|G��M̱wx��z������$Y��w:<G�`�Y\��Nz���x��G8�hTac��s�n	c;�Lȋt�`�Q<z�#�A��O-����ǣ�l0>Fp��D!�	���z���@Y8lRe�����mpWhmv�3�*�G-���������}�H�o��5�;����i�*P��@���>�;<�a��:X��K@�u��I\���#C�5��7n��q�xW6��i�"U�j���;m�i�͔�԰��xhyuLf�|����a�$�F"?���%��t��z,�x��sxZX^VZqa���tG0�+W��{�r
 ��&z�L+"�ZZ�$$G�$��� [1�������dN�����bU�b��6�Ɠ�CR0�[;>�dE	4�OoݺUk6?��/��4�lb���Slbŝ(o/�Xn��e>�M���i�s�(��Y�
�pt��� �߯��"�*`����F�sz�#���lll����	;�ܮ�$�oU���� ��<XSo� TH1x^���D$��E2m�zU�������:�z�7��ef��y����HЙ!70�R��i@v<�2���y�m\TP�h��l�v{�����]��`��~�쫪c���*:m�X��$�0*@F tjML�b�Va��Pv �ϥ��{����׿���'4Q:�VGi��� ���d��\ԞJ��!zw]�l�Љ@�aj��R�@���z`<i8>��kT ��Q	��Y�*צd��/e$�b�hley| �ՙe�b�8A,:B-�܊�C����$���P39��h��~�N�m4���Y`�X1|e��R�Tn�%:B��gRd�
��e	ˈb�1Z�GG$x���t@��	���͎��:��Q3�5��-&?����1�ފCUP���(J�`lKK��pj��J{�q�]���"ԣ�)�i��RG��&T�cj�h���Z\�`#�w�bR�*�j�즚)�eA�SdS�
)}� 1�^����Ц���7�L\�ʸ�j
C�y$�Gbb���,l7�8T�����8�#�˙�yP)�þ�g<o�2/__~|h�k���%J�FK�Z}�`8߄JR�qN�IZ�>�m]�������GO�<�(ǹ�ţ���E.a�(cқ��l �E���=}��,eE��4/�;w�( )K��˴����QP0�{�+�K��o\�~P��@t����B��&"�@��P��� ����x�k������U%�$��f�a��^kX����v�v�w���p4q�Ķ���+�o�ڝE����c�����++�s�e��W��y��0�C'-*߱�P���jM�Ӧ�s���H`*��j��M����Y��no\���t�ce��(��0N����p�UjR�dX����2�VCu���\d�UY5��W�'Y�c�m�)��,�4��Z}8�C��9���ǘ	찌�+�������#&��S�b�:	�Uq6�R�da��V��'E���LB�Pٶ��I?�I�>�]��,��i/��w��8\Z^61I���P�c����#�
�M&�0��b���7��}a�-Z�	�Ŏg�e������� �:Z�n�;I��GC�tgg����Q0�0K�"�98��j�D�j�:�T�'�'.�8��Ty�튅^дݚ�¢v(������q�(���E��j��Z8I�=�:Ƶ�,��q����z�d�g�ঀ	A�����Z���aM�c1Dw4�C|����[��m���Z��1����|���YҰ�h�/IV���H ��~��1�Y��Ops@u�\*\	�^�q?֩ QLr�Q�M�%��9o��x/���Ѣ�&�P(�¯����#qYh�p�0p0�� f�:Ŵ1AR�$���6��:诖3ė!@�a����Ļh��D�~mi�ZaR$-����'4�Ļ��4�"�C�_A�*+k`H�\¼ �)�0T������oHK*�uT�y��)}Mۄ��5K�Q��{�-��Gק���Jr'��G���:eX���Px/�BS�U h���y�&i|���@�"Cm��]��l��zbUq`?~������v(�^���@Y�,b��pH�)���E�w�}W�6�����qR�����]��a^�8i|
Q���i�դ�������n�>���D$���EA�ixfԐLD�p�����y ��Q�$�(ӧ�"gS���"��P�Pv�j�h�s0�_���&�\<_�zd�0ܾO~�!�ܸqǒ43��\�Q�i�y�oQ~�h���7Sצi|�i�|�T�+R]"�ɢ���!(�1e#I�Xi���a
p��&n)�O���Mp{����������[ߺ���}zz�k	r��lmn]s<g-,-w���hOB��M3���c�|7��ul@VGHq!0b���F���ѱx*`BE�n�[�f�F���|qe�^s�Oz�)H.K��i��_	qaJ�fQ���;��0/Ϫ�Z�`������g�>}�P ��iR$��	We���.�p��̔�7h�*�0�7p���&J�3ľ�����0��	=�uU5�5:7ġ(Eˬb�\-CP��ؓ0q����0�����խ- ��D,_�,IZP���GС���jk�+������'�xqs��,v�����N�֗���'�ݳ�V�a�k��o�ľ`��sl5D6����'��og�Y���잞 aܾ}���M����6"ODbӪה[�ZM�YE�i�@��>�������Ǣ*_^Xܸ�ڪ˝v��F���Dx�e�8H��i	���0-lM��&���l�18�"pS)���:ʑ��W�B�s���+�f�Dy����Y'�pk�*�T,�bgo�{5��댝����f��i�I��']�`�n5�D�S�5�M��֝�XC�p�b���@ՠ�;.Ѕ�K�*+S����eno�`���c���+�Ov���jmu��==8>���jwWm�Z�ʪ�$���8x����%$�X�JǼ�uٍ�G\~�høl�����TH\�ʱeYʪ0���X�'(�?>;׭�"A'�/ᄲ�L�)5�$텖�����
g'�F	�ܨ���@
@�&% 6qU�$�y;�g����=��<��|N�yF�Z"��4����|���p���D���S�_��`�.�ժgL�9�E!�L���p[��Ŀ���F��.<:¤0C5@4ס1�1��~ cIE�'5���
��S�|��]�-��E3
 %I���H�,B���42Gt( 1�3(����h�#�$���ʠց�w�0�'�1I�F�	6�btԜ�dѰ�o������'�|r��5JK�>7bۘFzh��K�6�mQ��1�#|g�A@R4R���ק�~JwQar(`
'��
7�.0w4E%
N#��T"c:}:���$��@�<i$ꩽ�V���z��CNNx�"{뭷���u!e�_����C�|,FH��JU#a2!""��Z�2�$�#ƀ�c0�s`U	!����0w��Q�F���pW�R<�-�Y��!�C��G1;�@S4�ֆ>V��;�Rge�]O���@;��/z��(Qȏm�e���,���۲�"�w;��O!�P�-��-�Zoi��7��Lⳳ����3���_ߺY�6�u�� ;AwC읲­5@�'�>ey|~���$�Lccs��q�(��u]YZ��zJ���,���,E�Z�Ą7�,��;�,t�	�y���Rv�g�,-�8ϱ��� �8b��AO�k��,������ώ�|�Zl�Bͣ�����^�re�լ�p#�<��4맧�([�@ k$6��V�=
�"�l��㱪�ھ��Y���: �H�EqQ�ƾ,��U�^e8�s��"��p"I�j\�ILcP�q�U-��v|x��8����\~�F ��o���b+և`5�E啵��X�iC���=:R:NWV���|p.&��R��ą>� K�	UE�Xb��ơc;{����k[�>h4ąM��3��EtϦU�r����"{
^��P�-ۢvF���l�����0�����{O�ٲBpdU��m�H���ŶR��V흷�q�ll{!i�35�A/��t�
Q��sL& �A��d�G{�A��L}�z �
������'���l���'�E�] �Ѱ��N�$GRP�D!V?D�kk��x\/E�����,#�����^ ��]�^��LB9/�+�mJ���!-��N�#qbW�-�� ���_��B��j����V�vJ�s`_P'�Cbk��x��{�������J���ö��2�!Tc?b��ǅ6T���C�IbwJ���}�y�1X!EHߣ�1.����}q�!���2 �H���ww)��Eb��F�I(�ɴ�u�L:����0�N'AMA���XA�HqB�p|g���e��y���JJ�;i�O`|�
��u!�(���bG5Qʌ+��W���W�a4ES4�[��i����� �L�*�� |����ǫ�� ��գ��{X�O�*���4
�L<�J94����zMX7�� �^ �7������ L�]9J�4^(�[r�"�����1��"����
� ��`h	]`�hǥ�7rм��b؃jo��6�jd(1<*oHh0���YA��]�w����-�����.�$S̋�T7�uCY�.�3�5�4�G=~�7	MoQ�޽{!MΨ���a��[��Zk�W����rQ�V�Qa�(;����j�E�+�2�\O��4���6�u��T
�g 2yT�qR����Kn�bіű�\��Gc��b^�aH�.�C���0����۷o��~��1�A�gO�:���Q���|΢�jܳ)4��9?ƈ�?�Q=�W�"l�`��(�ʩ��z��n���+�8�rO0����E�(n������i7�5q�Nq�A�����;H������c�x�5����?��Op�q|ϻ]\���q�U�y��j[�u�$-���,-2��DbX��NQ�H���)Z��-����az��ؚ��S�W$<x��H۴Yc�<��=ǭ��]L}�<y
���yE�٪���E �zI^�-WW� �0�Y�:h�bct��(�)1;ƱH�ԝF�sL5��Fi����XmX�����f�No�[x��q�WWWQ��l���Ա������]���~]W����������fTt�-�YP��O���I����O��&�s�tO�H�n`z�Vs���d"�4�WW(���"YZ����	��n?~�]z���T�i��������ZC ����2�2+�*���h��tǧgQ�,.-u{=������b������Q<��\6���S�:	��\�Q��v3�y �U���ZO{��1��0Y��ć,,,��~������_�������9�9�B?��G��C�(�%�����$YZM$�瘈���JҬ&�O��a�S4��+kk����B�((�Y��H�g����;Ti^Mn6p�ku���WT�FPZ�ӳ��q��?���ƍ��+�3{|�Ӥ�8���h���A�*�"\Y�H����DAn������h�2�(/Jy~�{�Ȭ�"���i�"�R�@���}L�wv���D1�J
�5x_`$��j�djL7�5;t[šǝ���x�� zpIvvv�z�Io�&�����n	H����E:K3��/�����9ͽP�ЀQ�4 4����쌶Ҍ�[�Σ�N�-��"ähm�F'tz��F�2��+S�i�q��1a4��a�������kG�� �P����S�ݑ�5�q�1���C�[< ���W�� *%��dµ]�R�9=}��젡4�6/gFS?���02L�6na�www���
n�0�]dL�=�V��PE���Ғ�L��3ޔ$�$��F�FE,����Ņ�
��86�����2b��t�3T|o����[����ZщSu��$�%Ѻ�|A$��d]�-���#f'v-QtlxM����/��(�V������!1̥&[GT����E�$���C����dI���U�{_�jk(�#��������[���B�����𻛷n��԰�DN�~�O0;7�~�l���-�x��EJ�ٗ���`��xiQ���\< #�;B*-��G�<Q~�ĭܸ�%*S����Siv������u@���]@���y������d�`4Y�k��wB�-/�~��\�5d8»8� WU����_Ա�
���U�f?�# _U� r��gg''g��/Y&b��h�f��9H���?�q�
\�I��Q�ffQ:�U3*1}��z��g�MK��Š&��������~�q����$^Y^�,w6ED�]�T�jT!�`�ֈ�DA��� �ɰ��(��P�E��#[$]~m������F���H<�M�M5u�?#�i')�/,.����Y� (��pwW�?��/oݼ9򼿷����\�&uO��~p���E��G��0��R�;�em��u�j��F��'��sLd�6Zm S�0/e/-�d��]�IP
���?x�hu
��'���db<�Ѥ�q QP�����|�Y��Mq̐h�j��jdf�~`�a"hүٮ��B��1Hu�����͎���(�Ƒai�D��N66��D���A�� �d.ya�Ǿ��1���]PGR&jLQo6P��8��4L{<	�E���&���I�&�@�����3��)����� ���S-G!���z���X�Ƶ@D���d8U��(3_P���b��&��d��m���,��(������yH�Υ+�Ď�4Dj��Y~�f �~����,,����/�Q4�-סc&錚/t�����/,��v0S�[Ϧ�����m<hp��B�`���(0(�.@�����U@��۷Aw���H�ը�#H�>=n2ч�͝;w%�4���S��GdM�Ӓ�16���:Ú���gI���$�h{�����Ecyx���!%�<�t�eo̘��i��8m]��1����wg�� ��pj�oeuI�O�)4�p��\Sj�%6A*0ʲ�o�_�M��>�R���Uw��V ��O%XɄ�!��hK���S�����#J�������i�rTծ��	�����1wZ������d`XimE�AayQO4���Vjd�@E��k��e�������21�ɨ�C�����F}��웼�'8�e�i����#�l5$H����u' g7�_ch)J텩����� qni5��q<�@��]o4�O���"��g;	����(�����%�)�"P�]��bj\m�
$�>��NIČ#��a���^��`vdb�{��C]�0gg]���P6���t��$���PD��mY��g+���c1QQ+;����������W�}��7���-������,-�w��Ə��rh�[ĵ6&�BF��є�R]7H�ʨF��z4�0����ݓXk�%��Aogg��L|���j�+ת���֕����U� �TY��=���;� MF�?���]o�=P� ���?���}���1��щk�z��G'��Q�8ad8�4�?��V�\�y��'�|���Ju�BL˂h�<�՛ iEGW�^��XV�]������v�[n��L�+O��͕��j�?�n��<+�
#{ Y;���7o�;���-����"�ʋ��{G����J���6�i�B�:� �s썭��bay��`ԙh�>%'�q��L��35ǵ�<�����X���<��������\{4�D�(sA#�Ƨ�gx�W���<ǚ���DY�TPu��?P�����}���7����㏣��
���A-��W�+� K�"�5�`'{����%Ѹ^���vgaks}0����㊐�ȫ�b$�K����ӧO�����Y_b]\gR���H�O��L�۰�rue����}�7�\��z�1��l�	��Օ�2���,ڽ;w1��Qn�i*Άfu�`�� ,����.E!���N-���M��iּ(�>P��<�ʋܹu�6�C��F�(�dy���늙��s%�0�%�N.��^{q��b���ᴨ��TX�O�ޠ�3m7[��^�}C�����A�s`e~ww7�DVo	�V��xS��q/J�ZLB�cC�� ��_��J�lt���d$�뇿�8~+����95�t>��c�6n�^��cPD�ã���+k�˫�"4�*+ɓ{��e~������e��~6��,��,g��7O��!�p�NOľH%5py�?��#����Ν�@� ڋ4�{�.(M\�?��6�<���D�a�PI�K>�?������w����7�LH��/haLq1�L�[���i�XY�$�B���v�*EV�A�H�P��on^����z�\�����_4����F��A�v�Q�ߑ�E��	"��=;g����H��p3��h7��msKzi�:?��ς�>cX�P�8�Ja<.�m%ǃJL@U�cmIҒ��Z�*�-�*�Ë�z@zE��_h=�͋����s<�~aK+�X^��kk�tS�O���T\��y2�ù���f�
r���n:��IJ�P5�-,2 �Sp�pX�p\�<`��($���9��%l[Hr��o6��Q�2��*���`��ӟ~�������6;-� ���A�W�^22�pʂe���Ҫh���E�!��c�:�D����+�6)ͷ���e֖�8M��t����0\U_¯��q.*7���A����X�AW<�3M�"�꜏�c`cT�!���	:]^^d$2IT���}1��2u)л�t4����:� �hx�]�nJ�����Xÿ����A���hc��h4�h��Gnl^gHA��h��bٽ凌6t#�K[5�1��Sϕx�T!2�0��SS�[�%l��G�������L��^QH�2��O?�g1R�& ��``	jM����Q���ަ��-!�4|���=��PZE�O�Q\���u��K0�
�U��y��DS�T��u��ϕN4$xvu�nI���Ǐ�b���y_�!�ē�G�D����oa
��ƁB ��V w@n��ҭl
���Ķ�fE~|zRW')jw�z�]�����CN���bj� $��
G��۪�|�g�Q?x��s}OH���Ң�Pfi~ec�&@���8���TPt�,9p%nd"�hR�J�%�\���ĲA�w�Nc\�Ls�Z�z��ʕz�O�N�H�k"1C9:Ql�YO�c�� ����&c�ڻd���Ws�%G�ǒ��	d�tp ����d`�|$�ΰ2�[#6ٖ�xt�$d�H�G5�(z�,y�-F���,ǦŰ�3�>��+Q���<�+%�ʴ�n�N�!����1|=��0�t�o5[~�!A�՝S�����'�B�{��4[jw6V׀6����=��7�r�:@9 �#	�&ю'QHc����_U�p�ȡ���Z8�%C{b�,
�����G�đ�&��D�+ok�`����S��z��j�}[���}��f�}Az�����׿�����;w��8����q��g�����|����C1�)�r
�����뇌6���	�$�F!J����N��t�� �J�8�7n�R��'��(EŁ�w͟�5�EԔ�ҟBRp�Z��pϷ��iɃv��&0�^�'.�%y^s@.����3�ˠ!�{ ^"9������W�TF�"C凨�j5q-����ƚ�Mc��5E4��J���"�++bD������.:�J(�q8���B?�*,��L	ֱ���MaH�>��<I�	C���16���Ƃ���^����
V�Eʡ���2
�
��ƙ�����`(�Lu����H1@,Z��	5"� =��)��Q8&7@��v]$/�Y��2^_]#Ĝ��h6��o��-xqf˄u�J	� ��?Ui2#�ƀjt~V�:���`����b��j�LG{q�P�).��#\i.�yuMh%�h�İ�9���Y�S:$��&������o#W���"�s�\2?����T�p�,�K?]Oc
��Z��(�F��O�ȫЏ6�4^��9 l7��g�:��1.��4��NQh��XS�S���&�,��	�0\1��k��q��ok�����{���)Z�+F.BZM����^�//ɀ�<H�^f2��z=T�? ����]�X����&��X�����>��$J��A�sz>��?���5�� �'9(�p�����{]!��I��H��S��W�D���Q��Y�Y*�4�*B�@ (�'���wj�hӚ��B���X3&�(H0�NАH� �8� U�H�Nb��������ƓNg����Y<:�mCeh��)��%1s<5��]����4�g�g	��ӧO�#���"s-��V����p8�CY�"v�3͆���qg��$�x���"�������������Ç�iqvr:��zt��$�|� ���"�|"!q�; om�Y��\���"��;���u�wyQ��hK�D
�L�' ������o�#f3>��U��qT������X\��E�]�fYX�$�4��z����@q$�o{�����" ð1�^�OQ��� 64�e�J�F ��s�4Y���Cp�'�Y�X j��@�{TM5ϴ��*�b&�A�fU�S0� :�ϞF�4�~o<���g�"�	��4���=����k�m3{�q)�8v^d�0>>9���ʕ߯���I��5� a���bq/I�oܺ�!�b#�+�+)���-M�eb��.`r�<���E���"�L�nK�żL�*tE��n������4��n ���\J�ڵ�B~���?����Gؾ��o��o~���O~���X�z]ٟ�<�G 2��T��%B�i��GR�@ߤ\�+�  �N��q<x� ��u��X�D$Z����:�ޞ�V�|�0y��Up8� ��1�%-�I@��	�4��Q��ɔ �dh�fC�4�٣G��YL� Pp��z�),��������Ы_PAd��h��48}�Č]RQAP���H�Q�/Tÿ�*�1A�߻{w C%��1����1.$�y��}Ǳ4�A|1O҅�Y�K�ғ!3.l�f�ʣiO���Ti�u���\p��lHljSi��n(,�=����^d����ÃJT4���.cʨI�#��ȟa�L�K4�U�C�?��}��l���fC�rQ>%i�$�TY��݀�G��D����
+��@�|g�.�s��_c�`[��|AS̤��Hlve��C!�{��`D�0��G�SƔ� �C�%�,�<6�]�:�Q�C&�ub�vC� �0�~�Q���x�����B��x��a�[-ZO�)L�Iű5̱�P`����IpM�B/]6�&�Ub��Y�0i5#�0��漬��ʧ�ov������%7I��M(�"s��1���'O��:�I�/��/���D��ƍ"�+d�1w*,L���MT�J��o��%0�1M�W)�g]1�O�@���Ҽ�ฏ�`������9���ͫ����n<)l�p�e���Z�'��iIt~\�)�%@mii���~���A�
�-h" D��kr��Kr�6�X�x��7�FE����u��V�ODOH�c�^��xx �E5���I�j,¢:����om�����4�*�q'W76Q���Xb����^����8��O$*��b����p)���4��C�^�R0LE��1�<�7�1 �1Rց�bJ�f�AQ~=>>���^�u ��N��O�����!��0�����n�y ��CkҖA]:r��爢�?]Z\9����M�D3��8�"?:�ꀳ���B@�
X�(�	��:	ާ�_ P�4rl � `$��� �!�ڶ���L<���" I �<�~P�7��0�Q$߉3,2@�ҩi"�Ɩ�q�Y,q(� x"����Z7�8TP�A��%�J�nyVYf^���b-Z`ʩ��9��ְ-Ƈ�I�{�;y��
�$���_ۺ�lK�K�K�s$�}�{xt��l���Ŋ��[#8��hc���bm'ZbM�KCC�R�����F��"���z��c��i��ǻW7%:rwJ��T��g
VN��lϯ����s�0�H��w��������������?�}�$g����CL��M�D�4z�����5�����&�RͅT�@��nʨpr$E_D8� 4�F���������m�@���m�rM�%]P�S�Jt�u�DCLLF5/�g�*�d��|y���;4������CU����,R<J/������4hD,y��uWt��C�(���&�U��c�#�����Xm"��`4 w���͛ 1�LF�@)<u$�������j]��(C�=
�rͯЦ͌��(��8�Q��w\�t�uѴ���4q�80���=�1$��BpZ�UW�����/��K���hR3�.�����t	���:��<��ree���x�&�[�B�fm��g�%Do�/p!}_Z�Y=	�}$i9:��&p^�J/�:�O���ľT�%�����>���3�P�� c�>-������$��y`�[	���*4�.�8���PW�Y�C,i�g��G��D�x��ݻ�i����������&����4� eIv�ߥ2J
yhف�� ~�޽{��k,^�P��i�QK���,)��a�����~�tga�+<�I�RI4�??�%�|���)��Bw�4�ts��R!�$}�?1cXb�I��vK�i�'�lUay���'h߉�/[W�2؎�ݽ��~{��:������Ō��x�+�6�fYy�.�0��鷭4���L�$������ށ$ˬ�;�>�%�yoxv><���8U����u���Y��3��W :�-�ʤ�H��Pd�g^c8��z˨����#��{����T����B2����q<@'���|��v��x�7p�?�.���YOL~�O?��e��%�fKcq;���*�x��T�Ah�k4kY��Y��������4E����ju!�����#�#���JҺ����8?�41h�LB��x���a�ҡE,�@	;���V1P�"..9�N���`Hep���O$�a?V�߂R��0N,����v�>O4X[�s��)�{�0��P�T4[L�����<9�Q���җB���9�+*�#*^�A^Z��t���u����"5�����t���s����.�C�����[�	�#�VWo\�� !�1�c�Qt�)b�M2O8�8$8iT�o?z,�EW��Q�ڎ�a�0��C�b��J4Kkv��x��U�H[ӳ�����$�n�����Lc�`������n^���^G8�����@sG�?������d�Xa��?����Pnݺ�>T�E|g.�c��W;Xq�-K'�� ������s:æ��쁌@_����17Y@☽�߂)X^Ya5��z��rEp��;"��7�z��qw��R��e��G}��i�7�x�w�2���T>]��5
'�^�N�_��*�H!������Q^9��UeJ�Py�8�(�&���zO||����y��	�h����>	pR�h�J�׵/l(� �++�;-l��\@9N@�X���i���H}Y۔����h������.PN���#2
	�V)�ѮF�`T%@g�0B�gS����+�7�|cCw ��Ԁ<�ܫ)�3��h�%���H�fQƔq{Y0��{d�I��?N����64~}�� }�y�I�f��!�$:�zS�c��rх�z�S��N�tq������V����� :��ښ[R~v��:W�|�vM�c�%C�5��d2-�P��j��3�Mr�'�|�֮�*M���(�d]F�I��5�^�N�2b��ˁ����	 "Z�ƃU����d��@��ո��ɣE}	�-	,b+�f�=\,5=�2��n��l��2��	(+�4݈�6�����Q��pK<$�Y�j{�	c���"z`d��]>;9e�%b>rc�	Ǣ��$J�,��-/m��l�R�\������ȏ�tj4�d� ��G�z���,�?U+���y&֤�{�S����\"O/��u�2X��X���l���o��o�S!���=�E��8q�����0�B���Y?4����fEN��4E0�� q�����ԡ�����/>< �r����U�j��՛
�@�1�y�N3�ɮ�)/!�*��QX�F'%)����]��̮J)���m=��<����st���f5T{���AB�e�dˤ�?~|tx�.n޸���P���0S�-�� ��F2U� ^��3h�%ԝ��V���G��@dh�Q���..VOCRg$�e�n`��+*a/M����4:���+*,���L�uc�TVP���Cq���m|�c���,!�G倍�F���<}�j��^� I1*ʵ(��V��b���M�qR)1*K��|���:(��.�b��{A�1-�0
˨/B?�E�����x�ݡ1fz��[��ux ��bp\20^w<�x<�J��iu:��0N"�^Z^Fw�ASjt���N�5ew�2�sܸ���Sđ�@~�z���$��E`G�T�>ཊ,
%��]Qkc4��&F�����"�S�P��qjV����8�@R*z�|q���� h �	�|2��4γ{wn�������V�O4����*�$p���\Y����Iw����~��<϶&�b8:����e�7M30/�`v�5e}&c�5͡��k[W�(�w�H�l7��ȯ��@�>[��a��V3Ӱhz�F�JI;j�xcg����_N�yӬ��e�v,>�8�'O�b`��`�K�������6f
��c	���Q�V� j �818y��կ>��3&R��&�ð�t��ꂠ��=��j���n�(T~�'QA�v�N3W,�t�o��vY=\�w�y7GC�.?|��I�h���O�GK�/���P_�̈XT��q}�By	�����������񌋴z�N��QC�"�,��-9���y1�N3[~��%�NPKN�
�)�`�Rt����Fwx�a"�--�9uԔ��g�:s*?�\; ����K����H뭷�̥��}�%���F,�i&]�HG�G�T�@����� �L��/�ͩ��5�ϱw`�T
t`��`!�|U��8t����@���]���e��s$���~ݻ;O	g�u�(���<n޼I�niM׊�><U��k��b���HD %ɩ�a�&^��B� ���c���,N��h���PqY�-��0��k77��S��Mu��u%�? 1� V�e����׷x��S�芵:51�h�+����-�f�d@�Yڞ��gD}t$ٛ��6K�y���?�땵U�.څO��߅rl-X�p�`c�;m2XdG$��#��T��d"gui�����7����qkc��M��W7����dS�-z6f����"�9�A�\#J�����q������~����8�o�m���$Lp"A��ߧO����B�]��7+*!K �4+�r}mC�=G�i�88L8��4�n�Tt�����G�H�7��̿����#� zp�����n�ȻO�n���M1������&ݚ�}�D��!z�<��)M�ݧ�����L������ʹM� =Ej���DȜRN���h �2'���20�i兰t����Y)i��31|�|5��H|X��G��ivx�d�՜��~�/~m-�3D��"��IJy��%�)8�R�Wj2Z��I-��p�u��fV(`�k�n��g?q��o?������@\���U�'
�FC46�y��-��Hu�� �]��Z��N&e&G.�'j��ͽtx&?w�~Lq��1[�xr<��\^[�y:�n��U��`��)�4���U�+@% �/�����2�!�.���������`�����H�hl�5PH�'Gد������:��;.ةIY��O=�ƞ#zo�:e�\|>��*�� $ww!��סY��R�������
�/�Ť��Z^\<;9��E�ɠ�;��!��͛c�~���}	�_k6n�7q���\ɾ�DH+�bkk���`2fԼ�`��.--�����-��������U�qv���A'��k��&��L*���[j4g�+�Ht�Pg�~M$���������J�:�5�-�Yj�ͩՖeׂ�㈀�ȍ��ީ$������+�����t���cA��q=�|"�����\H��-�%�|���>���uܽ�D��Bb�ol� H��O-)Z�Ӏ
`]�JK���.�Kp�v�̇�����)�X ��П��1M�cR�l{{��
A��wq�9�ڧ�:$� /Ҫ��e��73G!�-0��ø�TV�.&L�W��b��F��5�f�I�֠<M`��Q�1�VO�.��P����m�Ţ�c^H:B��&}*pդ
C�U(J�9ʋJ�i��X�0���	�X�b<�����ڮ�Ѥ(�����Q���tb����E�3@-�$﶐��|��zQ�3W!������5D3��2ʽ���v�!~�I��3��v-����O>��ŁfOLz�\J��/a��"�d�f���l�2��R�cc�4��H������HY4��hiiM�d�q�kBAB+���hH��ҼLT�/��D�8���N�b�OO�sP#� !�="�>3����خ�,5��q����5�)�g�|�G��c64R@�IA(O�\��NZ:`�uͤIߙ m<���P(�Ņ%z�S)�aŦ��U�!D� �"���Z<���W`�6@�,.��M��=���{�&���J�n�ys_j/,v��H��춻?̄���?9&b&�Y-�mY�DR&) ����3+�=��s�S������1D����}�g=�yzm��'�|��{܊��ۃ�bݞ"
؊�A�7���>�o��������#���VƱ![�$�<eg�z�j)�����l�;��/_��F:��O�}��X��x� �<M��L�@��B�cu�d{{��͛7n�(}��`�3�R�3H[ٞ�.3m�K�|X71&�ݻ��C���~'Cyi��1l!c8���g`2����ʂﲞh�Oa��"&DƓ��LFR d���zB�V2�Ju�Z\̭ewa=)��I0p0v6�g��21�e/bK��!�).�B?b��/ѩ����g�}6�o e^T�H]y�"���F�.>��(l���`����h����?��Oq&_Ӯ��X&��"�Ƃ�^�#.�L� ��v"W�O8�{�^�c�)7o���_B���~�f�p�Jic�Ӟ��Y<�Vi,��T������NV·��ɞ���*�����A�{�.�:��\j��Pu'�<���ML�0��}g`z��l����V��]�5�����Ր�bO*���b��z��\��51�v�Ĺ���^:��C�߿�9n.�/+G��ã�k�XoB����B6Hx���[�'���	:a2e	]^_�M��d!s�,q���CAu'��s�K��!|
KO��{���i��=N]�;lCt{�hJ�x�,2uZ�����1ix.]�,-��������N�S�h8.��30K�1�3���;�woݺ����Ŏ��\Z����j<�Dp����ϷS�|�����?̣j�Ջ�K�U���5*������¿��[���֐��}a/���k)O���T���F��ӎ$�,>\�����!��D�A��YyU�(4�Xs�����_<x�@�R�x{�4�7�8��ѐ�v����W����	Q=i+
a{K���>=�s B-6v����;H:8�!͋T�>36��hʻ��R=0���s0Bl\@�{-���nD��ǚO��+j�X+U�������i6,HB�q�P�r�H�2e�&��wt�_�JRm<��a�]��j_$=�7�T|O�.���:�c�����v����j	���:d���� F�uY��UFI�ׯ_�,-|��K����o˧Qy��dJwK��*Z<���3�DƝ;w�G�ie��R�x"lzF��st�ek��)�ʵ� fF�aE#��N�!崔d�����,�$.,�(�06 �W�X2qM^�zM��+$�9���R�K(����b�K���&
�Z[Yq�@�&���R~r��鈜z�W�;�E�I�@�|�S�Wm*e�E��+���\D�+H�fCgSJ�3��4�� WX�JA��Ю�M�6�(-���C໐NW.���{~A.r�LEf�A�2��Ϸc�-���Al���~,��N9�ϳ��X��{�>�G_$�|��wG�������4�q�Q�����������m6�]�qc�`iw}�Pʥs�0�H�OK��_��~g4J��F��|���+������v� '_���l4:�ϡ�ȇ�����3{�����d>p�Wd9E�����$�c����k�E�o�^U>�]�U�q��ryI�.L�#���`���͞�u���@�W,1ڰw@f��p:I��t���["�����Z>9>��'�{QX\Pdi�:�vϝ9�6�����I�K��Re���������ƣ&��'3�%���u�wv̦p*�A0Ǟ�n4t�l��˵�S���gB�4� }�MG���0��~�
��.Y �$�l>U(U�%7��y]m�J�"�x��
-��X�!��r"�d�:Ū4h9BEe�*|�O�tm���us��,�{�f���O`$��+�0�z�t���H�
���8<�7�$<ǏFѰ;���a+'�s1N����R�$.�m4�%v��G�Ѱ�8�}�z]ȸ�����cL���1m��,	7�܄�|�|8���hIoH�U^eV���%���WX`�y�϶vĜ���ި��f�'��UcO��IA��X&?1&��F=�j�ͤ-RK.>�s*�����f|�D]x#$�ZZY�rw�n�Q4lw�[^^�J��V�Of�0M��϶t.--`��I��a��n\YY�t�*)FF��~E���4ZM�]�0���"��d�����G6���n[(T�Ȉ(<Txo�X�b���gt�d"����b�Q�+�1tD�g��0t"hjN��V�`6q�Ȇ��-o�=�>>b�/��/:�����!|�^���b���uzN���>�Փ�YI�=/ɷ���v��������9/>�	���=Ctb�ǎ�I��i�=��#�C(FA�efB�D�G~�Q4Q�z;+B%�R+�}gg7w%ii�W��"�ق�ܣÞ "
�L�H�2������.������d؆F�##��K�	3p;ƾ�z���7�u��yVE�Vׇ�j�e�"�����`�]t��!_�CO�}�p�Lbύ/xy�'R٬EZpc�r��M�']��Y4HT�h�2���w٬�'d-!.]�ճ�c[U���3��bK�GQ�H��r�$�Q+�;��ǃ���
YQ��0-&1!�,R�P�I��<K�Y�w�eT�U�CT#˴��X��Hژ���d(L�A6��"y��إ*�����������^U�c��yY�J��%r��U�8V��A���'G*R���
/'��1(!����8B���$�`����{�h���T+|T��|�f�K��p�h��-�LT�G��b,�7�x�����\&�)�!E0��1�������6fcyyQ`
) yH
@iu0+��{a����t���^K�Ì11;�$z4���K�����4�;�wP��J>ȡ1��U��1��F5�`њH�P���{]�p~���7q�/^���{�r�L��%:Sj���8t���o��0-*����d��ÿ�3 y�u��� �:�5�_ia�lG�+�._����ちE�����JElPl���׫˄�;4Y=�=�av9��P v�{�2:�H�t�����-�^i&�Ew�5�d�[?�����e��`<��ّ�8��T]���ޏ���<�|B&e��q�1V/���=1;A.�2���$̿Z=y�r�Ƞz!�IM�q���s�֫�8{؂D�F��U�G7�K�li���}2%�]�.�Z۠/��q�jJ�I�j��H���a�3w2=�^%�%0BY���P�T�"��l�ﵻ?8g��YȂ�q�u�Dw��*HTC !
����H%�y8gI��Z��R.t���A����P�6D�����OXZ��6�1���_�2u�R>F�l�Y]`!,���U$�X��ĥJ9�	��	�Y�TI_�]�^1�I�P���@b�#�dN��+W.)���1x͹U!�(~u�����P'�d	���K�Kr��G,��Kr	��2u\�#�z��d��˃�����uet�q�m�Ol�)LDE�/A��>|�O�ϭ�L�}סK99�<U�ܠGn\����A�W����,/.�3�ÓSl38�2$X�#I, �T�83]H`�x�Uٮ@ۊ���夞�*8�{�5�.{�\G�R��<���$.�Uǧ�-��ž.>-��0�ڜy�k�ꈩusw;X��f��J����c�_�������c��b�dg�#x���U�~��� ��d:�
q����[�m�R��'���~q�v_���5�OX.����ׯ���?V�W�R,F5Q"�V���Q`/��"� �8�2�����Q��c����J�&�X���Yf��Pl]�Tl>�^1��ե��se��UZ8T�5�E�wV]'kH2��IV��o����r��p��]ܐ��ke��%�0�d�Du�&;B+>�5l�ʵ�%����
�`�*����b�����uCW%��� ��	�40"�f�U�F�Z�Is���H�[a�À�ѻC��&g`Y�hj���'$I�	C�;RZ�S3@s��@���{\������>�L�s��R�җ�XE�R2��Ed	�i�M�ޗ��`ux�!A�|dq�"�bUl�RVU �ǊCq�|��5O\^]����+���a�~�2m2ꕟӋ��F����R*�� Dݨ���L=�p����5�X��c��uI�!���X-��WT"�k4uXݜ�R�Y�Қ5��"�s�2�����KL��'s�'��f�����r6��ꫯZ��$�L�Z�ĵ�KJ�`uQ�$���}+��beA�9���~,�q���&񇝶p�*'DeoO��47�/g�'�*�*��!6��4R��P��T;%_��[:%���7�7�]����;��W��ս�l���l�ظ�L$�0� $����|������+�� bj�pC�Rf��?��?�ˇ�K+�tv���\���đ��������D �h4�_.��c����fGC2��5
��h�t������
��J0������5���>�8���y����2D�
QS���/��z��8�0<�|"�ҭ��0��
 ��ӱc�^,K��``�*�Ig��$ٛ��T�Y��2	�����a�����*���O�pi��(��
&�|������&�ozx@���k��}��%���̇t�0��(�3�	"Iy��G�ސ����K�
%ʥ��E6ޘe>noo+�(�rb͔T��0�Lr��Υ�8λ���TC7;�c�d��bh� [n��������x����,������\�iq�1��_�i����I�U�v��}V�G� �d�i2h}�2VW&�T�"�5�\�T���k��$I+��Z=_,(-�t��a��@�g�9��r6��DSx$�RQq$�,X�+�T1�	���`T
�9,obX�M_���qj�������H'�͕���Y���vyee��%���f��� �ż�� ��=r�I�E�AhD`Ƅ��յ%�+�F}rt�_���r}��fs��~�����&]ωf���)�l�Ӯ0&^8��Xv�[�o�3�
���F&Bc�:�|y���ؖ��յ55�R�aJd S�3�W��&��R�1D�A�!!����;��z^�%���ʒQX9�	1�C̤����Ig���r�Z���O�a>Lep�^�����l�2�n3��j��-��֩��I_z�/�KY�h��'�|���b���n6�f%�\N_DucK��$V��E���a�d�&�d"rCv��#�t�Y8��pL�P!��N*����#�Bc	`���Lu�E��*�k�Î�9��b�����1c��z:���o?�G�ݽ{�`?���lF8�b鶌r� d�P^
�R=Z#��Qe�p1ݵ>�&:r�[O3�&��ؔv/H��b��V�C��dr:��ź"{��@k���I���<Wƻ*�YQ�p��^x3c�o�lO��R}�bb�2*��M�,���#�y�Ν��z׋-�*��h\�a��oܸ��p�O?�T��b��ڵk��k�!(�CvU����Iī��jH�y����R-=^SwSI�8}%�a~�
D���us��������ű�!�EC�7�"�%��ӧO�E;6b`�
,�2�=��/�]%��9�(��]c)�a�q����u1�Uu��2ɕ����������!��<x��Q��/�S�2�u�,2��M�cN����T�(�KH�@5?�L�YR'����jie�a�À�	�omB�DWV�Q�֋0%ݣC*/M�p�jb�|T�$��R�:;Z�1�c�K�*l�"5������q���Pf��h�C�����ln�,��A�o��V��\I;;�Lv���I�h���/�T�54����Y�I���XT�a�~ú���[\^�@|�^�:��.�X	��,g��_����Xi���l<�\��` 5r0���͛��f�}&��\i�"�F��lW7����`��b�Uqvƕk
�x	H�%z��H&��i4�qj� �dy�o}vV�T��G
��l����p�M�����g�|���
�/����ӯƓJ_>�N�͓�����f>�P�^�2��@ಢ��(7��k���j�a��2i���G_=��f��q��	���jbcR�B�,%B�%�1�_Ŕ�E���~bΩ'E
Fq�Le/��<U����0DfNs�^(W�"�j� ��`}�8�mUA�fs֛�_�Ď�i7�|�,���K&B)	\F���/w_f06&�Go��f��a��\�����'C̞�CJ�omm�W� ��]�������5�I��l�HZm�[-�I�v�m ����dc#�n����aK,,,�jx�im2K�n6��(�݄FUB��5�N��F��BA{��AV*���e�P�79��a���0!�n�T����%\E�L���i�%v�� 8f�TƻE�� V��VF�� �l�qگ7�,�f2Oe���5�g&��$��t���s8Д�o�ƜCs0���&����%�
���f���v^����U���e,���}ωON������db;	��lw��a0�K-,���<��<�������i�޽;������67on�������Օ�Y<�n�2s�+���>�:o����X3ԇ_=!�s)��qxx$)��b:�e��:q
/�_bi�m{������s �c�P�e���$�$�oݺc��m�>cA�d�Ν;�Bp�����-�j��Ñ�Fp7x!Jl໙lh<���L��?����Yh��Y���[6��ʹf�٥�x�G�� jJA�1�5V�%l�6K��$���_��_�YF�1{�IV��>��]���$Oq#�y%��y_h�B�A���C��rc+�~9�Y__e����ɞUsyK�"�E�{A�%�C��ZR+IN}l��B��}��,`�ET�BU��
g ���w�u��
=��*_�0��*z����qj�[U�{ekK&��E*�_
;&B9yX�3��N�+�vA�0�����V�.zu�T;�'^�X`G�I��X�-e�]�v�}�
�[�d��%��ԭ��h����P���(!Ĥn�F��g@]R �(�Ɋj�R�J�4��Vڟ����Y�.�S��4�7�����T� �E���V3d@C��7-����1�%��P�"P$�a� )�9r6�Q*k��E�F8�򋐐�am�S��/_�N�6�D�U����̢rƓvn��
!a������LI����Pg����zlxhG1�(� 
"�F�����^�0)���8��~�{����~���;���7�6���qfs␧�O�n4�O��T>�ݗ�����1��@l��J_�v�b�8��L�Ҳ�z=�C�l��w�)$j"��q6�9��X�k76��jw�	�����d:����9L���GT�Y���aai9����0��s<7����@Uml@cu�<yU!;��"	�����4����K���y��]gת����zpJ��I�7K�<��Ic^\^ʗ����O�Μ���p����fH>�������P��;J��xb�$�l8��@��� 7{�}��k���I��.�O�L^�l�j��ǁ!�JQ���'�^?ch+�zɉ�i.��߿�Ӣ%�*��s��n��(���2h�:�tx|�l��@����t~��7�x���EW	h)��'O�T뺅\�l�䠊~�pP��z=a>
V�A�����>������DBZ�����,_���趄%�t.�k�''uI�uժܛ�%���m_&}��-C�l!st���oC�~��'S�������DPQ���9�W>������^Ǖĉ���4���������=�/��˅�|:OV��J���i�`
�C�E���X�K��w�0�8��6�-A�n���p<	/5�q��.7ll+���|�;pmh�%��k�6��7&��,~*Z4��oM!�G�	��EX��%p���X���	������FV���M�����{���8388ب��Rv=�*��uɫ6��!�68�R�9y4��{�V]�;�l�{4���e���gk��g؜�����8"S5<�Z���
!��NN��3�^����o��O��Op���h:�,�&-+>�Y���|��oLm`
5���?�Η�l��敷k�?��sh��	5�#�����/��b����������!�T �I`V����wp�"BY��}!� '������f xDj�V�oR/a�s}]�N��(x��V@f4!tJ�8(�Q��[^�����_�U07sD�(����� `m�Hw�����)5WS۽=ҩ���"�KM�-k�C��tH&��N(��c$�
�^�qj<���e�܎y)��E���jdݳ���b�Q&�:�6ԓI�LQ%����T�J�6�P��Y���܎�Y*B%��30�	��o	p)�,��(ܤxB�T��<�����-4��ￏ���_�J�1]�6��Q��X�a�4U*
��n�XDQfI�.��ֳm,�_�W��K 
%ܧ��"�0V��%����x
�
�����o~�,�&e�ga�#U_�|�*��V
M���خ]�6�;c�T��I�ۍy�������4������ �>!p�*A�.Z���X����/�D&f|n%y�����2R���Ұ6�iQ(�"�1�gX��
��#�ϚY�I!n݋�������er9f�\���	Ӯ6�l�j^�K�Ż�n�t'8��Y	;���6&B����29bMXU�նI�s��\K6�246�X��1r<���"]O�<�y�S�����8����1|�9��1�g����3�樁�����Oe?�98��bo90����0&C[�-�-�M��M�;� �D��������:��O���c5P�r)��a�Rٳ��pX�����Ӗ��c'��w�Ev��Zΐ��c�I��D*�xS%�u�łR��;�,rTDV(��{Nc0G0@tT:���R��A����g�Ήf�	%;��:���M�XP����1��D�7+'󙜚��(V[m���$��#��sm��K0�h1�s�j ᦦ�HI��P�1{Р�����0���a9X��p������*v&q�8�L	�ܻ��j9!�X�β�h<�\G��H'���N��x�T�bE���T,;
/n�(��kg���W�b��Y�r�I+B1G�y'�����x�=����ml�t�h���v�l�.�����5��>�S��s"ܾ�v��ۛ�aj�r�ɵe
�ӣ�;���.�4�FbIԙ�|�d��L����!�Q�kėJ�+�%�#P�^�V�2@e����"�;.���bi:b��ܾ};���G�c��=s\m ������c�
��7s��F[
���}6)s�#�	�#k�
��s�:�V�͊^B���ų���Ǔ ���GX�B��)1�`2�t�Z Q�Ю*R�0�����i+{������`�^�x���{���
�-�sL�\:L��)���΋��b&�eL{FBj��"h��frq4��$�0�;;�+����g��.`^m�O�B��%�=������1o#v�9N ���~��i`������B�$?a�!��䋲\��?��O"�/>X'��,V�k&�#1�S�4T[��Z45j[����c�0�Q�cޢ���$�bs�
y�qϭ�����2&��Z�At^�~���l�m?C)�09V�)#�&W�	�I�j��8�/L�M��76Й�S�Y~�P����2Y��m	7�w��V��<�ұ�X�5�glX-ƭ2�T]H�7�x���?v�ѷz8V�+�L�!n��f�/���W����6c�gl���j;�Qʝ͵��EiX�t��&Y���Pܿg����U���!��+ܑ`-��d�m���*�p~�=�˗/�/�+�V�^�4FX>��	L�/�Fc+�?(�,��(|w`��fk8�J,a�wE�M R9�E�@|BujF�������#XX�U��DU�g�q�<�v��R>��Y�n���� cu�Xcp2Lѽ{��2�3կ�ԙ�
զ-
����N����BGFy�r�J����◖ب��%?J�f���C�%� ;���"<X��D� ���aJ�h$�2�\�C,M�#I]�IS!�<c�d��Z�5�ׯ~mP]Ux�G����J�h����B��>�6�����ě�m8
���S+e��`(�+�3�ޥۧ;�1��Fh=�ږ��sBa+;��A��4�'>��S��?��E���m^�t恙o����D-�t[G)S�_�_c��;�P����biѸ�)�[�N*[2�h4q�T�F9���T| �5��/Ņ�@}�����<O���3v?�슦��տ^��N�mFx~ф�� \��w����_����� ;`���X�#5�f�oiG6��ۃ��7��W����ׯ���'�	E-\�N�߅C3NT^����I��o:�)5:�����|̕��|q2��ė�\��K8K�?�@�qs_<�{m=M��ZM�Xd29���t���,�C��b���Y	]2�������؊�W�F�KO�Z��>:h3;bɌ�E�"Vύ'�#]�y�99�@�]'�Ht��M���uב�ǋ�S1Y��D?�
�a>H�pZ�N2��N?L��kA4�K>��{��%#:N:�Ū`� �!)�5b���4����[��}�~U�����U��"0hh=W^��9s��������O�WX��1�����{�A������WVo^��۱H��)� ��O��(�{��i���L����v�U��`�Ƕ	�V�Cͤi8Ϣ��o�g��B�(������C�֍M�W�׍Kń��L[����>����?��_���b1a ���]��^�2xK�I��0`��S��'O�G�t�2�ǘ�X�iB�7�XI����u���V�,��T՚yznE�G_Ze~EǼ}υ U	'�aə���S�����bb6�r�2��ibAK��ˤvQ�^�#��2���!��C�;����,���"�r��Z
�G<R�:�|�����u���q�H�u�\s0�,���z��qe��/�*�R�0�f���/q��~��;�Yy4x���{���8U�^b��ѻ�����7��F:C���޿��_*?�:m�S�H�Ȫ5.�����T%��k��(@���XBib����I'Θ���`gc$��$c��XqY㡧V�)��I�5++k�P��۸|7�K,'&�TM��!F����k����F�2i�Ǐ�U��1���zQZ��|�^ob0�L�X�8�x_L�*	$k�K�Z5��G$�fY��W�xl�Ǐ�pV~^0_!\q��E�9v�)
3�� �
	��"|�ez���������U� /PtX�8
94O�s�`�@�X��6��0S��X��+P�#�Wu��L��"�.�,����u�PC�2�acc�|T�/��m �Qr��&�L�Ua��Rd\��J�*��?dMOH�����
����3�\SW5m�?�N#%�mw�7�ъTM��,'U�`A�-8�&S)"��\Z_w���­�����ٔ�L~�&��އ}��HH\� �z�}k.��]�j�vjޥ0 Ԇ�ʼ)NoП��x��YS0n�m���-V*�Z�`غo���/�K�}���G}k:Ҭѩ-��ݕ���źf�g���C�j�t8��[��e4uԮ� �V��q�Syrz��;�|����?��?�qު�#�c*���ި�jr��TK3@zN��%]�Y�J���[����g?��O�5�/-��o�J��ϐ��tk?`�|m�R��I�����j�	��N�D37�N��I�¥Ņu��Y�>n6�2o��o��H���W���馕%6������	)�䰮�"8�FI��ظ��2T4I$��3z�2s�Y�����ǻ�g�]#q4��0u�`qqA48r�à9`�� ��zY��p0 ���αn/�B«W�%\����	�^\A	;<Q�̱�<���B�'�����x"�>ʼ>ε��%񭐘��L6/��P��9�Ztn�,y�����c�<UH���T�e�b���0�\�L��1�B)���Y>8,�Q�)T��Nz#��pPU��k��j�Y�~��L�O��q�^���L�$�aNp�''�X�+�?'�R�nL&B��U" ���w<6�-��R3*�4�$ȫ"�@0t2�|eC81\���7���`~�fR�EC�f��3���)���A��s�@%���h<-W��$ �/�p�X���3x}(3�4x. ,1~�â��L*��/��p��d���VV�b�L�S�p�t{=�j̮g�uV2`M���`�^A+�L�6�u13�o��,1��8H&�=B�1��/�#<�y����{O�=�{�����5H�BQ�&��HbƖ�Vq��f���v�_'6�Cų�j�`�J�rr��w���fS����<� �[�����tV�W�)]c>%n@py"��=1*�o��pK�$��>��vv_\��w�ν����2�P�MB!0[(�#3�R��Ru�����X�q��\<#�s��S�f{{{���o�=o���_����0`������!��V����c��\n#��c�T&�����pyu���%�J�	-U3�0��O��~�X�Tdq���u��w��8��XB��lCbK5V2�]��j�,��Ј����ҡ�R��d�5�R����\�$�	%!Ut��◐S��"�w��""#S:)�>ɋ���o�� ��P�z"���G�jD��s��Q����!^YEfc2������?���_~�e!���˼��:��`h	LZ�tv^R�	s�V��z6�����Vt�y��ia6p��T0���jY�13��fP�k�D�\J%ܸ��v!��ǟ0�8��_��{����}�#4ϟ�
�ؠ����0�(��ZdY]�t��I�D���T���1���e�߿/)�~��"�3܊��iҸB4���V}�̺%���#~��mH����^Ro�y�D;H��v��O���I���ro�jQ�[��j����T��'��Eu�s\�rZ�=�قA���xMHy��lI�A�h9�/4�Y?B�"�(�D�7���V�Uq�!�;^K,wǼ��<c�.�8����&��^�#j2��?��][����8��R>�f��=�$��/��B1.�mu���r�O)�c3��&f �%Ԁ,H�R'�cq�BY{C�����������n_�l������˿����G?���E+��B�j����NΪ�����J�ل�i|o&\��I��_�W�����o
:�F�o�?���3�s8�p�3��������٦{�}���Ӧ
�a>�b�rq��(�Q�pyyswzR�U�`��S�P��2��{��r1�;�Q<í���q�n�$�L���?0��nf�N&�t�W�:��,�j���Mz��Rw�nw�أ��_�1����r���F��a��%Ɣz}"Sq��؁]�%�N_)ܜo�B=3Q�~2W..��N�L�A�Cټ�+0�����!���E�������XY�ڇDF�fӒO��6��K���B�L��uH,�����?:���A�����I���Ck>����a&�B6������D����o��Oq�a"f�4�X"8�ǽ݄��&á���#}E*����!"r]X޶��f��D*����i�!�m��q��^�KM\.�W�O�����c�/=�*K
���wa�?b�{�+{#���N4�j��:�����>���2~"m��3q��>02(�cr_[!7���i��Ѵ5��C1��q�3�l�T��*ck�؝�\�ڭ��U��z�e^ƻv�2+3�l��I�pv����^ ��ͧ�~�N-�n/�L��_;�� E����v(�=�Ǫe¬�e��Xm���d*��µ��e��^�O��Gd���;���6�'qeqi���E��f�D�r��H���a���"��+a�aw��0�n�����O���I����*X�V��������={����͛7�޼��/�B��EG�V�}��w[����69��\<�ߖ�s�z��#S�z�~j�#AJ���� #�N�^2e>��FH���F>[x���N^o=�V���DF\^_��z���=�v�Ep&{e�����B�P̕�B�=~����������d�S�l3_5��`x$����5�dcs �;�g�",'`�AX�`7��?���;WK9X�������2abg���H	$�ر<��ܪ���[�WBp�4a�4�z.!�*� ��<>m�>�N����VE+�S�&�����8Ὄ�����v���ƍ��
S��8��<��RU&)��0$�ޱ۲�n��Ħ?���jb�]�M�&$Ys�ϒ����ƙM-GGJ�(v�(TH���E:�D��8ml\�����˄:���
.9��٢�d;;;W.�Dv2X�����C���Ɍ�9���k*bC����}��H���@�ԫuÀ)/�b�J^EK����|Q�ڳ�ԓ�h�����o�o%ҡHJd�'�#�c2]x-�=�[aj Д����U�Y"�ݒ�lF���em��X*�$jV+Q=��u^�t�j�FތH���ъC���h�塚\,Rrsq�D|�/
���fi^�L�UK�̔cWm<��񈸣d������+2�V"���SX�$�=�Q���h���fx�����k`d<�N�ժ����Q��`��sB�:MQ3�8���� ͦ��P�5����5e�&ӱe���9b�.��V�j��\(%0HNcd��JU��m=}�s��ʅ�>�]���D�V�.S�O�\v^��j��xT����O�j�V'�Q#��n���(�Ng�!x:��*���[���<��ZS��jT���_-oʔ�Є�ƀcѥ9�����p��;�0�0,�(��ge��2l�M���H��?��3S��
U����	�l`�1�0���m�j0��F����秠3��<���p����R�Lg0�ԫd��I{J�PAڪ���؎��l�JoZ%��7\I ��s�I�9��,��� �
��
�:=� bT�F���N�<<��o��U���ٜ��b�pL�򯽮�5����<{���?���^Z�6���4�VY`<v���m�q�u��:J
�.6������BϭU�B����=SN�\{���B�>�:�w�^�����NjB
X�1��T�OF�qF���+�����"��ϒ�եe��u�]�}�&�����7ް�!��f�kB0qM�I��б*��?xe���Z��	Y�������� ��-�E�#M��&�
�G�b�|ÛE�x4Gc��sB<ך�M�X*BT� D��-���a�S�Ky�@ZE�9W�"$_�tɱND�x���B�O�������-��\d�cܘ��Њ�{*�Y����R1ۢ�����c9�R��B���e߃Z��s���ES��WD6cz��f�]%�܁ąc��ml��y0:x���~5A��n<��O��.I�Ix�L_OF�l��cl����~�����bz�>�'˫W��4��RA�`B���}�k�1���~��e��~����#��P!<1J, d��׃�Qټ���������GS��Y�.È��u�Ʉ��u���ԙY_H���2��"L���XqőQ~QI�����d4H&���
�����
?ꈩ\ѪP�v�^����n����3��L�勽x欮��p�ʳ�p��?R��ZO�)䭑R�ӟ�l��r���.\,����֕L$y�wH�Y��r�Qcl��0������A��>?�0-����=~ �s)/d7�u;گ�C�l��";1>"����}�a_7̔$��6���G}���4��7���f��o���~���R8�8W��Lm\'c$�O㻱I~��bx[[[A2T�2EuT�b8+J����r��%H��DU�v�#�_�w�S]�~&�U��-VW�1�gO��iHg��>�e
e�+-�V۪���K("��t,]aD���_�Ǣ2=����V��34�\�D@bm!�S���D"[GW�l�P*�G�$��*�\%ŋ;��X,R*ᗒ�� X]^Z�i�c\�Z��߿�rQL�X	�HL��ʪ�i������Z__Og3r�YK�'����m��}&8���WOK��ޔ�}%-�dv��~B4�ÐO���H�S�岵�5�b��gu/�1��À�,c�"�nzGY�B�Y�q�o���њ	��~c�h@�~�+��
p��Y{B�)�"�F{@��Ap�X��zO�;^�~h�J�w���(�4�y*���?�hS����*��/�d�zp�A��&Lw��2H"�%�G!�!�SpLy2?�8K�Q�E���<�	�ʈ{Bq6k�y"'L5�:�9��V0c�n�������\*�v����?���6��Y<;88>9�F�d��C��_~�����ݻ���y}彷��DҪZTb��2���,Y��K�����(H�^��E*L�ʅ��
��8�0�	�&0ݹl�����HOfd�a����6$�8��d��<�*�.-TX������KD�X�O�z������L�]Br�'��d<���y[S�^<�;"�ٻy��O��8V�A�	�������Mf�ʵN�U;;���gA,b���p%���W��������n:�';[���A�G����vڴm��2�ju�[c9:��ڵ� L��:�J�O)X+�-�јȖ%�L�N�tCxB����� C��o7��U+�����j�T����3Y'�a�$�
|��U��ME�b�Y���ԖB0�\�ز��yO���bJ��z�T�t�N��֥���T�@%��3;&d�u�j�L��yti�`?$\���ӑ|� #~�De����������p�;;�:�rfl�WU�&tt�i�PȄI�Ȥ,���S@��d�b�z}K�eD�ikiq8*�#��\�M�@�F�قS/��"����~�w��݁�k�j����tj<���Q�\*����Lh�����[&�a��\h�պ<%��p�V��aR,Hc8����8PPcj����L���v<?�
'���{�t;3�C��D�v�c%�;\�Q1W�t�O$'�,6o,�f<���WE�l4C=0�h�  F��b̼���y�'h�`��q.�Q�I�y���+�.ep��\8~�����gC�#}�X��"�TZ��~q�������?��7�}��[���n��b	��:���4�>%Ϡ3b��*Z��"���3y�Og��L�a3u�^�{a�_VTP:'��D�D���7��ۗT�o�ܹC�n����� {n��=�Z�iB^�Ce�a+`ukl���aV$7�3BI��N�/:�.z	�,�NO��EP�d�|�9trh
G3%�/�u����f3V���8'x4������֎g"�#�$�b`!F�PV)l��=�ˊ\�{���R�� �WIY�G$�=�¡�՚��+�"<��ɱǸ���b����zMYͷ��'�UP�����Φ���w?1��Pw� ٤�n��lc����b���v�Yj���M,Ķ��U��]aN��:�	���*-��3#uG:��1 ���_�Y�un߾��b�ia#�����+��B|<�Y���noo���6�X����p�VV@p��� �	cVov\��##�eki�ϫ�ff���^Q�Ov��L۝��-�Q�+(�E�5�P���߆w��%#�5�"ӢU�(���X�$p�]
O��"c^�p��+�1���	m���Kf�ܩ9[� �����V�1y]j/�75r_U4��������[�NW��۰.�L�6�𴍓l.� 
^��zݞɈ�K@��DJ�ᔮ���wW�X�1N�uY�2�>_��cV��t�ƍ���#Q�s:L31��?
c�\m(�v\=}u�?�p*O�3H��!�9϶w�S���;�R�LC(~��ͺ�}b��s+��hVo�A(]"6�؉ �1�Z��ሌ0�)�Je}u��X�k׮��%5i.+�=D96 L?zD&����'�%Q��m���ƙE�Ņ
�J�%����b@@�He��h�M/�$ӭF�FӯX���i�t���T5H^�j	�8�O$1����7sssa����Nvh��䤢p� ����\�ʦ�1�0�q�u0���Nf�|NIi���8<5�;�ɻ���!LX'?5�@vO�����ٔ�/S� ?�4`�*�#��-^
�@f�BZ���4))�ĸ�GPV�J��9˷��<�iF�L>B=C���o�K˫�a���°M��rE	p�_!Ey�Qa���2�v:����c��?�\�4��6�OE���BH&*�5s��8W.�������q��8�t߃��0��<aN3*^B4�'p鹢����q$f��-B����1���S�A��=��/����qey7�Д���P\��lK��$L�R��ͤ���$�%{�7��鄾v,|��C.)F=��b7� 6�"�'�
�O�5�xQ9~��R�,��lΈ*�Xf�<�ﺷn߆����վ���@\^Y�i���'�Re�$�D2y�!?��wb��]?��ƳH
9��`7;���=,($�`kH�n�9ߊ9����W�
0Ro���
��te�U��Z�TAol6q�j�e@p`�ߨ�F
7�䷟������Be���Q2�Y�,�V�n�~v�?�R}�Y�?��p���Z�L����}6�lu�q���P��ܣY��_�x
�ߙ}T���|�*&�2��b��+:	�����\b}nר�Z��lb|�9������L��oJ~O��ό�(��de|����p���LC�b��+��v��OY���Pi���U�� �s.O�A�mB������+��h@n�^��/���H����==3�즉�*�
�������� ���#c>7����U�[�͊	$g�mWx������>p�@��^K�x��7F���I
�S�z/�D��W����O���� ,��� 3Y�;��^�N�D�2dB`� �w�'Yܮ���3�p<sv�.�����[~�蠫�1������=��=��X��b1��jq6b��aV��%��۪ě ��VU9�	��p�P�G� ��	���S��*�!U�/�����RP'Nqvq��f�'���j�DN�$��ԣ^d�FR�*���]�r��˘���6��Ҕ�¨���'�?�D[�zB�̾�_a�l���J,j 55�������l��mL����g�M�e/0��chEA�h$��(��=�o�J����P,˔'ñ�z���Ap�C�N.�ȼ wAu`�g"�`�pK��9�S�d3;xeʬN�\&����ccC�9�d� ;�����?��kV:o�W ��R�6� d�%"7�F�ǧ�����<H�d�J���V%y�J���/�Y��HlG�7a3�q'�a���ۍ�6��۷��앱�j)*J7�[������@�BD8q\07�l6o�1^�;�v9��!�f�'��,f�9N��qA4�����#U��bfxW�^V�6N�Й��{ҜZ<���ȱ��D4MF��+�S	C�К���z�]�ݽ��7���ފ�xM�؊J��]��r���,z/�NLa�n6��ˋEȎ��5U��/�XY`[�Y&S��u,3,�	/��y�!u��C�OODc\�M�[��ds��y߂��X�s��I�I���'	�Kl�+x�,bE	0o�H�����!H��ibںhՅ;�1/��2����A�c6�M:�/�âluXؼZ.�����Y<�S� ��$���Lr�䗥���z�ؠ5��K�b�3��+���'͝T�M�1�ƭ��#����������(F� ��:�Ѭl(��i�
3�aH�'F��1`{а�KO�.����	Ox����Wخ"N�>��^���)�=+k<L�w���9�-,M�MHy�p���v����!_`�us����>����J�ӌ]����������w;woߪ�����_��&~�6�2']40z4&�ɓ'*ȗ�{l��bq�*�d�v�(!6D����bR[U2�l�-I_F�L������l+`4��Ё�cZ��~#�;��Z5�Kx�G^����jl�ÓcIy�k�0�6�󶵊y*�j1�4d�O���#������������F������deqIk���/�&���N����:Ն��cί~3�`�W����SP�� ��#�\ vbix9��Y?�F�T3�`��ܰ�x@�� 'Zz8Le.�GίBϢ��(��7v��}��Q�:����+����8i�Gl��h��c�;=�nd�>�}��l%�V�M}C�k!�}�-�튐��.����v�3|V���F_`��s"�����q��2�/�Ҫh��������ˆi���0e�*���q�ܼu.���Z� $m��Y{��2�:$2Ĕ��1�W|��N��Hrɮ׶V%�x[�XzdZ��?<oI��འ�TE�,H
-�h�(�P�R1��(�$��ȉEՅ���$|�y�T,���|M�sR���0X5T�Y$��l����B�"�=�a�#��>�&3�13To%.�=pv����`�O�^�G��)XA+-�`���C�KF1v2)�c�ǆm�V
��E��BF�Oױ���;:����
������b/�_bZ���PhfC���(,�Q�U֡Z�a�J�~Jd����%|5Ǣ^��W�Sh���h0ZLV����i�	��\� Zr@Ś.���i
J#^�c\�hE!%h�W���7�BC2�ڭs�q#2C�(q�𣲌�Vë�!����F2�Ӳ��4��ٖ-�BW���]���d�=0�RZ�#!,I����(�6�_���?L�BMI�O�3`��Nw$ҩ4�ʴ������U�d��ȁ�d6Tn:�v_�TrR�9c�'��x��գV��R^��JQ�6<�ke�t��m&r�5He�]*��N&���jd~���A6f����o��y����a���;6V����߄Y:�]��;�?ĮbNĲ�ӓ��KJ)c�66��ZY������癕�
;eQ!)m���E�s;�.vl�z�*d"N�)��������Փ^o`x�<$/�n80{V�ىf��5�g���#B�2g��bg""q��k۟N��E�:��Uk2����笾1��J�L������\>�u�O����a&�J�&�@���y�����O���L`CxA���@D�w�W`Dbo��y$t���{P�0/�v��k�f����,��+ˋ�'�!r���{E�pC��g�Ň\�j�g���A'�E1�OA)D'���Q�F�	�ukԄs��1ec��cHjx�G�'����y���@u&����ʠ|��7kGr\�����t�}���|��n2B9aVAAu��N0+W��qguM�3��U�Pᗃ~��V�M���`V��G�8��z�2Dۨ�?=:9=�ZJ���C��l����8P��*�a�1�;$Z�±j�^�7�ן>}*�4�hkN��מԋ+&��OeaѮL+��[aW�Z@�6��V̺��09gu<CZ��cė�|��h��A�=ǖw2Nf2�CՋs��K�aᰬ�^�7�5 ��>c�;Rb0	J;#�H1��q��t�*�g�|���q�凿�;{�ڍN�K&j}FD�9�#;�c͝���ͣ����.;�`�����itD(�o��0v��%\3�'��L
C<bB���(�,g�C7o �D�ޜ��!�%T6��Pjs-��ŷ�� U¢8f����Z�׮+f�1�����,�\�rC:2��i�.Za<�o��6`9�f�h�cX���9�a�[���Z5�*��%��Ӆo)��q2�y�O�+���V�sC]�����b&C۲0kXW��"�=���# �1���W�	2�a�3��%���'��'�g�"�3A>�p@�{�L���L�@C�.]�<
�#�a7I�*@���DI���)�7��3e58��X��ÖŊ�2g6Ժ'B+fdm���<�e5���á��<Hqd�+2b�Y\�f�K�ic0a|MxM�����z�7���i&��U���*տ���l��1E����V����]YY�p���ۆ�LrՅM��X��3kI�rD�4H1|]�P�ɴ|*L	Z�:���Xߝ��sIQ�K�k
��)O�J]4���7O�H���Xrd�^�R�8P�n|���Œ9�r_��s<�f �
�Ƕ�˩���0l�sղEE��Y��?Xk�u�x��J�ZY��,{OZ����J�S�_ŀ)٪�I�:����\e���4߷n�����K���d�/���B��Җ�^��R;�-_���.�U�,���D3��Z�~�4��!S>[[[��[7��j����9�w�!��/�k�|ͷӒÎM�}����S*�T�5(�0�/Č�_���pA.o�өUzGW7.���������!��߿���\��@�ﺱ�	Ӆ<������Z�v��p�,Mj��_=��WW�K:�ƙ��b`�~|`���GS
�����/Ȑǻ`�냸YXZ�L�F����&��)m:gF]����!��_&�[f�v�W��j���j$�Ux��l������B���n�����|>�R��i���$lC�G��豣Y��Î1�ę$���p���5��ku[r��6$��ccTݙ0�=�i�h �-�����xNk��l��Ėvճ:��Uxi�$���%�U>eG���T"	c�)��x�|
��L%��
�(�M����o���)�A�-��<ϵ�;s$76��m=��٬lf�媦�'��p�ͣÆ9N�Z=��dg&�׎c��hr�0H�=Q�|/��db`�Nk|2.�Ԇ��"H��c"jp���q��a�z$AZY4y��"�MD�A<H��	wR�*��p��.~���^���	��[Ce<�e����4P�K� �����������~�j����w���p���.�Zu��û���Hl�XK��K�AO��,h;�~�� ��M+�3�GHJ��9���bs!+b:����n5�+�\F	'o8��vs:at4.����pi}5_Y<��(�2�_���g�,��*W�EΪ�H�������,/��]��NFc����*��`8��RQ��l��rS���d���ߨ�g�J��S��I�:Xw�"����;D�.Å0q ,-��V����Lne�rxp��O��O�ŭ��o��n ����$���u�N�!T��b�T�/�������wɐT-�BY�*a*�G�ԙY`����	jihx���@Bbc	T�ǭp�p�����O�ӛ�6Uu��,��[w�<"A/C[�,"1�c���_U����L ������1NU�]�Ư�F~`�##E�A��%g�IƎ�H�5��gg55GcB�vj�W����p��@�T�~x/�(��N2ͮ\���g<�d�S.��ф3&X�y0��B/�R�_�2�[�`�ܔ*g���	�+熕�݁	��(.����x��,�`�Z|f6�+��G"^�֮p�xA5(��~ a�jo_�2~Y[�D
:e����$��,�Q:]�X��r�޺����+����`�߼q]_��={&�b!h�h�𷲠����0��K+x�2A�d���+T��+�
�'��D�$� X
��q��lh-����,A��I�*�IKu|�,]&���4�h��Ba����%����=�1 !	Un-� M��)��C�;Zyc�HϦ�l�V '��f��إ���<��}V��6��5~�h2U�
�g��t/o2���U��(s���N��V`Pf��6��/�Q�z���Fik��v>��������_��ݱ��Ң�1Ϛ�S�P_���R�ƪ!c�&j���L2Z�Cew���.HR!P	���P�S6��T��8n�|� `���8�I�b���W1l�ս{��� p���_o����m8
�Mz�5��r�u�l%�^@�i��y��`8b��T*ؙ陱���#X���C���͛�AdC��6lI�x̜����^.��>��n�\�7��.�.�f)�k��|�}'���.c�!=>=�鍔��{Y
��E���ؼ�A�|���:\Vʱ�l���%�G� !�E*�|��F	��Z��yR��SX8�MƑ@~�` �+�Z\ �(b�g¹��z��F�qM$��5�k7�p%B+��E&��b��߃e�	S�)�h�(��%�M�)E�}Y�ԥ�m��	��	ݹ��F�;�w1�{w`�����d|��X2L��

�������XU_ҍ�0�C��#E�Ę�#7a�kǡY*���{w:=�wf�ө��ׇD�I��ɠ�L��c8Z̓�� b ���Lv���5[D�7>Ŏ�bKH��ӓF���}�_ggU"D\B�GF����l��XY�b*�5En���⮮��-�R�����t(`(��.��.*"Dj�?�)�L*��q������A��B����Wgs�F�z*B�#���~.�������V�"�D����5q�b����9��P=��6����#;rj�븡 -�VX�hʲ&�V����xJi9�	�A�ݙ����G�K�bI��̯\��E\�h,�	���B1�w�E&����,���	r��X$�:<'��t���&ˤ�"U� �ZH�V9W~�<�KJu���{[; �-O�-#���f�b6Mv��Y���ܭ��'�rc�l^��y�2�ܯ�����m�ze&��X9^���X�u��ট g�x�c�ΰ���o�Xƛ�,��>P�1,��X�E)�����䑕�]��~8?���0�4��Nǿ`Ws��[����Sň`.��>Įҕ���@��'47�!���Ȓ�)�G9	����c�K��?R+VڃX;� Q��./��H������q��ľ4uj^񅰛0�?��?��}��W$����c�5���s�e�b�Xf�8�g�!����=��0�_3L&l�Ǌ�a���A�<�m�-6���"���ҋ��u'*?�����=�\9�+�L$����^C6�f��zC!�gW;��k�����P�4;=j��&)���{�L��Ld�9����h�MM��q�B�o���9��؅Q���Z)n+�b�rww���V�+�9��"��X%����L�p�b,�¿}c}����Y_����|���
G�+P����KA��v�9֪WzH%&S�l�]�?��?���կ~յR,��/_�����b��p�~��Ĩ��D���P(bH�''�?�S�W���K���)���u�;w�\�qRS J�Z�b�lR�)�����V�\G�fL
����Y9*���׬�j9�{jM'�vv�\��=�Q��Kq�l2eq2��3�wE��c2����+�L�H�����u�����]u3���c�nlF�(�R�pe��9�<NU�xF���X&Hҏ>���^'���i�!Z��� ��aN�ŌuC,P�WD�rX�8�UT°����j����ɪ�������2�lF���������2���@�R��.��[�n�����ݬU������+B���p����s�W��˸�48��ˡ�����F��p|KUm��I��0�������|q�h���^%�I�?�@u)tvr���v��/aMn%6���9M�	��d��X�����n����߇�@�;c]��d*�r�q�C����G��b�5�ٰB��`}aY{�	��ֽQ*a@s��p<1���\�8?>�m�g�T&}���ׯ_fr��$hu8�R�/t��ݲ��޲�!��L�ϸ����;�׍�8?=�I��䳬L�}����(8x˦f�P-V�|��?WX <�����{��ā�wt��l��`��|>���H���7�M�݅1����m��gO�c�J�r��z�)L�T�?��'7�]���M��
�t��y��d�;1Z��wѡ=�˧���B�p�T#Y��qF��0�
��L'�Mb�s/n5�V����3����������!�������d�>U�HgrQ솋8�MX2�̃LW�@�{��&�P��'����k�y�GS�K���^g�8\�D�� <_�2�L���Ȱ5z��77	�8=�(W�EV���h���p���>�|���sL2ưQ-Gq�ek��s2Ʉ� I�s��W_�ٽ{���ݬmΧ�#v�"M���\�z��{�b7,f��}pJ�}�&G���{O�����]�S):PS���\4�>;��q��q���8WpG�q<����T�+O��V�����(I�&��4x��U�T��d;x�L�w1x�x�J�(Y�d/��<N���i�O$S,Ԙ��7�J�����L̼M)l����g�Ά��E2�.�T�q�܋#��T�uOԘ��� ����Dr�'�B[�J��4p�'����>Z̃a�$и5\a<���| -��K;^j�����>�}�Bvé]�;��`���=i7�	���9����_��񤌳���3�X��%H�T������t�Ѿ��Og���s�0/s{%&\�֗v�(�2G?ӻ�'�O�Å�%L��Q�Ƣ�-N�I�}%p�'�_\tXH;Qlo�������J*�j���c�I�k`�e�ܡ��y��R�F~��6���sWwf>�萵����3�޻3����É���U$:���m�"ڭNK�H< ��}2��Ϻ�u'cX"pioʹ���Uw��xzz�'i�
�ݞ����ao�d��<�4��և��<�=���������*��2"����.�,������w��>� �a{
��f��qq&b�1��B�4�pg�����PQo���*���Q,[X0Y9=x����*I�R��7>|����T=+��`��zbEpqe�w�lY<`B�W��Ch�	��w�����
_��R����cQ�<;�a�,��:-BP�F=����<y�B�nTJ�pe*������x���SA��>�πg;���#��?�q0`f ߿���>}�T�Y�P玹�*ݷ4u�(E�4X��/�+O=���D��Qy��*�ؚ؏*�7�+^o��%�3ˮ+�#��c��^��|2�W-��B`���r��:V��]*�d`��6��nc��V�,���s0�J��xXuIe:d���
'�`�Ʋ���R)#+y�f�;��W�g���G�)Y������B�V\S�A����K-�{\^��c<���T��s=W���5���s��!�Mz��?e%�SI���T�Op���8n�d�SP=|3���:kVb�.fn��70�m�D�q(Z����WG����ȕq���51�.ǘ2?��������7?��Op;1lǧ�vI���fsb���uu���Xr,�ޥ���Z~1�gN�g�PO�����v$c2Q4��%�u��(�o�����==k�Q���9u�4�&���82֗����E���[M��^�צ���g��l6Ǫ��a�TI���V�P�=���)�~�-	���޸q�^<}�T1'P|OE�A*|�*��m;~7�_-���y�=X�C6�h�riE��������Yd�@�0pr�,�>��T!��e�������e�1H�B��s2"\�|-����;/��xXv��%�uHJy���C��m]�Ǝfif�a�)�)N$���ZP�&ZapPJ����>>�L�`�e��d�e�}����㜩7Ś&�M��B�����eӿ��oO�糺�Q�r�+}������Ӆ������B.���u���9Hz����4`P�X�7$5�Ӊ*]�|�X(��A8\"�U1���	�ܘ�͂x\��<�4�L���)��B�ug��1b�d�CRV���=ƈ`		r�����w�#�� �C(�t�6x�w�-��0q�S�@u����J�67�<;;�o�xIl3o�lX֓�C�r�]D�L�74J\�Si�x��Q1,T�!��W�^qokv�L�!�I�BNkOv���5�pՍ����Uv'�;�ǣu.�����������g���Z��#��q����5�]c��'Q��G�@��tnMp����P��,��^��v�V��owr&����0ux]qܘLŅS��O���歉ńT!�D��������u����#���r���р�Ӂ��R���T%ƚ�+Ƚ]�V��Pk�Q��b�$�T��_q�'�y2�QZ��}���}��%���Y[�����~��T4��Q����$��n=[�M,+$a5�\荰���'�':*�fT�� ��]�6�����-�Lf��eD5�T��>5:�z�>,:�ъC��8˪�#T�p�Z҂k	ϑ���hO#U��~�J�2���1��٭2��1�+�mL��JN�Vӏ��_�2?���k786�g�t�~� "���v�ַT*߱�\U��qVz�.I0�Bc�U).�[��_� �Kf�<+��W�W�@8'��5�g�*X� oZƠ�i��Q���,5qR�>�bT�=)Ձ����.(-���z�!*4���`9�Psi|N}�:*=�q���_��P3J�7̯^���z�U"4mQ8y9�9�?��S)<9ΪՇ��!���t�'��e��f��AV-��u1�5l#�F��66*�E��i�a�פ��VL���C��f�6�TA)ԩ��LؖXQ����p%�;��恰[���i�� �V!8T��o�H��Pk�,U�c ��aA���`���d"��.��[ki��U,Ս���P/4ε�!5�6|�"�>��sL(�J�W["Ĝ|2�*��rym����P�R貓��[��T3�DYe5�����;��k0�r�cͲ��D�bkJ[JU(u/�!,�L�KUݻ��Q�T�fU�����b*���s([P#�\hiZ	����Vc�#;��� æQ�̴�c	ѭ�;?��������oAW����}gջ�R��J�Ǯ��6��q$�R����%�S����^�ф�����y�c��j��@����^�X(�ҍT��
��
6���Zʚy���l�p�UI�x�`Ίc*غ�������T��e>|�����-÷l���@N����q��vn�y���������]��/{;;�{��r�#h/�~� �d�MEK�lGݶ9��DW+|.<�-�ܹ#/;aM�4`�,�.�O�R5UD���p9{��M�^��9�;���g;�_=\�X�g`-����	Y�'��U�Dڒ1��b沰k"Nc�4A�X��5�q0�E+c�����^�#�����D�F�.p�<$#�B���1#	ɪ���:G�����x��8;ð�b{t,[wy���V��ޭ�р�].��,��Қ�m�6���&5�Pg�y�3ΤӘ���SxJҠ~2�	ġ{�b���%-�0��m�ı*w������?Qp�b��.��Z�z�j���NY�4����"��시CR���������M�R�Zn�EҺp������������n�$U��^���[���䊆�fn�P*�n�{�V��j�/.Z8��aH׮\����х�rw��e")�+Wr����J���G@��%�����w{}?Ɉ\�P�U�Jg�[����XbXR9�
��LI�|9�Ck�Ĕx>/ ���@&���?�ܫ�l����)��c�^�`�r�W%�B��`���;"�!X؏�p��<�`L�D6��=��p6ݨ�	nh��>�ˢT����TO�"���U8Q��%i��(��(З2/g{��8's������y���KMjO�|33^�2	�#�@�",�:�
�PE�V�U�n�1����0�l�8�->|��ǟd��O?�����F}S��|AX;�s/!��V�n$��xl](0G'L�es��_6i"�i%�16�x�SJ�p!�i]3�[�q	2��ý�ĜW�q>��nM� ��;�𤬕Ԇ�C�Ae[��	��D�:1��gϞ9�ݛɂ,��j�(p��f���$�v/ǜ*կ�V��7����.�_��CЦd=j��/�rS��w޼~]��Is���+�y�(�DJl���@d>�Z��������w�>�%شo�2U��(��]�T^A�٪��lPuvYW��LEy�;+�,��J
��+�~pK��
��[T�N8�X������?V����v�����;0ZqA��qk�F�}and~��`<�0��4�5��5���1[*u5Q��jYF��Z�$W$@\��:�f,�Cfl� R����%d��kX^��:M�7���&<�X.�ux�_~����.�.9r�����%�X�bZ	�g������T��aK�qM�X1l�+b�޽{��C��_��r�?���5���8fnf*K_(��X�c�U��I%���c�V��eѵHr}&V0(�rb��۪W���:�ԲY'�g�ߕ���O� e�����ݖ
y9�7����ȕe�,��y����bB�<����2�x_�Y�\�Q�M��'�K	��|GQ���}�o�90�t.-?�uH�$)�3�2!��,tUn"�1��Ȝ���D�lwO�
����a�gD�����/��/�?1�w߻#�Z��� r�����h�ⰻ�R�g�w�����!x����N�����@~�d�n·#�/�v��w�K��Q�C�戮�{;�O5�X�N&8�Ys6���c�C�,\�Ӆ;)�*���������TFz��L���x�fk{'�yO�=��1Nu��}lٌ��	l�n���Z疹J7ެW�G��Y6��������(��}wpx/�?@�+⴦�H���YO�UJn������0�)��e�p��B����L��4�i5���q2�s�J��ݤW̱H����MR/��W�P�!�r�X�TJ�-��},��W��Sa(���ى}�1%gg;9{�v�$�Sؑ����ɳ�>�L14I�Q��l�P ^�����K{����/fp���2�ӟ������{hd��m�9�������6���$��3��ϭ�)�bV� 	M	7w�J=\��\!/����`W���N� !>D"l�\�+��]�d5V�U]���1VYU��QF��,�s�j,ܲ�/蹢������/�;_��n�GG,c::�
���������3i&�䄎�E5�\�:K���u��dx�e�L�u(eE�w�%e�Ǩ:/�3��7U �ʤI����h�&��sn[��ݻ�A��x���d,�k7na�\t��>s˟|�	����O0fu\��[��/m�`T�}�����&#ҴL�6 zn8s��(D�n�Eߗ!�|�VbҀV��d�Y���Xb�����he�JC�g2dmb4���c�R�X��!�8�E0ݍDmi�/9���D�"���d�l?L����U�"�zS%�
���b���޽�,�����PF���?��?��G~����oݸ�)m�[[�[Zz�(p���fZ�E�f��f;�l�l3����,t����>��2-�]jls�\^�p���O�!����H�Z'­�:���6~���t��V�8L�Az+FUB��3��m�:���|�g�?p���E[磏>z��9���%	]*��7��:F�$sX�8R<��D$��q��Tu	:{jMq��U�
��D�;N}��L�F�L?F��"��c����ɭ�6d3���wa9�A��T� N�]*���?�#H�'O��ƻ���e����v2�)�Ėj�/����}�$����ɝ�Q����%~�rbG�e,��55�L!xj�V���+�	�������|�ҥF�By�lV�z�.*QVH�-=X�.�wT�`i-Ҍ'bG�4�aDB��U�	�'SF,�G��_g�tH��YY~V�+�z�Όu54�Z#�oj�p���#��<��&�}�Z`�0��Bafd߽{wM7B)`4ˌ������y��{��ГZC����h�	�z5�<�}��-��/�"��\D��\��T��5E�=!�O�q)m'(oxQ��^���l�s
�i)5�Ut��U=�i�򖔯�㧌C^q$����h:�1�&&*,vU���<^ߺuKL
TZ�&fO:�l�Q�t����q�Skg�5�$"���/)Y2,T-e`9vm�لMB񔪦TfTy,�.����R!��;��2��r��*�M��s���O>|x������+8��*Ie0��^���I���?���6~')E��V���NΚ��ݭ}�H�l�H��v�;�-,�Ru�(�ɪ9�G� D�9�����uR� ��Ų�T���3eM�\q����D��t�&��a�O�Q�4$#rP�hA�R68y�6WWiC��&}6��"��.�,��f�E�5��֔�!g';�lY��E��>�>S��K�Uɱ�w����M���s�*i�����ފ{(�+K�/ݾ}���E�2:�xF�G�ƥK{�HXϬ������;k�̏r���/�q����?��^�?�t�L�z"0�u/D2f�ys�k�9㊀�(D �T&�S�G���?����;?�я>���s�.����h>��1;�KE
�;c{��3���_cY��t�DL�&�+v���2p9Ĥ��1�Lu�$��o�;�c`I:I�Z�V��[�6=#Ǽ�����Qْp�w�Y,�Oxp2������Z)���l������x���&"g�n�t��;;BQ_��,��B�g�[����������؇�Ǧ���3&�`��aySQ�Z�<.��sy:	.|w| ���Mn����#Jzq2�Q}%	��8o],gf_�S�"�<��<��S,܄ca@��T��/���$�2��X��3�!��D�-�l�"\��*�e@Xig̮U%��uǎ����4�o6>�7�v���	��͝�(���ϦsZ6p�qxfU#ʺ�s��)oC��b�T���E$����&����T��a`ET�{�;I�N��/&S�2I���K�ʿ�Y���������o D�k��wL`��|����g�l����+��޽{a�sq��5�.�M��}�G˿o�6֩�&>��\������͟��g�/_��!F�UYS����s�ΒΕ�r>ieD�������M�S�d 1"m���2�jn��]lXE��"�������F�$<NDY�5�9��=T�!����i�k�$DĽ��Y^R�i��DU�Ɗ�P�t�jl��(܅��A-���D�a��!�	�]��V��>Xy�5B0R�(�ET�h(e)�,N8��5%�����΋U��T*� ;�L���"jo@��ι�:pwT���v��<���ZU� gy]�+H�Do��M�_����,�L�é��p<Qd��;;s�܎��k/�T�"e�x �om��.�J]EHTE��*X�J���S./�'�a�ˤh���F�S��o�uހ���l�^�ӶѤA)���ʕ�����`50�E%��z2��F��]���fa6��3�B-N:˖ƻ�Fx���R`Q��}(f���&.J��\gi��2��p����������P��hZZ:�x!��n��|����{*<^=�c���t��rS��*���0����
�p�*d*á�z�U����z牓²/%s�B���K�����[�Ô���ΐC���1x�@�Y�<V}5�ǣ |9�g�8��7�Ų��0����(ؤ�lk�hsn1.�����*���r�TD�V���9V�?����
��P-����u��?��X�`%pD�����|u8�̢n�uo0t��驔/·ĐN��×gm��l��6��$�����,Vס�vm�;}���bac�Ď�i)\3�9Hib�Z(�Y��Q� ��`8���4�D�̵����>� 0e���8��װ�������X��f,�5?����AD���R��Qq�P�	�k�W�3ܽױZ��� F�S����������M�*a/�7�i���&�[���<"y�ZU��ͫ�p��߹�AZ�J��ըRV[�ĭ��֪���&#FcU/�yP����R�J�[�M�F�(��[��3ʽ���#������=�VQ�A���ٸ?��K��5�w8�'�!L�i0�d3J�f3y|,��$����
!�P6|
�)mCU�ωjE K���R��$�U�]�Sb�%m�	��&�LTl�SU)�gҥ��E�� 5%`D(Q�@匲�Q������d�p����<��C�h�a��Axt|�Dk6U۬�g��vk=��XA�=��Ն=T��p��eL9�aw�2v�%c�
����`������҄<��Jw��u�/��3M%1�<�[�:f��|g��ު���b�,̽��ª�b
A�Z�s�ݩCx��8��й��
ޚI9��T)��,�.� ���l��v<׉��n8'W��V}Q���F��]H�ޠ_�؀�Gʨw����g�1�* .GS*!X�9�%*H�c1^�1��$t^���q�
�Ρ�D�ݕBH�E�2e���$0��|tS���2�(���_�����!ֈ�u�	v/&��c�Q��8�|�e� 
��� \bg}����==|�O>fao����K�o�68V*;���_��W����!�DI���ԈIs�R(\GEƾ���&k�%�8f�0]��k����y� 4,5X1x�Wae�Jhw�9� �����;w��L�F�%b��7��0h��[����a0w��z�0���b��T�����.8C�f#.^��K�*���	����,z�d[;���-+�@`a������۷x�Z�Q���x_�3e�)���(�Z��7+�ڵ�"}�5	fs�q�d��Ue�&��-\K�ƩH�,e����Icy�x+�rawQO���ۿe�a���i�\\�
�:*AW��5�vH:L�� �A�� ��F�v�hw����RpI�h��Q�T�ױ��(\:Rx(��)��eÙ�O��I�aE�B
�eC�Ԫ/LƗ�u"Y�#�Y�Æ?+>W�Q=���Ey9�p�j�$�8��Ch�P�4�t;�x�����H��0�z=�Ή*���8�D�NlK�� T�g}nhL�R�9눮�|��T��;,��  k���^������ˏ�����	O��Ŝ�v�~U`�@��2�,��h�Eƕ�+d��'��sϥ{ں 5K�T��Tc;�ɣ����SO6�6b0�զ+�F��u�dm�\�?ʪ8Y�͙�%�4Px�8��Ċ9�����S˄��Qm:���r!��W������6�����l��g�#ʖ/����"$}>[PUf�����T+M��||z��Z������È_���i<�6��s`ఢ=!A�D{�:�1X�$[��F'g�EåXw9���t���g�I��c:^�?�;���K�lF��8cv��x��S�y�"��8�'J�B�T�~��,4,��E�ޟ}�Y0a�� �^;�U��y����Yި�����'/��T�cm������:�e��i�����\�|Y���h�1�((�*���Â���~����駿���<H����ط��b���А�ЉR.��~��J>�۪o⑷ju<��]=��������xa0��Z5��:�5����C�\�p:c<Q	�i�X������Ȼg0s%T��,ץ���bI=ib	GΧ�;��Q�T�j2�d�)%i]�Y���� Ĭ�
7�;aߍGSQ��� �Ǘ{)�DHǰ435�1g���c�iùyґѪ��i��߆��#X[-ҳ�ˉn�ҹ��x	�9�F���}��d9��d���&S� ��I�a-��r���Luح0K�ӄ}x��]�K:���m�݀�N��1�O��Perʘ�K���?���%(�E�e9��:�}�}�D-�T+l��'3��"N'p�FCX\�yuw��n��ugf{{kǔ�+a������ǌ�ڤ#y��mA�g6�9��d8Q(x���F�zqњN�jЄ*��&+G���8�Y*;g����`�R�'�Gc�>�<c`)O�����e�&g�d|�Q�k��ث�[�E�T�gx:�ٜ�_�	�X�`R�$��-|?��ǐ��%�7�\"��X����WA`�x{�+m�"�/T7���۵�Ӿ
H��Պ�k��Ȋ�����ͭZ��Ɗ�Ճ��-���O�yƩ�q�N���zrm�L��G#�������/_����h.٢r���n�*v�ڔUrIn�lj�H��_ʜGhe�fӥK��r��&d+\E|g	6���׹<�zqz|h�&vԂ��t2��*��h��8t��:�]�ۇ :9x'�KϬo��ꤍS'~�"���%����.Tn@���ȞJXKsen�Ϙ�4�T`J9eL |���~�#�Zd��e��?�b��s2$�I����!V6��C	��Z]�cd>y+�q���e�I^� �2����"zg�{�lr�U݀��ٛ~t��>��L)�C�֬YJu(C�[�fl ���֒U����D�֪,�n�� PG��H�޼��7JJ�
I��X Y\�B'��zkc��pB�'��ۜ$Qoi�9ƻ���mԚ�*��Zn:Q�Y2E��_�ߔ|Z�K�)����;���t��͛�L�ɓ'�9�M���)����B��B b�JT� ���U?MLT�`�;��LꩈAh߈u1���Z��������gح�"iF��DǪ��F�Y�+Nfq*Œ�;�7��xb��1�x�G�ȺI��A��)n߾�L0��ml��*E$����W�Le@U+.�K�Hŷ�Lr;��Q��nJ��1]�	Y#&��.;���"iJ�.V�3�ϥj��FS�{�mO�ǒa�0��f�,���ɭɜ�hA�s���@��9����h����B�>��Z�G��L�J���l^<��Z��
�E��矏Ƿ��]�6��U.�]�s�|� �8�8:�ΰp-�v�'$�cӈ�
�,D�B�������,b��v/` d�0�r�/Ch���f�U�נ�C'a#$�|.�2�0����G�u@�)^˓�x�۹h�`��޽u�t�b2�$ ��
�L�ө�k���b&����8a��L��J���P	�����kל���\�Z�]>g�>��r���2�H��iz(/�}h[M��������� /��'a5�h"�Pn㔍�´�,���a��V�{��ɶ޿��s�!�^�"Y"޼~��0n�piw�j�������� �Jy�d��ʒ�:-y�f#�����?	�6��I����AY?o)G�S���J]t;�vK��[�j�Ϛ���b�`��q_�Vs�)�L� �3�dP�=Z�3���ىI҅��RBhE��b�U�oJ��X�8Y����z�G~2-�Rj@W�mm:�5�fYy�q�Ȗ��[��\.U���/����/��c�/�F��`0n���z��GF 5�l.�����͇��z}�62��K��6���'��x*�8��lZx!S��l�eC��������x��	GO�+{���jZ23%���i�߃y�	�	��������Q����Č�%��Y��S_��p� v�3�a����Z�{SF�[r�����h�גl"2�r�t�n�� �/��t��Ier���Q�Qj���X׎�CU�hN�
�DV�^v��8��QX{lK��ɚs���β����,�ܣ�7��JóB��B�e�	je��� �8O�ó3����.��y����|���	t������y��,�����g>�`�!�}��e����� Hg@�b�RY���6	:)�]��6�_�ثc~F���7�'�ffU�R	ͯ�&�,��NKNn#����Y۰��L0.+&}4`��Ɲ�XAJB���y�����d͜��/�f�J�x||�1߽{�r�n��D�5\�}�펄��9���u֕
o_���0\Y���A80!8��bި�|��)����_��\̬�Z�W,e���D���x����`�ɛ7�on��'?y��q��C%���H06�S�	�s-��bםB3I�qq�|T�A���Z��{�����Oz�^�d�\��L:�NQ����z��-iN�B..�a ˨�UT.�p���+�æ,���
�&k^�9S��rI��4T?�!�ްd"���2d��Ux/B!&�{�J)��X2/�r<=O���d�l��E���X䏿�ĵBb|U�า��Ζ��9�Pr� �U��@ĥ}�e(�y�@�L�x[�Tu��3,NT1����Ⱥy����tX�E������eZT�Fwg;�
��fT���L~ ��JA�K<����H��F9�;`6�e�+��$��22��2GaL����˙��엜	O�ތO�YY]I<�-���|��,~�KB���p2��qT>b7]{b(аuX�؁-����V��yE񱪕�@�JJ�8�$3�[�D��۔�(��?<c�}$_��	�LS#����{���E%�Î�Q�*��/~�;���ǰʥK�|	��u�M�[+j��S�wZ[*ND�^��6��߼����OJ�+qz<��/���A�L�am�Y+����=��s��F���&��������:ǧ���G��� ���vJ�!�܆���?>:�آ��(�Hy~��_0Ct�&Sx0��S*Ce�[c?S-�Ǖ�
H��H�[[�f���Ҙ�7�9C�Xu`��gSօ�,(	=71�`Ѽ{ssN�6�0�d:a%����/^��p<���~"
2i�Q דR��')?S,UCK�.�s��޾w�6������9I�a.4ޕ
�L��;��+��A���ܕkW;09ˤ
�(��S�gϞ�v'�ϞF����f:�x��+(�R� %�0�F�&�M���n�>�� Ծ���B.]�Ґ�7knLo=MԐ�[�s
e�~�ryn	�M`�Tsg�y�1v|:݁c>��P��3��2�Pn(|qH��n,�ЂKqYd�*�r~�-����#9�|�(�Y=�5!r�jJ}��ԫ�6�r���s�ͧ�Ao��*䕭�6�ħbM�0(��J���Q�X�`�)q)fo�O������#��k&��"�MF��AP@�|���ytt����o����}rrzlqm���8��[������������lz[ܚ��ۏ?���{����#6{���f���K�ξx��1��q�J�A��'�E8�X���ٰEYT��q��(�'AM����d(�f��>ƃ�>�h-�R8��j.�ouب���+X�F��+bG0���W_��5����g�&�
��SX�	Kg�T"f��g.=�Y���%�d����d��ri��R�b�y8R$�����h�|uhF�rp��4S�u�JNb�z�z(����g��ͺ��G*��ȣ:�;S�e0��R�ڷX(f2)�IΛ�D3�׿��Đ5J`ܻ�>��`^���j��N$����j��F[�p�e���J�?ڟ���Irt�Z�Ѵ��ۑ�`{��ԉ���c���Ȃc4q����Z*�\le#J{o߼����U='eުO�߷w���m�`r[��B�Ck�h����/_��;[ť�f�͈y�������-�+�R��0U�J;�P�ܬ
G?����^g����A��;��Ӧr^��HR��g'ggF3�;9n��T�;��ݢ����P��w��99|)��k��'��x��'Ҙ����xC;a㲟ڜ��^)Hu`�,���M�KP���8B@��I�n�a�q�D�@�|3�V].�AH+��g�Wp��wo�D\��NK��������E$�*a��ӓC��/��/������"g�V�J�O�Vc��uQ�˱�K�j"�	�v�L.��S���	�t��}|�����@� ����}�6�$"vV�>���Ĝ����l>e���G��^(���'+#��P1P�J�bu��(���1�P �t��U6J��
�dE^�2s
�Y�e��c���E�b��6�*I;~�ₖb��
]�����A~�oMQ�cÄ�dNNp
_c�0���&qk����ڽ�\�u� �x�1	�ǟ����u�U�tHl�>(=ڪ���2|��7�Jܕ.����Q���]"zg�ʥZ�5b�����j��X�]�/�;	C��s2zHj�J�J�w�9&.[��+����G@T�aTQ����'���mJ��9�ɠ|z}��	�h����uD ����|��ɹ�{����6�q01l���!)��������B{)c���X�����w,#�P���q�P�J��
�elMh#�p���u*��n�O��,��������X��wZ#v�e
�;"�h��j6Z=��������~��o;m���`%A���~��/���x4�z�3[8h]k����"l��kc��t�2�*��c���E�M���g�}lnO��з����{gxn0 ;���b�� *Gm)�9Β��0м�[�����%���ϟ��%wt�l�DaH�� ���Υ�
�q�8�ڽd��I�����p����Ja2������r��{1l�񨷳]�V+8��Yrrt�ޝ������\Z� a���Q%S��
���t�ژхbC�Z�Z2����{Cs����_*Γ$��ǟ�����O~��4�s ,��l��TC0�v���\
���(�#F�٪I�ҧ3�P�+4���#���~dFeƸ�?��?���A;��q��;D�Ŗ	O�`�̴XV��U��yʺ(���I�D�6��`���=m`P�a��3$>4T�(|�J���T�M.�R��`��[K�i�
�7�cb��Y!�$hEu/:�o����u���mCh�g��V�����e~Rb�m�[��ܥKW0Qb6�?�:m܈���F���~��m&K �����R�I�v��y
n'M������T��o^�a�'��HP°�]ľ�{0�ő  ��IDAT��	���[��}��{�A`��7�M�+�[%ՠ�0r(�++���?�*OSl�9qׅ)���l���
�`_�'X�����6~Ca��0���ξ��r�P�DF�/몤l���I��Pi��k��L2�g´�q�4��E�=�$��%�.�F�3*���/ٯ7��]0�BV�0Pt���y a�0� �T2|�B���F�t��X��ku"5���I���|6�K��q�?,���[���j����������ϛm%`ם�S���Kd�|�Ҁ2�4Y�kOA!�lRZ��/�ßY�w�lg��|&#m|�&Z�����`sE�� �+�fI�l	!;b4�Ax,�k�eShHʄ�����I���������#��~BE[l�jm�q5F���¾T��z����>�9�,��,I���+៶F��-�wi��ha���/Z-��}��!���ׯ�ķNN�Ek#�A}��=�Y�B.�������������?��O?�T0LG-��}5�֫Q�8]�Rs�vc�Ab�E�1�$ỘNO���g>|�1o��c4�ei؅5=���t�TT�6�9�4S�~2�X�$�4�� Tѩ&Wʴ� L�K8�:�)��Ƞȭm��b r�U�M��zb
%�"�"р�9+�<a�����-i5�%�Éu�� ¨�x����Y�=|�>�x��x���LHH��q�^+ۡ����JS	{-?C�a�G���L�&rˤ�@��ΈCMz�L��9V�BV�0����i���4��մft_�T�*�8���p'X�I��m��T*�]�.Eg0�BS�Y��'��Q�
k'�R��ls_&���#+��c�z�U4���B1�2d0M��R9!�Dg�8D����5e	�&�ػw���׮]��n�g�T:i�qQ-�t�$���|Ոh���U{�^�#&�КVh�P�F�g��V^�cb0.|:����'߁�{pt��3��eY	��⛪�h]g��KO
��'��*{	�ˆ0��N��ڪW�L�!C"�*f�I'��k3A/�]:��H��j<�)���vӞ2|�rܨ��P�/_�$u��:�r�����c��
����_ݬ���#l>[�����(�L�C^O��ReA��73~ʰ$���o�z�t�L�zHSk��j^Y+��7�:9>��)���-Z:]�=&��;{�	$���ƚ�fV�GC9[�J�s/:펱5�������d�g>dKe���
n�t�o���i�j/������^ڈ H:yޤb����"�0MN�?����?�Ͽ�ַ���_�Z�h�N�+	<8����X7��Kђb+���^Z'3����$��@
X��d�2�u�)��Y8���YDI7a�����hޔ��u�\�u⸥|a4J�wz�|.�\rϘ���6�+ggs��ɛ��I���w�y��s^�"|7� �ZA��3�Qv	�Z��^6�.�E�j���o}`<|iH���$��h2Kx>�����> Ù���
���K�p�>{�i�<B�����;;�O��t�ՄO���6��wv���3hL,����ʪ[�	g�@nZ���;r&�ꦬ�R�W \>����+�v��w޻�v<�d���,�\t����3�
`���׷`"���jwZ�p��/b�Üc�`ʇOi�B�:�Y̹C�%�#j�t�����XP�=��B�9�*jO�FO�Z��������fV<��r2:�vxSI��Jf�R�uC�i�5Ղ�ab�~2�֪�AaW%�b�˹Jͫ���5��{��#�/�g�w� ��X�%%$�:�j�j.�$MM��yЙ�Ǔ�Q\(�z���#��qZ(d���V}��������m�������|�۷o/\�M=�����ȩ��]å�<��H�����Gm85�l��.i��ކ;\F���+��9(^{|����������	Q�*B�ٮA�:��`T߀1g�	�f�Pb[�nvI�,�(�=6��q-rm5EN�E�g�c ��l.��l}����p
��8��j���d|E��M8��k��1P�14*_�?�K��N�Tqe�
,U���*�6a��B��(��{�=���ϙ��|���|K����Ce��v_}��������>=Ue�F�$#�1~@�
4�������&ŨK5����H���A* 	Y�&D�: N:�-�Su�
|ͦs��Xr��K#�إ�1		kw!�_m3I����p�3�v�:�r"VV��l:��1(&�$7��\�NjY�J�ռP���G0Y�o�ޏr��o�6��j|��U��+@>��b#�^�B�)���&�ׯw�@z��Ǌ�U�
1����U4C0Y�L)lh��9*�6��)�o�"�U�-��T��3�	,o�H�!je;K׊�I5.���l��h8�:7JL)m�{h_�$���
w����Ӊl�8	���tH�
fr\�+�e��)D����QxJ�
cHm�V]��Sި)i�c��!7��@�9�!�űӤF^r"mf\�.�ּ �Ӥ��<�i��(I"�b]�"��pA���{��x��L6w�X��]{H���� ��r0nd�n\���/1���r��O�. W�¿M������.};r����Ѻ����um��<8<	g�����߇p��/�h��Q�
M��:c�2N��%��rn�Yܧ�����b�E����kb|k5F��:��~hֵ�M���\��n�XFV���,�rA�˿���}�3�4����Ȭ`��+Ͷ-Wh�b1Fo�g�%d��y�V�������R���2�Y���,bi/���ӳ3k>���͇1b*fv��K��EM'�Jy#���g/^�$F�l9���\�=�8��+�x�6�	?�V�-Ĕ�.�S�c5�8�_��1G�m�ڷo^)0�X�MBs�J0'ld4\�
����x7*�N�͍�$[*a�q�7�T2H���EI�3�$��@��u����d(��1�4�D�:'���O*da��B(O��Ƭ_�Fd�s�
�ŋ�uj���r��ݶ1��,f��f
Z�O�Ii�uA�o�e��w�0�������Z7S�N'���
W�z��i*��x��d���\.o�7D�Ŏҩ��m�[�ӦR-��a���Q.'ݬ��]�5�2�he���|p���O?�Tiv	Dͤ;ڽ:)J��h��ք��KrI=����nd�z����F��0V�(��p�ܦ�+\���,���&� �g\�`����F�\j��˝m�M�-L��;w�?9�"���zL��ߵ��"�ZwAre�*H��� �ǒ�6����|��ō/"H��٪\w<::���{7!!���20�KWMÒơ"ʙuZ^HzǪ�$%�Jxǲ}.+�_��@�!DX�:C�k��Z�Bx/��9�9m�b~i�Z	v���l��]O��B�?9(n���B��,��_�	ο����6�8R9qh��`'[�h�|5��e���'�
|�xB��|6I��g�:Q�7�U�l�8o�U����u<�={�,X�!��ǌ`B"R!G˰��� rWNZ> �j� ʯ~���ZA'���@E���f,9���uzB��"���N}�T��H��k�CJ'��K�]Qz`* �|��RA�Y%ef�ז��bX����JWk�V�٦x>�s�[@�$-�)�_��c�\WB``��j\�"׮]�`pބ\�LBI̬ �:�!ae�Af�1�ՑE�M)LD��n�K�jqEI�[`�U�f�w���Z+�.�8b*���Զ�9U�I ��T�� �J"�.�Iɏ艰�R!�je(a�H�˒��媑.'���h���y��>�~ծzf{QB)�mGt���xzz�����3�)�3>?;���^��b&Yh����a*��T��op���~��f}F�˗/�RZ��X7"�Ȃ��O�|
��MB���Vn�p\p�a��)l��gS���]'L�'�[��"���+��7��q�#�,W¼��5��n.�,�`�`2S��Z�Q�������"A�H�I)L�G6�[��	W.��X����R[o�5�KU2�p(?�d�E�
zB�J�0e�4�`����Ζ"���9Zҕr6`z�9xI�`	3=�v��aQf�Y@x�ϗ#	 +V@�-xg4*�)V.��C+ey-k�-n�������o�+�Mz"�f�5_�g��Q�����"�K�,-΋S��M�Hg��B��/'٠���#wz�d	�^�D@F�8t���xҝ�i����Od[˃O�;8���.]�l�x��v6|���XY��P)��5��ի��� �XOo8N�)�`�v���� h�mb�jX�[x/��V�R�Q�_b+���d8�q�����)\fL���^m�κ�F��E�Mg$V�99��BQ�6\�\�����\ڨU7q�OT���7Ά�N�Ero�J�`v�����R6W����0�.�����b��hL���we�(ķҾ����qw�]� GQ8'?i2r���.��"��v�}���i�3����d�9x��I�I,��h[c�-B�	ۦ�i�˅���T�F���cn�&�	V�Z;��%!I9G��A:6�>φU|Ƌ ���ƣܵ�ϖ���F�OVd��ё�K���6MШ���b��KXG�F�ec�����-fsl�t��Qּߢdx���p/�狂��/H!9&A P��~`��L��%�O���x�)D���"�e��[�,���tz?"سO�<?�+|��OA*���?�3�����%�T�Jx�UR�$�rI�Upu�(��⊫t�@���Ժ"2P���,S����&��۞T�*�W����0����̊�*8,�����3�)��VQ���w.��	���-���4c:�_�.������5�?͘[��4����ڽk���e�J��
Z��
?����⃒>��*�*$�����c�x��j%��{\�<iႾ���i&�n\����l~�=�ǰ]㣋Vd�B�06��!�_%�Y�r�2�B�3��� ɇy��A0����@+B���F��u�e �s�ܿ7e:-E 5���ٔ��P�ǧ�Y���"�b����~���!3$X�"�ݿ�z:���ͭ'O�4���9��^��$�hV����.J����2�MeUA:5\����8�BA��j6��4��Q�\ڿ�X�K�[���"*�b�Q�o��G��X�5`����Ga���L�E���䥺0�;��X���Y��!	kٽh	T��Ǒ+&WgE�8R�^�h��"�eY ƢΖؠ'4""PS��!WRm�hWƃ+�*[\9���ػz���0[V�M�[ȗ�UHut��y_$�,�Ogx
*%���3 �ƻ�UH]hA��ʆ�UV֙�}�2�S.����m�� ���2c��d�&S�\f����q�����-�c/�C���H#S�Ib'�I�(�����D|�C%�iO�V�<�1v���<=����ξ�I�R��AM� ?�jU-GJ�o�Ұ�F�������a���1���q�S��#�L藔��\�/֝�W�Wq8�F�N��xN���~�M�[t}�]e�Ź���X�(�>N���X�mR��]Y��Kg�ԃ��t�,$h��nĄ��E���`�p�zF	��/dWh�q`®$'G�����ׯ_�1�r2ɭ�f.)��|;��f����R�#��ɱ������ɱ5b[�ٰ�Ņ���0{0L��-XQ�u|���S���$��#s���S�O�+��L&�R�@q���|KV���遐�Z�n�`&�f����("�x\�F)�dg�����9������;���P!�b���y}�hvL��Y)�p&&��wr�7aC����nhl�is-r����4�<�%�f�qdt!�gb��Ŕ-��E�f�af�$.�A��V���!��xH�w��U��p���w�j5h�F�M��O�f����0�F<��U�|l���Vz�5��6���v��?(���=?oB�@��9��F��;R�&dY����7|�����ܯ�ݗ�q�ђ�aS�Tv8�.,J�Q��^�囷x.qn��B�|�\(�� �y4X=����z��\��Q���왟�1	�Ϩ��tk6�snf���H�HGݓӃ�dԳJI�J(�cؔ�C\qs����;,7�x�*ڍ��gK�'K�ዊ�ȔV(+��T[0�>���v��Q�XuwX�s3���@���୎�kiŬp����Hq&[́6��Jr��c��=�[��	� &�db�~�A�'VA�ld	��-�*A?��8'ɨQ�y�J��N\(�B������'Qn�2���j"���`��V�b^�!uo�~���%�{<�ުcH����D3;n~��� �p�Xg*�QA!��n,[����.MC9D�sUp#��3p�S�7��0r0�~��,�c�\�]�6�=#�M����C0�f�� ʕ��4Z��&9Q�]\v8�C��0�>c�}�O��ڦ�'-/��if�g�+�/�JJ?X�&��k�#뙊U^�@=z�Ą�hz5���5D�hV���1S�H3#�r*��Ek�8��F�ϵ��1�d�C�S���^����]�۽lvVC�aS�+bl��P��`m��{z�E�e�!W�4QaJ��l^Χ19��C'¥&ڟi����x2�L ˈ�ة�`x��.���E�{������6��H�%�m������/^�P������q���TC�fǜ�e�.]P&ʢ�ia���h�Ï�;>>%����V�R��U�$m��؝t����&1 ��"6�|dn7Q'/�� O���=�ߌ���LQ�n���x�B��B�!����{{���3��+�sfE�X3($(���m�9q�y%_x��ya�e�ɂ�Ť�������l>+܋�q?��O?��O?��믿�B`x$N1��gIo���k�@��#3M�1\'�bdd�|~������VYx'b�&S��Y�Z�X׬����t�y�ܠ�����]՘(�T�$���P�d92�똀��BQ�C˸�.(-/T.=��Xȼ5�Q�:c��ʩ��9���ER.<5��)B������s�u��ZR�
�IR�`̮�?��e)�%5&�8_�	"(���R	XbOm-��a� K�k뢥X����������v/��|wm?X�Jbk��.H)a��ːw�<igϗ�O[f�I��_35`℥^g��O'�@!/H0J�LZ wR7���{�n$�
�,f��g���`�}����lW\M-r߼y'l����E����n�łR*^����p|$�ּ�5����Ŭs!��h43�u��<�^��0x�ajtq)WW�"%����IuR�f��_3n�����6с͢Ƌr/fH�Y��JD3e�Z� 1�����,7���$i��eG��T{���w�U��8�+<�d��<�ں��u�)�����h�2��|�^Ş�Ž�(��_�|9��5����Λ�������W_}utF�������@�P6�Lz��'���MH2����)|�@Y�r���ڠ��Q�_�z�֭[��޼y�������eD%�clD��/����"�r�ݻwǣ)�r0ą^����O��_~!��v�sʕ��ېY/)-�������1����b���[�ƍ[�� a�+��13]8T�7��������#��"\8q5�Q-�~�˟��^i��;Y�	Ͽty�Cb�0�z��a�8�ޜ�rz�� F���� N��&�5�|�2������/�'MíÖ�Wo�7����Ф�k��]>���F+؏���#��J>����ԭ6Z�
:9+��t2��Q��^���sd�L��j�����ܿ������W�Վ��K��G�'TKi�z���ы�(���t���.|�`��g)fk��N%�\ޯWk0PԓC����Z&*)H�%`�s��/���vvh�t�m�lr��K�BP�����aS+8�J��y����l���hs[b%0*�ݝ�M��ʩɋϺ��+c?�:]fG�ic���f��\ފ�r#�e�'I^Dݞ�e҂�D�,��uxM�x2�)���A���g��S~F��̒wV���/~��߾y�ʕK����X��D�s T9� �O��ķ:�N��jy�b���`�rgV�q3���P�w�.�5�i�Ց���3���$%����OUc'C(cg����|��)�zW�ߡH�`?Zu�gsQqT!�TAi���銹Y�D�ι�}�L��2Ң5���
>y�\�/��^�eE�"
9�c���s���0�a�򻴹!mpw�? ��ٳ��h@�C�)2��$f���0�����h2�^�K�Q���V��A��\T�$ƃw���<��Km�Y�Kb"q�`5qR��/]�zU�Kr��}��l��c��
�kȑ�����!_ �h�E�"I�k���f�'� V�IAdLgcMܗ_~���+Ƭ)��!����ZũB�F[�,�r�7�x}tx�-���D�x�����-��QA7��9�V�k�v�.��V��a�j����m�xF��">?��2�*nI\�+�	���Q�����D4���4Bb�q6���I��P�b%Y�\�PX�� ;X�d>�_�=�/J�b*�y��w��{=|�pa�!g��9��@��ΉO�bP5�p�j��Y��X���c7�N
�5[�����)����~��P�
°:��Ŋ\�u�IƑ~?ʲ`�m�6<;�ë�����d�VU�EUi}�Qu����s�'*�a��a��Т�"���Q1�B�rg�t�:؊�s)O5L�b�Ѭa��l�9�;L�ٓ��@�5e˱!I/cf��*&u�X �;w�`�T����0=���M����ԛ�22�U���ʠY3��y�\��Ԫ���lCլ)ή�|����v�a�cưu�B��,�0�N�:}���΁�¿�)�sߣY0c +�.1
��:�bV�X8L�"îz֌>�������V]�z=&�1E���/eJgVr_x-4�c��+�,�,X�2Ȩ����ڔ*�������2.u������U�pDe+�t�C+�����K�J�������	W��>	D�+�����]��B� =)7Tk���N�?���&�5��u�\q�] \�ljQ ���$�'Ou����.�zj4[��C������];`�����S��zmk�R�ݨ�n9�b� L��Z�M��t���0
�Uuf���E��%�R�\J8�Ė�<�ܘq�v{4��j��%\�v���,�f�����fO�����q��ܳ*�����l�M)�Y���(dM؏~��#�!?K��D�k3�#J��z/�k�}�zq}�w T5[-Ɏ��lf������o=���+�*Ʒ�a���̨s;�K�i�0{rrZ���!�alT�0q+��ᨯ��"�÷�+x3;;7�Hm}<�$�v��1C2�{~FfLs�Z����,V��'f���^'_z2x����P|���+�ge:�s�v�����/�������UD&����H��_Z[���k7o�'�̵�(�	9�;_�e���n�G�W��,��c����z0v��C���H�l̠���v3��i6F�@��q]#�	� �W)W�(�95a2b�[a@86��(��
���X�m�9����e8�����W�e��5�r8�� �b
���ٳ��'I��Uo�*��B�B�@k�F�2��(���-!>���R��ac�)�t��=��� �۴0z�����Glha",63P��X�8���!;O���pRE�����&R�����92G|Ә8�#F�S�k�rY�ܬ+F��-d��|;��;�@����O~�l��Z�/Q����
gB���2F��MF�b��r�]#�Vk���n_�Ȏ^VԷքT/�A�w��}����	������"̿��m��c#$,!��ǲze"�$�&˰���<~�X����E�e4h#8�*%j����s��9��!�L�xe.��*6�)j,RF�emm2'�ݩ�Khp8T2d1�8���.4t�d0h�8�w��o����s<"�s�[m�n����!�tz�n�˖���d�D��O�o�jo��=���O Ri/��0ƢP,��<��K�:��H�}:7vH�yN$~�F��7�ĩة��w�<,��i�����a@���C��/-k��
�'^\��<υ�:>��裏T�E$���t��<W(i\T�Mr֨�����̄$��љn^��o}�[����=�5���$��d�����������Y�D�����R5Y*S��A�v���4�X�kn��h�B9K�L,f�~���6qۇ��ծmm(YW>JF�U�Lx���	�\� ���>Q�򩍌a����G?���W�9V�X��b���V,�}zRW��!����R�0G��n�H�^%���.�pAD@���+V�^Fyu�s�\V�0$�bG�\^��qVF����@�=�fJ!����B[��wH`E��Z���:}�l�����ث���Z�y���+�7�8�l(va�Ux!k:ӵ�Vu���V����g�]^�5#"B���Y{+U6��FK?W=��^}���Ӄ�E�W�)L�p0VvAV�"��86�c��Y	;�:�W��L�N�VHa��?<��c�>+[������,e�&
���@U������]�l[M��3�1�Ԇ���S�4� ��!?���e�p����������3��P������l�K]_e��̊�7c8�`�_+�~b���E��i��G�
�	��.�!ͤ�Qy��e�tW�M�\�ãG�\���B��iczuϊ��n�d5��,���ڂ�$�f���ND����T,�:�����B��X�V�����t�<7MF�.\�:���Nry��sGgǃ��ν;r�rafyc�~z�aj��_��s�qo���t�^��X�����z�bG%�ذ�Z������AK���>��51A9��ö�����'c��όz�=�+��qe�GIc���F�J�6��^��(���N2_��^:�)����ƛ��2�`8'��j~����)��E�n!��v����Me��" 'q�7�	!����Vۈ��tȮ������+R�:n�/21�j��ř�F��>|�r!�S��M�(���}z�N���Sn˭M�f�+�$�
ť���N�5����av�۷7`]r7�0aa�b:��&$N?=mXEHaggg}}��U1����]g�m��ҲA�bX��a��-�����z��u!<����q3��34\ɳYV�;�y�l�&������\)7ƣ�6�x�[�X�,���L�u��ܼy��>(tj�B�Z�������#��{�ԇy�wY�i�9Ui	��� ���Rmk���i��V�#p���e�W:VӺ!$���9������>'s�pt�M|��D��Df�Ns��Y����N&T���'��ǧخ�'�^��v��3�m\Z���"0��~���Kƃ�;�X���KG�*��a<R޵�ѝ/3�6���v��Ľ���� f?� C���or� 
[F��;�Xf�z��V]��G�lx�$�l%0�c4�	��j�F���
$Ȓ��c��j7�9��h����776(ǻ�A��vת�A6#>�f�c��W�V!-e�v6/�/��8I'�=F{2�W�a�déwvx,8[~ժ�w�~�ݱ�X?�$0������=وq�����y��!�{���b�Z�ۿj7f��0J&I���Jm�X��=�R� �	W�b����X����e�"�����8��R�V4���B1wq^�"y��wqZ+n�r] P�Z�8���u���16X��5E��^�ٹ��Ǯ�"\[O�D�g����}#a�_}�5|N6�ﴻ-g���6�0p���O���q3ew/G�4-D��UF*q��^w�F�Q��c�{IM�~�e5��Xܗ�!��y�x\��_��_):��[��O`D���b%�]V+6Ð��,[�34� ������χe�D=3�?.�Y2rqN� 5��N�zt߻u����ũ��l���V�Z4�Pfz�m��6�u��7�z��ǈ�F��k�dU��9;=��[�(��=���C1���B|�	Ά�Q��r$j��8~�.Zȱ�'����o��YуEX�%�M�q��ds�
8Tʤjp�o�K��#|ԊT:���(z2,�1�"GZD��P,XV�`�c1\�-t�$Q,�$z��U�),��EC2���XP��.S� Ճ�$BΖ�7����.n �觟~j\5S%$e*����櫯�z��-�Q=3g�dזa�_)��Px!gH��;��Z��X`Q�Vd�;V��u(2D�q$�482�Ů���U��FD�U�ƺ�j]����R[�Ҩl��!Q"��%BdMH�w���f��ǰ�5+E��r%�L�����Z�<j���;���"�90~-�W��ys1��yC�.�v0y3M,�IߢӚ�(�X^�U���
v�DN��@!'iI�l|/T�N^��P,�ٺ�3i�	�,�0K�h� Ū����
f��y�Gs|�n�a=U��a=�`ŭB���(ZyE���ǣ-��\��dM]1�5�T����4���h��j��૊u�9E�-��m�H��b0�ijɞ�RPrXq'7o�T�L�
LiU��Lam[<�7�%5��0�B��6�D�B�*���qm�\Y]&p�z�l����eX�]���p�����\g(֌^��WW�8�]�����3J<ҽ�wsf�v��\�Dp`9���ư��q2u�n�͞���9d�$�9�Zv��g7'�������T��1eΪ����{-��� ����u��4��� ��0WW�ggj�8u',���5�[-G���UX�WM�na�**
հ�w0��K�����ϕ�%��c����U,���DA��$NG߷�����kk��^�� Gt��u�4Y���ܹ��C2����H_����߳s�tz��["��X޾��|�^��0��W*�V�*5b#7eA����(�˕�$\�.�a���.:���o�V>2\6���d<��L���S��4z%����TlH+�ܙJ����g24�0�d�V���-\(	�0���7V���e�J�y�F:Y(j�Z��"��l�!��k�M�WQ��r����U���9�Wm��u�s*����(�O��*�SZB������wŚ�<��c�gC
d2��[&�*2�$���Ƴ����ë�x��D�`�q�l6�w��u����ƃp����xHٴZ[�e�'��4��xK/yJ]�T��%)Xo8�r<Jx�(���B{0h63ÌC�N}�%�nh,�)y��_g0��\����{jJ��A���\���b����kC�]^QATZ���p�ԭ.�^p���~�B뇅�l��Óö�Io2��R���(���s{
w�����L�䃌��<K>��)!<7t'���}�T�~����F�tL#���-y�X��J&��Q�&����Z-S����&ԗ9���'=>9fp��J��)ג�	͉�FpXK�e�3|'��5VW(����|��1��r����3T�/�¼���ؗ��lUx3�|�������){w��6,[�C��\[v��׬�y���2�+�:V�^/Q�EP%��j��ٟ���lw��QZ����K���x	�`���j<!�+�M���$�=�E{3��J�H�|���;Dg��`�^���L��e���ؾƖ�sk|��Ǭ�08��6W�0ދ6J���۷�s���+	k�޽{����L��[�\:�Q(�Vـ�(�n�&\��UL��a�KY���q'�V[�-�����*F�j���m�1I��nD��3���1��� !��V[W'�A�M'�d�4I�1����5�
�y7�7'42��Sݕd���]O�_�9�U��-��ux�T�8���>#��(�g��p�5���-V\n�p/IO��1�^�����U{(��h�n�nT��	�x;��U6�������r��`��@�T�nR�CV�aW�%<�\�7�Z6*��Lg7�0��e�%�1�)�qM�TE?���pE����N۰0�\��E�������Q@y�x@����I�!�Q�3�߉���=5~Y����:�7S"� �� ��3�&�N�d풝�뫔2�fv8lj�e-�dcb�^��+�K�:I�r��~�m+�x�Q��ZI�f�D�4�GC�-�/���|<��B�LHa���rE���$��hKk�Ȉ����W1�]Ov�I"gS/�^LЅJUZb)R�Cn�`�+��{����9��j�J�ARE�Pr��^�y�D�5�ˤ?��C���� aֵ�$g���vX�,�S�Z���^3��̫<ef62E6"�ؙewッ���ck�jh��!H�
�����K�2F�8;S/"}���3Z����5Vx������a�X���a�ݏ�L:I:�#޸q"2��X���'$��J�@��N.��yc;����7ϣh��}�m�4�d��N�3x������[�%��L��s�^��R[_�fܣu����.�*�t<&IF}���L �R-���%��n��$@��f���~�5��b����v���Gܹ�Jl��^� O��NM�g�� �j��S7x��y�N5�0i��1�t�����^��B�D������e�y�8�����i2.�!�;�n6�r�����U�*f����1�ȼ���^�����p��C����9�����g3/�>Ɛ���I��-v"�v���ZG<�i�u"��Lo2#�ڲ���j��שZ��_��k$��u)������|�F�*�U!��1��}�X���X&9���l��x%zz�Sa��j`�6���O�D�}j���_�U�cl���h0<�d,NgS^Ա�%��������T|gᮟ_^@��mG�G�æ(�J�JiZY�5Z,~���}��̢d�z��w�9^:RX�S2��b	�p2����8���N:F�ʅ4�d�CXo0�$n�C������F�.n9��vw0%�������l����p�TXu���$|�\[>>��}�dF�<gb�F;7o����f��x�UkVGY�<�����3<�K�� �I����h�:��'aHb�а�v����F.��ҩ��]?l֯�\<�Nv��zX�T��/!� `��W��f��Pp��Ç���W�
����[R�Fh�fr�ͯ�(d�`{�He0���(h���������O�z�8�/��Y�+�.���=ߕ�x����O��Jd,bw��$��ӓ��Ҳh٨�&�g�H��0�2��ژ~�m�-}�Q(�m-�/.
�ѱ�
�M�_�T��K�O��D�ݞ�B�rDX	<Y�>�w����p�X�,Y�YWT�Q槬檱�� |�(��$ry�y�S���FE_�n5�P;c�����.�#���}�ћo�����w���G���Da�	���Q$�q�$H��ɥ�eR	��4�8V˿������vw�Rjw�f��58a�ْHU9$]7gV5M[l:����Z�7Q��#ks��O���"�����O����g]�a�@��l7V��tμ"��J��[*W�簖��ݒ�DF�Ll-Y��:d̴;㬎�k�"�jJ**�pN!���!���^�Q|��t���[YUhKA'�:X���g�JD]����{wĸg�����Y!�E�mui�&���� 9�j,�|���y���c�Ƴ[:;�h�u�k=Yq�`�ꠀ�	�G�t��Y���)(rI�����,MU#��[������*���E�b��5LF��& t���O�J�z�0��d`)��
g��waW����4)ㆀ�#���^���w}cY|V�Ab@�>��߬ԑ�Z���>1�24Mr_�c�������O�IgO��}i�[[���_�?�^�XR�퐳��ܿ$�r�2�
��bX��5j-YJ�tL�|�6�[�k
3��@O`�>}��S��t��͵./R�ߚ���[e�\��I�ui��Q�B�5\"�U�lq�
7@X�U�-ju%ҥc묊郐�?<x k�q�&f$}�N!'A���+������B"�i�����u�9�BP��|�Ȕ��H.r�y�wpzـ��Ev�O��lv�"����Q��\�N��`�g�We_I:�<������hp|y�m+�ld�ӛ:.�����Ɨ����UV]Mƻ����moo��.C~�X��E{��V���OG����S�1�/x��� K'G�g�"�D�n��t&��n�9M:������r�(��8����é
&��Óf��db���l��SŻ��?7�����&�9�g���Lʕl��}��J�3�|'�^67D��cL�_��b�e��������>M�d�� "B�A����҉
3��e����4g����K8}M�pG�q��Y��,���;l1T�-5��ҢT���T��~��V<�W9=a�H)��X��v�l�Mi�2���z���~�<Z_�ue#e)yp{|vy6I'���CL.N���s��V{QΩzo�d>�Q��ق4��VAWa��8�� �`�ֱ��?c4��`cYk]kd��C��w���&g�8N���Kl��_}4��0�%hMV>���m\�bhW!��U�Ѹj9�5# 1;�����F�^�Vk�f�s�R5�����sRF�h���`��'��A5��(
�%�@bU�֌�Ր�/?�<�r\��o���p�X�e<�\&�{��P&��ȃa��2�Je���[�_d��>����kR�D�N�b.��FL��i�T��]���_���'���az��[��n��:�կ81�B��[#�/�P�w�{$~�����	6ݭ�-��"G�1q�%�����z���nݺ�%�����F�Aw���p����ӢW�qX���*���A��Cs^{\�1�2��8.��BuC	aj��ӰB��j^��j�XB�RY���g�v�Z�)ܳV�"���T�����0�~�GC *�L�c)F��$P�W�U%Gi��@H�1�*/����s��%Ŧ�����//.:2�ՔBJS�ӯLI���ow;���8�[̚/Z�ȑ�=�븧O?����I���e�Ӯ�p�o����T9~�bE!�fPT�Qj\\�9���o�6��9��Ds�\r�p����߇��o���0�P�x�_=�LqHQ��
��q!X) n"����J�eԫ���p��s�c#
�Y��}��t��cjLת5!T?�.j�w6�ܹ3��v�@���;�KW��,z�$Ϟ=�B��$~�TQ��l�!.��C�����v�7)/�7L�x+�w��c��kRϗ���:�B�*줊$Y�Fm�n�a�h���6H�/,�dU�=��ugl�X?Xp�f�l���Wy�F^�d�(«��Ç�I�BH�M��Uۅ�\JU]�!h/����JH���ل��,V�z�	�F����/�k+��
�e���m�ny���w�ƃMH��p�͍u�j�X�-�G��de~���IHl�tV�ɛ�U:��?�P���Tu����2��֣1g�9�,c�0se��Z�?�)�V��Ԝ���(��W����߂d$���W1ֺ���s���}�!���̓"��)��j,��S� ������}������bA/�o��3ا\����mD�NY���oh���:�v4����qVm�L��������o��$'�TJRY1�!�O;3h�+��"GQ�T+ӭ����D�d��%�yHW�q8l�|��G���4�!�$m	(�I`VA�N��%�#9��,oC/B����z�7^����f��\���O��JͻA�Ï?����<��R9��>���+�cW)�K����q�u~.���f�w�����Q�ͼ9))����2�v��Nmu��������y#���%�5���Z�֭�8g�I��۝�8W�,��ہ�\�qc�WPZ\]m�ݡH����d��	#E�l4�#����sgsec���N`�4j�w���Ӌ������#�y�lG?�p/�|�*�nܸ�lw��&<���ąs���J�4q`�<�>�-=�e�L������S��x~��ow{f:=Le���¶3^���ݛ�ȡ�jg�h�RM��F�~q|�MQ.��L�:A�@�붹��^=�w�fú�f�cGÁ�ǭ� �����}���� �!�T1��4�������J�X`�q
7ud i�{����q���]��a?������*7�Ɂ�Q�&h/<U���%�ٕ��9��ťj���ђ5!��R䘈�嚓]f2�����Q	��ϡ��9�2��[3ux��̰���О_���n�2�R�.u�<�U������b�>$����{�	I��t'J��씇5�����>�Z3����(ه��"�1�AK�?�ߦ:z�2�$�	���j]'�N)_��N��׷�e����o�����o_�a��.Y�U�P[��=߅yKS�j\�C�c Q6�6�Zx#B��,�7�w��ۿ"����'O��+@�����Q��K�?�����v���,E���o�.O��jcg�RX��̗��K��`@�ܾ�':�;HG�퍭Q�+g�v��c<��|�T�7\)��sj@�e&�nG�!F��r��]Y_c�N���d�tz]l	Ƈ�puPB:[�P��f���듟�X�%0¥R+\�ʊ�bÅ�.�]�\�bI0ܩ��$�a����>�,�3�̴?U�S,d4��ϼy�hh��>+�]/�|lR���v�],1�d��i,�5��m�⼄�$T�+K����@���X[��O�.��������A��)ۺ�!#������j�6�}�`�O�_Td�;�M|%B���SV�,o��P�N�ת^v��싱�ϳ��a���9��kRUvj\7F45[���X�̼��\��Qo�eŽ�X��V�u��Z�hՋ&ΔoP�D���:a�Y���?\Q��U��uq]H��z��c�,�Z���	1��2���MN��Q����ɞbX{�H��=+.�I�D����ƷpZ�S׺�}M����1�^�����o��N��G���8�]V�����"��"T�(q3B����'����&�T����+R|�x�hc��b�ued	*�͸���a3]�d���T�2���6D*#s[���o�^��b����vA�&�8�-S����R�V�D�� �j�"���+I�R��L���Ef&���}��ʆ���*es�F]ޞ��r':f��Uڒ��r9ԋVá��jŅm�X���(4��T�֔��N��V������XB��X�|
/L�!T���8I�8��	3t� <k$,0��ἆ�]Q�OYFM�t�r������6f�����������KJX���-� lll�!Ј�p�q ˑ��I�:����*Y��V��
��35\��vU/I^!nU�;��7�����"�^UP�X'�Y�qH6*��߰)�܁���%W��T̀�r� ʃ�u	�n�hx����BY���S"���No�7d[���n&�y��4�.���Jbu��n}<q���]��qL�N���������vڍ��O���֖B���F����y�4X�?�����A�)T�����3��q-�`6_��1�B�ؒ{�'���N߽Wn��c�z�����*�j�3m��e���s��w�}�ݯ={��ٓG���$�Ta��:I&ݽw��^[�>�s�$���'?"M&���5���k��c��l�,�\bIP���G�U;_,QtiA*�*�x��h�bETsw��]��H���k�*��_��yE�"9�����o��s~�{�K�Cl�0�������������G��ݘ6�Ԇ���-z�#��U�Z+!���W^!u�(�u��o��Ao�-�;�I���G�pggg4�d?��p}{�KRz{����!�?���AP
~-7A��F�q~r
QZ�`��;a�ӡ!�zh4�^X ��^�3���h�9� Rb3�#K�՛W/bON�0�a@S��m[p#P�I�:j;gdTT�^�v6���M_����U"n`�����e>]�!�u:��ˋ��LU�MPv���T@gg4���sDCb\m��NS+)N&X�X���t�F���:A�֒ _�צ5|�tWu�s�4iw�qf�.N�쌂�K��~�ٸh\��>#c�8���mmeehF5��[>u��t��/V�!�`�+��i��Z�L�[�P�^��q:���܍[�H��h*���'q��pا$�&�{��Пz��P.E&���l�q�~29i�°U&�����t��� ��Ü�$�So4Œ�;8���Q&n5��c3粏�<9\{��0Q�h}pUm3I��~t2l!)�!솢C*PI���1��4�}��(M��,KD�\.k]%g��ш�����ûw���!��E2�ִ��y��<��}��o�Y-�w��x�7Z�a��aʞ_P� �pg6Ն��&?1&�ZZa��؀�)dYcm�R��,�u�Ү�����5�1,�ıU���_}��(c�C.[�EשּׂBg���`�S(����ӟZ�(|����۷�y�\����*��9;��Mb�`�Glv2�K�輪�Z���:���%�ԟ?��0> B��4�~	�h�̺�L�}��E5؃di�i�f��B6��j��lg�L4»�����U��@'�/�Uԗ��48y�j��P���ƓLf������lw�x4)D�i�	PrE!o�}획��F%,����=�����g��%��,}��r@V66����4�#������e��6B��I�T�E�{"�/ds�'��v�ɣZ[#ɘ%��n���y:��(^�RU(>�/�����J����c�Nƥ���!�h�xBs<Ty��Q"�'``�@���)�ƶi��P�qY�J�(���Ή�T����S�N�9�/HÔT�@p��p �$:^ް�Qa7+�ak֨NPm.��x�l�:n�M>�P��F}I 3��b�X�j�,9+�4�+�5��c����~4]ȅ�������$�;�?۽�5ŕ��
��竁���T��U����	�m�������3v'���"5(�K�^��9�}�k��HV�Mď';X�^B�A�j��I>�}��e��k�1��%ӅoĲW��1Ϟ�`��\þP'Q��4��d�=!rd�0$=+\<�.��^`d����,�2�䆦[N�6���ř(� �Ɍ�S�S�s*א�1�E�#:vk�:�:^Qp笣	��Ӻ��_������E����y���	�/�F�"�v�5WY#�E0=<�s��"�2�1�����W������Ý6��i��/.w�o��0�m�e3���ȇ�3�����X�\N��f�e�ãcn����E1ϊV�K���$N����I`FX��qvv
u����vm�Na1��R�*���M�+�,iL�k�T+i�D�--��+�ܺIc��c���M�%1�c@������V����n��)�T׉��k��T����&Y
�
���;�b���}<E�Gf�`W�l�7w�s�X����f�8q�~:���n6?{�l2T��'���k�|��R8X�,������e�?y�����o����i��''�1ٓ�I���L6g�j�+����uL��
iD�Hm����p��LQ,,��?�����r�v�S+02�p��޳�a��G�Cl!ţ���~ e�� $Ux�\��c�^�s�Ȟ�[��ڰj[W4�����[��\,	jȘ۰e"�A�ְ#����%1T��0���p�TG SEh�a%J*A,�)Tu���N�#�m���vvr�0��C�^�N��e����N�M�fk������l�;���˗�ǳ��8��� 5�6�_�B�[�t���5Ȕr�+�ю�,��l�l��ťvƖ�i�k� ��K/� �:i&�k�� ����\��eJ��x{>�
��n7ȕ��5L��x}�I����X3�w�'�`������/�0F��L+H��]B�V�Lz˵R�'�Lm-{vFYl�'2�f������<�����US�+��I�VWmeY���%��lehW�JG��V�M�Vt�h#���Ѱ�ˆ�7����q3�!_�X\���ԝ��\�MѤr�D��4��{�4�Ee���h���{�����s�x���j\06Bb����XVoh��O?�K��k��X!��e0Wx96����%g�@�����G1�'�23x�T!�1S�&� 48�ͧ��l�F;�%����ڶx�ꫯ☽�6K�R���(���s�|W�q���H��|E>Lx9?��O��T`���C����8���e]b8�0�TikC�N��NU�x����<xBX@��޽{�JI�wq/cC��[o��Ax����}���t�((ת�w��.��zڲ|Ǻ%c
9��l%�Zs2u5;��,ׇ-��>FRF�`����� ��$X��s��-� �O�>'+p1�3W��1��d8x��7�7���������c^NN΄Qa�B�+�3����d���������?��߫F�1n+SW����A��;���O����E�yŬ̵�Y)ӷ�Mu�?����HA�q+L�ι��������1��T�61�u9�2؅]�l�&�N�w� |�0����gȥ�[0���з&���5eT"c�}�b����Cܫ�X�m��S}.�]��+U@
aG�TO��w��<�R��hn8_t�,���dtI�� 9ӊ��f]F���,�jwڣ�X���Ԍ��S�g��8�踆P�8 �p�ݭ㘖E8d���˚r�8gdu`j��$SM��jRm
��^Hحt�Ư����<��?o�G=a~� ط��E��zk�U2�BE*�J3L�iC?yR�`�K��@�8����"!�����oԌ��1�E8��rn�P��׵9�-%��#��*�ɿ*6�����Ǆ=�F#8'�@���7��*D�N�K/W�}Qm��*��Qʑxmrb����,�w�X��/�]V�)C[�A��ƅ��i�4l������{��(�b'������c,��6����n�P�f��;��i�c�7VV1x�N)�81�滞�P�d��ǅ���f����A�:����C��������p�&C6d��)�}k��嚥"q��K,kj���J6_S>�q�s�LG��v�G�I���I�oY�$pa��\������w1ͤ�J�����G䚽�0��xn�w�].��3�F��'�f�Bc��d8j]\�Z�N����G�Ǟ6�^\�X��ۙE�(�{�Z#W�?"�yLw�[?8~
�nⲪ��u�R47:�2@��/#�������o[�l�(�!y��W�ܹ�٧�$b*�o��0	�VV!vU7����흷�~��w�-�h�g���P�YL�\x�� O�O��xVt��uu��Q�*.DG��񱍭Ṃt�O&f�4q�������B�~~!���B�������*�0��)�������uڇ����=~(����0$�c
E�E�~�s[�k��)YY}=��	HA0<8�U5�F#�����i�BW6;^ �:���\�V�t�����83SA�L�b�Ɓ�ݬ�U�����TZ�����кf�a����e\����]����<""s��R�˚�M��qs2�)�L���D�U�V�s�t)�2�vk�Q����S�IXF �ٟ~�՜�y�B�M=�5�7/{�!���2�L�l��3���E����O�'��k�y����y
q�m��4��(�y�Z������Q�t�n��ٮL�,�|��I�\�%'l�O.Z�8�M��l@�F`�>����2R���\`�(��n�y�\FO
4	�h��6�$V�dk�6�X��-�ׅ�����m���q~��ըTI8(	a�ի�V-���rs؃����­�T0sKf�ʐ�E��*��L����ԭP0��.���]� �<�>T\��Hӷg��+r�/���D�_>Քčn�8�s�wC��M�����$��q���Op �rG��F[�0LY�X/�,����X/�j#ƅ=y���X'������dRo;.m����{2 �-C7�<M������>��s�Sh{���>e��$��K���
�"��ڴ���B,f�hS"T-Te��֔P	�8_�#��q>DF����D�I�#�B;�Pμ��b��m@�uz]���(�\��Ww������V-������ŕƴa���V�' 2���)�q�y��$|�ݧ,~��1���������󅾄lR�T(8������qB��V�0���ygX�}$1\�A����*傰�f8�m��­��_�E��<
D���1�KK$bR���(�(l]c%"ǢȂ�F��T��S35͊��W��̄��_8�:.��ċV�Z=!���Wk�M��!,��g�����eF�we�+x��������&�*T���_�>�*�[*���^{m8������_R�̵��|�8�$�c�ip�L�F��1\u��L����_*0�3��jb�����L,����itg�Y�K�\�	�H���C �"�eAcϥ3�+n�K��}ג[����	���+�u dֵT�2�&0�6kE%i����O�>�e󸫋ibaz��_?MV�'l�zz~��o8%_JTB����J,�nsYkJ�I�ׂ�	>�0��8⟐�05�n1��	T�L�7�b���O�����%�0��U�����M�������z�@KA�������ț$�o244`����jH�؁#�:!��(�F4ǃ�+��������q���o���=�8�+"1�6qb�&�-3ʆ^�ͼV%����7��矯,U��8S�v��7�����n�R�\��+���˫�~6�dh�i�e��!Ev�T)�����Y��⠳���V+gX���p�b���ʇ�G��#�Ҳ(��J�Ӳ^��Gd�6���rd��~0T��w��0��ap���nw�e�=e0}�q�0pR��YUc�$���t�$�Wq�я��$$^��s��P�=���˵��6���i.Ҍ�z",��x
��C�榖���[�ɼ=c�*M��F��,)�ԷO��;��e��}*x��a.j��L�	�&Fb�:�ę�1����Ba���*���a�C�Q��������������VkX��\�-W)UW7��K�NZ�֨=��b�D:�sx/u��f3���Y�v��Oɶ��noecsi����b�_�;��r!�u0P T�ܽ�u����dgXFV�V�З׭]��Aw8][�d�x�����k�����2���ä�:o�s$q�����k�1����:�FQ��`2)5=��D��:dI���(���V�	�Y��N����r�8�"eή�����t�\\�u���~c����LL�`�_��Z�Ѭ?�g=׵�TpV:M��
v΀S��'ӑ9���-V.ǹ��d��ujk�b~�B屷���w�V3q����P���s"��L�L��.�4�Y誽4�%�0���H�1����I�!��H|������`��T��"�9Qh�gO��9�^���dc� x��,���V�5�!�x�T���&f��u�푬����Bg����Ԁ�tD��t�(��ƹ����c6=?8�)֋[l��EC��������7�3fo^[_c+����X��<�(Δ�LZ���[Z]۹q�̤㤶�	�����i`9A0�������ʟ=~�xlV���r�qgHR������`�z���/�Rb"�ĚMD׶n`����CJc�<�<��#����_���i[�C�7��_��~xxpz�l��8K}i<M�t�B#d�l�٨0����_��n�i�!lZ^N��=��uz~@w;���zf9��x �-]�Ns"�)���ƨͲp����S,c���d��flw��\�䳺�+�ϲ�NW&ԃ2��j9�����W�jaa|�-ќ�L�����؊����|�H�_��7o�Hp�"[7�����ei$�=��x^���[�ZŨߒ�V;��L<���xQ����
�*/�S)���t��'�--1k�����w((�~�zT�7������|q���M
�8�e���C9!�o�^�Ҷ�U�>p-\v��Mh�?��?|������[,t��;}���:a#؏{{{����)>�K������z||�����eCp���وx6�_�+ى*�T"�k�K�3�&�p\b�hI]ڰ�Ti�sc���J E��5N� ����k7��϶���K70�1\��ȵ7�����\�6v�Ț7�bF�w"JPM����Psy���.�#�g�Ւ�,]j�O4&K�^�£�'�/������?���_X�"V (hsC&3���b⦊�j��s��^���sr_Y�D�3ZH�/�-gނ{:'�Ӈf,�ৰ��B�(����)�p����Z���J'�$���M�b?$0��>�#�Z�{Y���9�%.�E�&l�>X�EN
��7���?��WP ��'�+�ٜ����3≇j�����Q8)�����S�wa��8��38<B,X�
�0��n��*Wp$�ƣG�<k%��aa?B�����
+OSlsc7����ࡰ+g]B�bH}q�s:����0���s=�?��ŏa�Rۼv��g�{Dy��O�i�LqU�v������ܷZ)��qg�����{�;;7'��6�7p����� �3!9���\����ԛ�m�S������g�R��)q?c~=�&/Wj�������o���Ak�����mX|�f�\�he�r��ΰ��J.8��!�SR���S_���~����y��m��p<��߷��DSk�	����J'�)��@A�I�p2}yxp��;sq���g�ˑR�&�M���F�ajp��7�,)\X�����E�84t)�M\CS��Լ˹Z�ƅl��<�x�j��5ͥ�=���Aؔ�y'%��u�1F�V����@�g�������x睷U�{vr�u��U����}\k;�"�O�Znjh�h���#Q���1���=�]}��7��k���¢�'�?<$���P�$��^��7X��{d2��ҩ��?d��#�C�o����4M����0WȲ��d(����6�tmu� ��q�P5^���J�X�ƛ�`j�mH�.�Z�0��~.j�E�(1ܩ�P����Ijm0��/Ccd�P��Ǹ��sT���ӳf���r!_�]���<����~oԃ1w��h���������)^[���ǟ�Qe�DM�M�X��C�i�v�r����|����7�S8�6��i�O9�L^��[X*Zl
z,���d�/_F������[�iaN)�&�iw8^d��
&��$�dDu5��my~υ��SǍSRWg�I����;P�G�g?�я`^30�C�4�a6�w{�?��$��TVn/���(;���`��R���+�J�lϱG��l���W���?�����v�����T�ph r��p� 8��3X$�My�r�.��mߺ�}����>���3�"[`�Ƀ0sxtb��O�~�]�닋l	L�O��r�	r���1�GkU4���z�
����Sao$%1��M����%�.��@|�ls��( (.���]p�T�)>(��I���bGA����J�C'���[uū�����x��w��jW&-�_6��I�f�Nǒ9�;;����޾w�z	��X�1)��V}*k�rz|̀���2j�y��6��.	w���:Z��8�1��I��L�{���x�-H���ܚ���e���Br_�F��0m��m=]H�����R�A��Ɣ5�V�1k1y�1�JX�?��?�-���7�n������_�V�$)�h`5r��{��^'��(k�&�ޙl��2���}{�̀�N�2��P̚�c���z<�0
� �Y���@ID �`Hi%���
�2H��i{KE�7e1(Q�s��`~3����AI�J�d~�v���%�В��LiN�xp�\Dg�f��jKJ�(&�|���D�u܉���䭃/��A�b�������;�H���Kv���w��ڹ1s4!�}���O۲�iA���"S%��@�B��5Y��z/E����>�w[��0:+���Y���բՒ��y��ͬ�w�*2 ҈
&t<�q��L�4�v��̶�R�x�88>��+Ex��Y�c�,��ê������%�(d��Ǐ_�[��ACyJz�d2����Y�CѸ�vʵt���[k>$�ꁄr$�(mp���#z��*�q�P���\
����|�? �?��R t:p��2o,&�4���`���rb{{�J|��`�7����O|~|��mxq�����d�����p-FVI5y���Y}rn��_5�Xo� T����A��sfu��+5�P�{�ԩK�˿������4]��m);�ib��ҍ7���g�FOt��e+8L�V�����r��͛��Zb��.��a+,F��2�L�`!΄�kXAUy��x�lo�%[�ܘ�K��b�/��6��y\ok�B_PŰ�K|y/�N���k�����V;/E����a��~aX|��u����1���rdb4�}L<r<y���h�cc6�}߸�<<=����O�������?����_|�vZ-�T�9o%���<�H;:ܺ{3��G�$�I6�:]x���%��4��3��F�޾�a�	.�5��P�ش�����{؁)��6��jR�N��u�ZAhD(k	���D89f2�������.�^%��$"��ё����ӌ�ʕ�R�F-r�IٚvH(HK%�FZ\��F�����(�Bh��)�Q�V!�����{�n�n׶o�[au��������w���w~����ܾg:��=}��������Z��pM�C���S w�X���n�em��iٸ�����s�{��O���^���u�O\�_=�5��\U��-;l2���0�������s�d<�{]׼��:�ۤ�/�+��������ޓg�����VW7+i�wr~�j����O�������89g!� e��=%�1/R�f
�8�d"8sg瑑�5�-�������ϥ6<�Y�Y^
޲qB���X�
���P���z"�7r�5?o��񌊪��4|d�0�&�꒱�43���t2p`Fa�T�R�3�	v/���:��{�7X����Q�������z��G�bN&"���˨~U��F8P�m!d'��
?�|_Y��2�{�T��
	�M8蓰^�*�w���*��
J��	�ɯ�v��~N!UQ�?��6�z�9��� �\k�H�h4s˫�ڨ��gh�[pE�����\�1�!��=�g���1䨜�s�@,���\|k9�/'��.^�>ч�Ě�jS�8�i��(V��#�/�0}������3��%������ۛ׶�y��=��O~������˓��ٟ�ٟ��׿�G�G�(����
�02%`��ط�A��W�$���/T>Y�	��	�.
h����KI�x�?Q��������6�������܇�'���GP6UnV��fc���B� f�vjM�t��J&t&3�g�$G�-�^*�a��f�!��
eD�ڬ�4}�i�Sf�Hj���R]�x��5���@Ly;l(l��ʲz�M�^�{�]����o��\�g��x�f��Y��V��ò��W�L�/��/U�֖��}��t��}���N��8���d�\�Vb�����p�͊S뙰�S۪�-{*�(�E]�ƞ���δ�+&���px����K:Ow����j+*�7��'�	���>���ٞX����b[Z]�� Ȱ\�M�"��hJO`6�h�1��"X����38��9�A1'�ɅZ�0����I�7�������֧ [��V�h����<��S�v9��pE��_���Ig�uW2#�N�/�ؙ����F����5:Q�f��u墱*歫b�1��)�5������Q-����P��T;�?�Dn�R���&dX�� ��S[���g���Uφ��}���n�^^��gk�:�\�Oڢ�a���l�|a�J�����(6��јP��Kw��aU��S��ٺ�#�W�E�X0�/D��nZM�O�Iگ����G����W��eg�����a/Ι�Y��	=e/��lDV�0������[w>��Cz����&�v{Ϳ���tz�������o�������q&�$ͭ�f�>ˬ`����MXkvsg��?Ƽ���\�8�?FX)�����ىB�X�`�J��Z-$���_�Rf��Q�mIEq?EK�f0�AS�ز<C��[����фT*U,�,U�'�,��������9V	[o���Q+[l��c�3�*�T�c�F=����1�������35]�b}�!p�^�) %�/��=O�i��+����� .p>ε���{ׯ�������v���h8�d�/�)�^ ��sf��1]8
s����(��������dƦ�:s�b-<��/b�f�翴j}I$���Ss��y�8
��M�Aq^�Q��m�H��LFp�l�>:��WW�z����	�֏NN�����v���d<m^�����y�����Y���y뭷nݽ�}���þ�~4���0)#K�Cћ��T*�-����\�y!�F+V`Y-���[*uQ�L���ی4~��N:ľ����{���h0TG�?��VBkO�x�6�.-����Z�������dw�2��T�1�/^���!� �gϞ��W�R��(�/�y�+,@�
����2{Pc;a�T4+JQ3����qЂy#�y����b��$��bP����{��)7���	��4(5�1ʅ.ׯoY�A�fcn6�y̞���ݻ����31y��\�:jK/"�!�Zo��:�X�jD�����_h�+�� �����o_D����_~��z��_R9�����r@`����_
[�~�yJ���03Q8���f��+������@���c�����o~��V�����վXzo��LiE9��Pq;�Q����X��L6���F(����J�s�|�Tմ�y���pb����o͚Ty�Gօp*���*�2�9��pƥ:�;B�زߊ�`US�KT��v`��O�1�;�m����c̣�-�%'0��&�a�\���N�#�R��N�"D��;�Dx*�@�3��с�ȴ�X��DY�}�_绅|�5��n�:���{�ot�~� �3횞�!�>i�,�w^��3�|��j�{_�:��</��=�ҩ�"�8�c�`�nʵ>S3��qn��{㲡��c��(�`A������
?���{X�O���?yy�%�L�����c��{wȌP�Ɵ|����1*�j�f/����y�q����*���㊡�1eVZX���]�� oU.JOŝ*�퀵�5|~F��7�7q�����Cܻk��[����w�����%}_�`�ˉʡ�I�m�V�P�\�b\�8�1��{tr��S���'�$�j���e�������n���Z	���c���F�ɵ�쟃C�#���6���f}m}�?)�s�AOA��g5m����'O�1��R�כ�I:��r�^�V�~c{s{�����U��{���x2(���I�3~8�[*�.�f謶l�G����+��6��bYy��Ck~��o�R18_�r^��KǤ�v���/�g��v֢U�O���_�I�K�(,���Vv|��[�*K�����o5r\]����gw����Zǜ��ֱ6��s��(���{a�	N9�1����Z�»#����k/XQ�������U�܇u�a�'=~��|l�IY� �������Ź�*r�'�|��;�=Z*W�Z�ʠ<�r�Ĵ�:�3,��$�F��T�v.᪘��������3���M����f`:���i%�!�E8
����Yt�ip8����/��|K�b&d$��~i������k��v�P�C��G�뛛��;���/�XR�Kk�%��!��{�N���gb}&�=�E���Je����?�Z���K������El�s��a�{,/�UT��}��'P
 ".{�����j!�������'���dW�X��K˵(�>~��O>��_����o~����?��O��_�����]���$��G�ӳ�+�Sqz��#�T�^n<S�nv��E�T��j!��!M�_��	�������5�U}}�ƿ�W�:�O��OYtn �Fâ��I�ك{�����/���-���h���N}�5��A0C�K�^);�K5 $���LF6Oke�����+5G3�ǰ���O!2f���L�7"[�� mu��'�jEj��͛�6[���l��P�V[��R&L9El�_��☃^�m�\��u�P�3RLU�u!ۈ��ckl2b��7o�F#T�`5���f����Z�����/�ӟ]1-���֩b��uÇPd}mC�3!��FgA�T��D��$q3���a���QA������2Ķ�p�U��%$�\|�F,�f�-� �H~cue[iC:		�e�Z ȟPm�u�KU;�����9�N,��H��s1�([
'W�/�v�9�-5��zf�lP���j4����)�V�����gMNO0b�^�x{�������w�[)�������8a
z��ߨ.�bm�dʁ`��4O�D���|}c����{��!yN���$��B�m�D�%�����!����au�5rkk��<mKs!A�)�)F5���$�k�:��#R2��_�����LW�l������P��X$���Y�ҷ%�L0�N���Ee䳨�G�����2�Q��3�=����a�k��t<�LͱҒ��#�-��$�L_�O/�B��y�k����nO�$+b�兵�W'Ǉ������mZOg�����]�O>�L<j��0�5��ʫ�l����̃a����8XH�j��)U���29�7�,�@�V���G��K+����?���k����rrޱN�N�����8�ݥl��o�s���Y~�����;;7�w~���/F��Btf��<���ݹS('�1�]��0�Z-,3�"���9�w���c�:`q߿�1$,��Fl�4����Zې,�9=%����`�-h���ą�Lҳ+�n-U��8>=}.�f�a�]��c5y��٬U�z�����i���Y/hܒ2�V�1]p�)�"�TyK��Ҟ���5�Av�L��
�1Z<]�9��>������b��0�wyy:�m�]�n^�x睯A(<~��l=����һ�{�Z��	~i����Kk ���{�g���\l��S�әG �`H�3%J��+%����r\yqխ��Ȯ��ŕ�#W�rE	�H�DI 1���S��y�S���>��l�I��]*��g��o���֗�
~��i������h���1��0��i�I/�M9����2��|fo���z������1��W�^���9��4wl��q鶫��Jo��f�+|3�8�{��h��/l���pn��U�s~����+�
�U���H`�JW$&k�1�bA�>�l^hqZ�L2��8V�	Z>�t��3�~�T.�P"
��t6DX�>h2M&>Dx�G���C?�(��+ET��
zwgg�#($Jh��אo������͛7�u�^�� �x"���\��i��dh	�[U�"&��j~m,���!+!���Wq66d�x�:��ED��9x��s�hP�+y�lF0΁?�����鱉��8S|<�fB�t���<��'6l�A�8ն�##'M˾w���k��֨�!QԀ�Cv��G�"����)4�}ԑ���P����-��?�i��,��L��B�[-:,�J���m�n蝰 �����X
���H���Þ9u
�mik*�F=z�6UQ��UBk0��D�dR��z��7<�5E�����*���,~�()���:��VACq���ʲ���%|������a��!ꬬ2t�._��|��v�2���M�t�
$O*+A�=[�����?�����|��#=4�B��_��>|��W��e ��E�7FQ ��eI�F[��m[��p�8`��;:� ,�DZn�QrV�����9$�*O����!!T���٣��
8��x9�'����d��	��u$?��n��r�^�'r&�İ"\~��m�a�3�~��dJM�d	d�T�ܹ3�F���F�\X��D�%X��/�l&�b���vۺI�Ζ�F�G���I���V��4�)䳢#�bd~C��KE\���F��9y���S����@��9�sO�U�'{|n������S�lw�ɐyU�y��n���=|~��=����us<q�����vӑ��˵j=;=���Mg�ܹ5??a2�9B�c5[��e�JE?�[�~&]�`�)���:���ۆ������������0!͆d���ft&Ձڌ�ɓ�o8^IfD+W&۠F�7����1�`����S�ȑ�����$�<x���)$��j6�-�՘tz6LX�R Jîjp�B�h%�
O�<��R���=���n��K��x�|���p�þ��loo��0=|f�����ن�8slI� B��Ͳ���y#���ySß[�?�4���G� Ah���m)�Ƒ�Y�a`[������/�M����{+w�@hO./�\�z����ڟ�ٟ-?�̤k�7��zBoT��j�^ۓ�ׁ����	�±F8�w���P�GI7�-yav)!�������"d39�r��E������Dzym�Nt�����A876�8vM��X��X�� 'Dp��l�"�����ë�Z�#̋s�H*��I7F�,,�������غ�J�`*<�t*���2B�E�ݧ�z*�Ks8������=B�zs�$l����������Ԏ�c�Ј��Z�*��sO�)x�L�SN188���p�\*�a,�9�v`�,E��G�G�c软�ϻ1	K�O�"	�66��^���x[��e�Wd]�J9@FA���.ŞN@�$�����LN*"�H�s=��I#R��{;�ld�1Ex�,�qh<����uv�Оs�#'fc	p���.��ϐr��p]��@P#G�2M,�i�>� ����A�1�c,����
�Z���I�.���&N'�ő�S��`'if[2l�(W�����`�K�.Y	3��S��ۿc��<�Ӗ$��h;N��b�g.�Ġ�7j��T�矇������X^:���}���Xd��luhD��u�+�{4���,6@H�)�&�Ì��8�,CXZf��|�ʕg�}VFnך���[f��۲�$!�[[�j`W�����J}�(lS�!>����NK��ZM�iy���Ę%i�Q�[�f��*�L�0�t� �8��^x��VH��Q��K�ɫ^�
���K��-�0Klmm��"��nX ;�����Y�>���Jh����R;��:n����i7�P4Q��ڨ�,3����|����g$��٦e����0�a��0�'B�������GO_}Nw��� ��0�Dk�c�,���9,��RZ�!3d`-D|uuR�M���M٪4ỉ	Iz�����{�H��8�o��f��S��J$�c�N@�5���֩F$"YI���F����B(3d��J�r�p&� �7��yff
���N �uK�"�j�<�����dӒE��!�� (��-4��F�(p�X&����h�|h�`q����eD�h-8�G�Á�(�����3g�{�t�Yc�%��b�H(B�/^*e��qF��X�7��G/��W������m4̣�;�y�jC��?u���eZ��50�E�;���#��l�~�����̉��ۃ�>���07���z�֭��uH�ɥK/���ݻw��v�Ƞ.����aS2��h2rjj^8B���I�Bsapv�INCB��II��n���¬#�-�&��K�L.v C�%��-�p@{/;�v��m����Vyl���E�3#��hXa���c*�8Mu�^��ɰv���l��Xf����}	�ԇ�KKP����A�alR�u�=丁�'q�����d�t���Q?������l2�K�I���\y^<!H��5/J��~UH,ΜZ���v6�J`ź�mC���|JG(�.!�����n��I�Of��,<��m��uV
l?GY�}�r9:B�4�q�Tī����aO�T�E���5��_^^&u�Z2�=��Q��u%o��m:L�G N�KW	�CI�0�NL2ф�K Z>��d���CE�}���ē�9o�t=,����rL��d�xa҆��a���VY��P;�rV����,�`�$�M2r�'�d�.H_���y�P�����a���[\�3�=t��iN�SK���	�ʶQˊ����XC<�k��m�"�֥K����:��ӹs���?�q헿�%�����C�n޼ɾ}V������`@��ۓ�$��3 �dq��26��l�k��݂%i� X��C�$�={�l��$����
I���F�2�3 ��p������m�F;v����o�oᬅ�T�8�3�(����L���!%�lZ0^�v:���,�ތ2���?�?�i�0àW�d>�� !�Y��9��މoe'l�7ַw�dj"�Ó/� �N�==;C���ۃ��5?1u��� ��lV#i2J�$L;�����ϟ�2���Qw���_C����lʻ��d��!^���f>�ſ�'�����;�>�/�5��ś�ZX��ʧ
�r�R�]�q�k�<i[^�����(���w��hvv�@ح��z�.Ҷ�>a��
�(
�A?\Z�)���^����؄2�����(�'&�p�W ��g���i[��c%@������l*��q�Ɵ�������[o����J�OI
!C�`�1X���b.�<�H��IrI�{\jº�����U�7�vH�+QN���3M�:��ڜ�Y�Y��&�e����_�à�j�� ,��ӳs8ݽ{�z����NMNN�P͚4�
�V�1(��#&��Kn�Vqa��Wp�d.����>#��7��s�	I���YY���6����\����g��~��ng��ɖkt�Ǜ�C��x�Q�L�?������x�����lqv��կ~��G�^Z�Ξ<1?}�گ��Ĵj��c���~��^ؘ�>�����Xq*�d%�*p_�P�ݾ�>
J�����(���Dh�#軉X�W̫f	�I�\��mȪ �(�����,���[wq����h��V�p�(F}i�0�B���K�z%a�����&#�3d��G{
r��}�ZF$�˵;qzb��|I�z:
)��/$�;O���L�f��Q:�0&�	0օC����ȮE�XW ��"�Ζ�BC���.��JY>�a|��t��Q�|�}����6B�	XbP�.k�pMA��͙3gf���{�=���o���̌�&HBVA�t:��d%C�I&�0u�K��W�0�H����ĉ�E8��B<��ێ�p[]q���E�_T!o�O,�jeW����q��bg>��OM���[+++��[C(�r��"��3,ig)0{H���YG�Ҵ�K%=��L�T�_��-�2c@ba2�g��8"��1%�IXa�^��5b���"������S�w?��t�/���/^��>������;��.���?��ު���$B�i\M�R���k[�8����,}q3�<p4BfDI �a(c1���e�"����^Na1�"����X��2huJ���G��Z��I��aߏD� ��5�ͻ^fiyy��ʞC��Ib�0kS�l:�i���ː>1z�A?�߫dS�ٚ��%#[����0�H�Q'"���f���R�	��D����I�봻�Ss��z�[_9���/��ŋ�'���z�ׁ�r�rq�� ������d�$�賖�Or�>o���F_��H���t.���+�m�FFx�¹J�Zݯ 6m�:��R���a�}Z� �k�)�P��ݑ����l���R����Z����w�҅��e���G��������O ~0;�{����THIM��+/��vl,ږ(��+#�_�p��'7o�c���"ib��9x�^*s��Rd����O��󠜾gD�am�u�+4i2�������ZO��3s�B�Hy���A 1�0౰�I��'Sj���/�^J�%v��O������l�>�zF�צƏ������k�
剧�OU7w���g[,{'O_X\>��6ᅧ�LX6���@��NYRӍ��2̆��fǵ\H��b�t29V&���(q&7�A� �3Ns�u�V�ن'taz����8ޭF$���-�P��v"�����"e�|Hi���g��Ԧ��<��K������%�S���-(zAǇ�L4;�� ��<�����8�[�B$����\���hLC6�sZF' bYNE�q�Q__���=�$O�������j��_y�˗����ձrt&�����n#�;j+ۻ��C�����$�A� ��988x�E�!y��-xd����lF(�{���k�����JrDu�T1;+E�7`���!���Dq��۝&LHBX~3�8C�3�%�U�E(�N�<���ٳ�o߆�2�ˡ�c�e�_�����SS��U���u�V;��������gb�8����
��'�ɑΣ�.Bs���hƈL^�b���әl�(�#�#tK�h|j|�[����\�t^�/�|���@�V���7�7?�����O�
�y�&]�gO��>w�d0�̔�'�w��u����Q��|�(���9d�@�!�(��]�-�}@J!G��^��h{2�X�I�׾��Pg3y	�]�l�^��\��f��!�c��'��I�80z�q�'b�IKf�Z��d��%���lZ���$�a���@M����U�X���,�ˈΞ9�ӱ��,�p0�P��S����:���%-�WWW]��w6�8�d���;c���>N$k�LT������z�Av��%�+CC}���a��)S"�2',�w��V o8Lg� Y���z���LC-�݇�%��ݻw���x�z299U*�-ak��R����$m,i��J!�N��,�hZ�t�B :�P��Z��s��Y��N�X.����������|5B"t���Y���p��,����)؛�++�;;�奥�{=��d2R����?����q�#��
V]&���B�F�%N�}J� �&��+������冣5�!aI�0~M�N�kY'�w	I���oX�^ބg9Pɔkو��5)2�H�@,����dr��m�����S�,~��T*��m'&���/��曻����/-M����n�z��g��?}�Py����%a۝�x���p��=����V��Z����l�N���Fg����^�a&�ӥK� rp��x� ]�~�����ڸc&��ju;�B:G���%="E��:~?0"���ar�Q�^(�o�һ�=�r��BM��K�e:G�$������K�V#KR[���E��B���t�ɅʀY�2V�c�C���K����>��'Oǯvv����� ��ַΟ:�)t���}�/kQ�򑻎p+�����n5Gpw�z�4�M&�c'`n�g�<j�6��	)YK�!I���e [�9��4�X�2-aVN焮�V���v |�������	&J�Cԗ�i�C�/�/�
��^�>28R	��8�՜�q�taO/%��v��������̌�:]6��3�ĎBCtlc����1h`�a�7,�u]�Ĉ�T��ı�*��X�PzP�~��=6 V0���/;����V�W0�	������K/�������x���/��<h���G�y��W_}���u�-w����1�&�/���G?�hhS]=hj�"/�V�S�V�9<Im����)]�ڎ*�3D�>;!s*w7%�?vB�j+���C[�qI����D�s����a�Ү�馲9�q���P(|q�,)$)̙����!Kd�yD'R�\+!�ֽ��T�H��>!e�����Y8��ζT�k�l��w�ֱT��2{���r��o<���s����YoL����w��+�|��Sq���J���rO<�����jk�F�ǿa��N|��!~,�2������s_��D��k��2F=�ԩd�����m%��Q��rY?��#�+��W�Z(�}>���1i�U}�Xru����+�V\=�4Vf?��T� �B����U*+C�fg�dd��U��U-Qnl��j�:Cx����6�����^c���k-�;a��`f�K%[͎��p%�b!��"�ʚY��D��%�����n�� ��L�;B��H�z���<����Ă����OoЏ��B�piHpd]ܝ<���A��n���Q��q<
��G���7���a|v�b���>{�\pq��. Θ3K��s'f������j��|�W
E�����������w�����de]�ɽv��g��R�L��!�Z5���ujr&
�@�퐂[�����.�(�~&	X턃OFxnB�Ed�^n����ξe�X��uԨy����0�،�DapDb(T9�P8DoD�O,|J�+�ш�/_�������H@۔F�������e�������ζ�'�E���X:�����c:k ��F'$�F>ڋ/=�#�<�S��x��/�;cH����Ң1`em���9����m;��p$r%��׭"�%�sܤ��xKKK�_	1���e2YR3���055	�ݱ��r"��� Dl	!%<9�D������Ⅵ�^g:�(���n���2���ݻ$�Jg�y�3jt�}���Q,�;,`�.����ϩ��uf������hx��d�ۙ찱��8���2!�$i'(�`_���f'''q����d;0D�h1o:\9�ϐ��^ YX�'Ǳ|}��$�1�	�Ah �D���?��{7n�xn���`}}����������M��Yql"T���E��Ey1��N�6��`
N�n$�����YRD*`��?��E�!�����vd�������/�8�b� ���X��O��j�E�
a-n���T�\�����X�!}L}�~��t��� #�/�M5�(-G^b&��� �s*��>�Ú���a��4���lc1�:IC�����RY\XN��8��w�����w_�f�V����V��q����k�C���\�D��ala�fc��<��q9"Fz�ᬷ�Ϩ�w�q��7���|j��迉O�Ѝ��#=6f �n$뉃�n��g*��p�͈��h��q4�`��p��KS���8�����n҅�b�M��*uǴR��wz����gA�ĉXB옃� Ѡ`�� �ѨC�''�vtc
�C�p�vUh�]�����17��l�Yv&X�d2�E�C��6 
�CAڦ��\��͛�b�|D��j4�;�˃�Ǘ8������o�'בAR#� |X:����Cȿ�Ϥ��W�q���sk�T#cY�q�Ĥ�P�s�=�ڔ��0�X�&�0N���"�E^2dZQ�����0��������]������8u��A�?�	���g(H�X>P�y���J/;>�ū��K�����Og���Gߓ�e$�#�H��?��b��f�n~����)�� [����?�aa��O��N���s�Wo�}����<�?��?qݢtr^�'��z+�Y�����I�ď����\*���:�^��8lԳ�\�XJ�,B�H��"��R��_]]���A�p�����YZ^���A4��+X�'��Y��w��C)[��0f����`�7�l��@�Q�7,NEK��ZE��\%[Z���a��X$�P�TI�HN�0v�UPbٯ� ��r����F`�����y�7'�e��7��\̯~�+�0��4��S	q���p;�>���ET�
��w��l5m7�۔9�ZY&�Pc�rǐ=Z�W��������}����G�B:6|�pvV?���ym���Ij�S<�k�,D*�2T-��@|e2J2+�IȤ#���9N����S#r��#��qC��ଊE�z:�!Ae��[��)%���J$��#��ޑ�IO��fCHa��!x�+����."O��
�ˑ)�������aYjĐ&|�����=��uO�jy�rb���0 �p$777��R��(��!�}����<4�vq|,쀇����L�һ��B	8��
�%w)���࿓���e�7
��/���cc�l�Z�r%o6:R��Mo|�!(T�GS�t��p&��#�pd�O�Gt4ZxhB�{K?9�v9����V��V�P����#�L�"gw�ˇHe�.��b�o���ӗ����ԩ���~�פT�R)��o}f���.���?�����p���&��ЇO�w�"m��d�GCeH�ɲ���
ĕ���ϕIV���X��ѹ'��ҹ������͜�hҤ��&󾾅h ���|Z� �.	����UB�h����W�������%C?���Ԃ��qdxt����� �q��<#�rS^��w�{�`evz
�;aSS��VP*�%]�ڵk�^R��rz��O?�UJjC�Z�+�_Id>��Z��v	)TL�"dAb(���� !h��Lli��FQd2��(V�a ����	���LzdrR��Ç1�=��yJ�����5�}D$� n°� �Ga����B5&�Iܫ���<+?��xJ��Ӑ��Ê��%�9��B0LE���aj�ެ��8��&������J�J��f66����/�ă�����������Շ˧NB��+(Y,T�*8�h��]���e�]�6C�û��|��H"<?a����ٳ�k�����^���p@߯hJ��j�J (1�&�������0 Պ��=��	M�B�f���ݻ������VKZ��7t��~u�ܹq)�m�f��üq��ظk�r��7�jYx"�F�8�棑��t@�������s���G�9t5�������(V��ʢP	��vQ��P���:8�|xp�:|��*l.O�$'���;���?�=Ɠ�f'ۑ���Gx����D�����$���R�~�'�y���G�G�fK�/�����|Z�4�KY#SZ[[���B�R�6��X��^�\l$Ψ�~��8�No ʼ�%h�7�l������
���b��A��ر�c�{���I�#������4xL2<�#�,��0vwcM�`ΉYhjX!��!�`�\�/FF��'pJ�(2�����z뭷h�%9�m�D2}��p��t������{{;�%33.1W��矽�Gӂ;���N��(���ߖ8��F���i�mLCA�UU1
�F �A@L@��A6H���G�~84���RսIk4��'/I�V���td�#��:�d�&b��b¡�I�c37忂����q�/ Ȧ�+��gm��w6�q#3:ϊ���Ƒ�<��u�1qUs����d��ĉx	-qK�*��]�TW_)�/���GǺ4ψC���S�n[�P��f�C� �c:���'{{{��o��ʇ����?	!N��H��u(!]"l�v7�#4���/��lp��R��$�4�R2U�� 5��0j�Ő���?H-ĎN6���+U@�$�8���@rJ	�0G��L���I�㼧#�j(ʁ�9���5u�X�kh<4�:��
1��5NE5f�̿�!{�̵5�K�ah\���{���=�{�t�@�+D�ţ��^�g.��������w���?��?��K�.]�܅��ѵS�P�<����߼yӶaEFg� ���v��ā12������JԩE��{��U�$9�OLMʬ���l'D�He�@���:
��,3y�a�\�>�ML�/.@"��g�	0s3��ͭ\P�:�!�4փ~����9iN���z�(�ݭMxv8&�ց,�j��<����n5p��O��O����P7W��w|qf0譬��nc�7����?16aR���3�h���=�*��:b��*�{7;]�x<7�HC@�j�ʒRn��ЩW=.T�@Չ�LJ;|CU"ɱ��!U8�01�T1\���"�亪�	�� �hb_R4
["7�!Ԟ���g���"l����`��=�s�I���92W���%s��t�Z�q��������?��K�.Qy�NJ3��a��R&�RJ��W!!&���Ӟ�A�� �]�P*��-"Z�����ѓ�S����$`w{���SO�Ӭ�l5�(��0395^*�z]�|z�=.�tjr���8�Dh�*��������I�b�����S��$�{K��ɔ��N�O .��k���w`'�sؼ\!/,R:���@d�����V!#L
�M�g|>�\i�q#��n��#L�M�s��	����fA�Jw���A;��̇�[�h<�H��G��0>
$T&��E� cHT2�dk��9�g�/��?�4�po}5�;RՄ�!��2c��+9WHF��F�f�FN� ��'&C�U��`˪/>�M��͕�%��B��%��u�����3�$��7� i����fN	4���͹;�ϝ>����~w+��W��d:��J:Ӿ�zIK���,X%�6v%��N�7�
%N����d��pאOY5��i��']I{
�<�υ������g��hu;i��AX������A5P��Q��h#�Q0X$�zk�Z�zS'k��2ɶx��������9��<1��S��!�Q��9����n�c�O�kZ�f�$*2YzZx�9Գ\*������XKKKXf|pUԢ?����h,�%�F��<��ۆ�cABdT'��Bk�uM�H���:�nw����<��V��������ܾ}��	��KGB�d<��/�t��B
���vz�r��,�[�8��c��<&��n����os��P��LJ*��;�D�+7���i8p������Ү�l"^���P���\*j��e�k�!�	͗�����s�c�ن����PA�"�)�SZqSF�g��Жh���>������[�n�v��A	��}�̙���gp�fgE>�˩;]�rm��׃MD�Y����Y�d}M���O�H����d+¶_�����[<vu��w$��/�L������x���l���)�����M��qt�k�/���8�G���S(C��`��caD<�;7���l�����Dh�tP?�Ɛ'��8�b ���;xq�t������e#%�P>1��N��J����F��W^y�^�r��G}���OC]H����T|������6C^�)��&,�G�l���/~�h�瞻t�ƍ��RWH�s6�(�1\>��ER�:���"�<���"`�T�R�-`�NWR@V!K�N���@����OX�uݺ��D���Iz����Z�(쳙�)&:���K˧��؂w�+�s�N�Õ���l.�ΐ���}
�\�)��Ci�:�4dl}M*�B�"A����0�8� ;����e��k�~������}p���!�����3�^~��p�r��aG��'s����_V#���)�Ll��Amlnh���Ӯ��7]���71^�������4젺���u���qx��-����{�vF7ք�������)BfY9eQ&�*|.'��y�l��K����,{&ۋ=��?h��m��^s4DHb�a=v��-�0ڝ����.�@r����|��1�V���
�K���J��� ���B���MgK\��ݮ��F(e@(I\IU�j)¹T,�b�4��8����gvA���x�߇woÙZ�B�k���H����7�����4��k��������߿�:![dI��oNp�s�L(^�P�o�m��YGd�*}��-�?�%����L	�v�N9f���RrwӶ�"׮5��ݨK��
Za���1esU�y�2Źߝ��e����fC󄠿�#$Z]Y$���ܔ�L6uz�t�I�ch֋Zu�M��@H�.�~T�|D�Da ZL&�Xx�Mi�0?>�R�";-�h�"֑s�\/}�����j5[2�jh2�'�9�:��a�i�pv�������kxY0��ϟ�����)fzG���`ğ���ˇ�C��F�z���𩝙*YO����H`��������������ַzV��r���kN"=|��x^�s�����W�2��a��i/	�
�S$}�@8,�C/�\>]m����$�%�`�Br�Ճ���%�'��!:8(�Y?�y�P�f���N��"�y��W�v`̣CiU��b�������"r�נ&�\�^p�}��Ɉ�*$gĢ��WH!쭴�7e	|�b�p���z��O���u
�{�������c%�S��ah��ol�O.����s��؁d�P
-<e�]l"`��X�����W�bAs����!tK�g���I��8~���J�
���'�����)Zٞʕ�u�ׄ=!�+��)#��B��%d4�����ư����s��7����(I�NaQ}(6O*dݖ���?�.T�j�?� 8u�R��^Q������R|gWHg�S�H��hR�'qM>����FYl�,mw��J�a!�{�o��~.sٴ�e���:ދf�"��tըФw�Q�h��5��NnA>8TG�YG��������@�XN�8!�[��WP���B�%s�WF�L�����Xx#rqa���:��}5�Ais�E#Ĳש�4GR��Ԑ���6bi��I�^m�>C��74,$Y{9��(҃��Ox��g]�IrN����	���N�!�(Z�����o!�����v���T1n��&�����յ#��{F9��0�u7J�<����o�������#z��7�i����_��' ����i�PGq�𖱄!6��cXXNc��Kv5����y�Q�}qF~�Ǔ��$+�W �dC`�Uؖ(�*M��(xT�2��'�Uj-x�0��2�[2$gr��nu~ib��l���G�����gf��g�K��i�:�wla7��?�)��*1������d��R��W��-Gq�qb��2���ݕ����r���|����q�{��pg�{�zmyv�u'�=�v�G_��ۿQN��{�OL����(~��U;3������n���ڡ��33���{w�^�����UUc1��b��J�]/�#�MesűT6�ˋ�[���߾yP���|u��P�:���D�R��$����'6Μ=W�f��vz>����@�$+c�Q�+�̦\�}/�s���"��W�^�b)�g{��r�sX�۫k��Xq�/8ua��Jϖ�mGJ�!�j9�ܱ�~��j֒�>i�]���N�v���M��a(���ʌ�]h�"3���N�����5�u�L�������v��̉�c)a�~��$I�h6���0%!ѭg<wokӊ#X�o��ʕ__�I˓B�Ӑ��')����imχ��~�U�	���v���iOʃf8��^���9a�wmX�X,��W��dS��i�=�M�~�K�L�T�������%x���!�L�1��ͭN�=^+���1w�驙J��aY�R��j=�؀�D�h�l/?��[n*�͹^���Ԇ�͟>�nI�-���q�u�7"��V{���1�v7�2��L!?1;�����S+�gg�J�Ҹ�' M#��x'Mh�n�i6�d�G�F3�Ns�=7Q��%�u({'_������n�
����{O&��a<�plw�"q�+��0l5����%CB��y]����&7�D� J��>�D[?���KM6�m��B<q�]o�ᨕKe�ZA �T�tG� aă|���m3T�?3tx���8�r_>1�I����ɹ_=x8q���?x��ǿ~���dN~�v5��H�<�A���tf��ʽFCf�gS�~ի2g>��
9�B���$3�l�?�tlzvj{o��۩��L��+9'�&�=!��L����N���Fhi�c��!���5�����Qݫ�ZP��ZMJָ&� ��d���Bԣ����b*����:H-n��}��$���8���iH�ʭ;��ۖ�x���3/�+���*nDtۋp]A(æ�޽OJ��7߅�N�B��0 ��~X������?����%u%������q�0Ŀ���x�x�f���,����;�[�XF<I�[��g,��ӈF�W��z
���ĸ�����%�ܨ�J>$��}�8(�E�X;��c���9I��E�X�d�H��6��l��T)r&BN�#���G�2ׁ} fxz�O���Τ����jd

:�G���/]a��7��x6�I�R� "Y= �xGt�T�'�_ELm�c��l*-9(K��NR����^�H2���"gN$�,\Ĳ�h{u��QdIo;///�_��V����:v��]d�~���r%P1��YZ�� ���
�et�t>�ٞ�ӡ�MS�`��7,�=�������q�B�aRE��2��r�qڇ��v2�x�iOШ�#���ƈ r8f�<��|�q�c��0����}30ꈨn\�����h;�x��o���ADH�֊$�� 0N}��wk2ڸ|�������Ӧ'gخ!e�#���-��T���W�������5���D��ի�g�åK�^_��R���Lhw'��%^w$A��tJ��p�Fb�$�QRA�6�"M�<ge����u<����T�'U�΀ꥠ�|���G�͸1^ؕ�����q>8��8���mooo���$�C��n�C��d�K��	��F�N�Ս"��ޖ��3c��8���E���sr��4$��D��^�:'���j�O{&=,Ť*�$2�v��{���'7��k�:wW�r�������AЄ��Z>u2
�J��L1�o�z�KH��T*\Z*'��XcFqЎ�#d��L�iI&]�� C���{��L6<���촩�����5�]#e�gD��S���\/v���!-N�����T����Jj��@Z�#�9
�,ᯭN/��n �.��X��9��q������^o�j���5u6�f�L��'T�R	sS��z���T�#��:5`@��=�1=r3k	:�����{wm�)OL�iz�9~����֪q(UYx���� #$�����9c�%GK�1ܤ��a�Ed�DQEٶ`����|jj:�k�@Z�BBp?ڝ&B����8DH1A|!\�����'�|"����fØ\�sy�@�/�fW\�vR�Nad;�oS�žL����TR�a��+�P�U	� ��;��ΰcv��*���`�Ӓl:%�t2ްqś�a`�%�"��݃ h��$����n.��J��ȜƤ��)����Q��W�bG|��Wq���������ʪ�]��7���F6;�]?�$^:���5�F��L�TXl>N3�o�e��%,!��������p���(��38܂P���S��t]�p�����[�F�M�Lb�4-Dkss]�y��j��+ ..BV������3����f{�����6��ĒL�^1�7̌����%|%��4�R:/�q��?$�^1$2� �^���qc�e�vƍ����H'u�g�[8Rz�QG��s��s�Ym���%��?��<�+!Ew��a�>���9'��T"}����ڃ�
E���u<Dx\O?������������������R��}b�A�^}�,>%�����ggI#3R���${A��G!���L>'5�b�ג,s�V��
s�m���?�И��(Fmɔ��h7�?����`�B:ڶ���U��H�:��H@�Ш���H6feJ���U�CtP^���\1$���H�/e
щF]2��Ǖ%A��c�j*c��ٶ��I�6���#3��2����0�<�mq��a����<1Q����,�~�E��Bҕ�:B�y�g�
�'��V*�H5�6��ir��{������P�R©� Y��?�x��.�bpjVA�i%875���*��<͏�l����p�?�ĘQn��kRTPtɰ��i�o'�$��Z]Z�r)�q�&�RꕳKt���_�IX=�\��}��;w�<3˒�S�lS��#�+vSg�͞y�&.	k���A��^���*���+(�y��t񡤔6�n�X��û(��E($c�j����+�#�U��#I"�[�;��{�/�����?�я�W�:ȑ�Z`!��@0C�&F��N����;�$o�gE6��<�t5)�]�������/<�s�i�t��C̒ګ<lASW2fװ�Kk_�������ܖT*�j4�c2�%3	ƅP����u��d�ɩ�V���'�\XNgϞW"iG��"�T�[���b7�d�Jy3�f��ƞB&��8��a��h��pQ؁�r�_�K%
������0(ǊB?L8P��ֽ{�������m�{�+�
�lN���=���}���3������;��^�ph�� yLA�V���p����V]�Y�+���^�,��L�����ڝ�x:S(SY�� ̱���%��NJ�]���lv������j����e�0y#!���R`���L�a{�M|u,����4-!�L8p'aq`��Ȅ���!,� M'�tMa�G�㧒�ri�~Xm����:T�#ζk%3������}�4�mwp-X��t�819�	�J#���(��^��P|�ֵ�N���Ca�r�T�$<��aV�C��z���~rK2��8>!ɥ�A=!�Qx��2p�Z��=3�,.���N�ٛ���&w�J�F�@�I�M�� ]�E
t	.;T�m^K�X5 h��͍�ٙ� �J�pog�zp�kc� 	)�KN�Z!�K	BB��S�J���k]��؈�?���xi˱���a��d�~��� �q���ܶ�:��5q3���yż���A�jw�?��#|�ư�o��y��1�gk[�@�SQP�!�,�˖'�m�ݯV�?���]�,�}	ްتZ�|�t��3m��CM�I�G�4۝0F�7���6?���pz~[�����^�X�A�B�d�p_
��i�I��	��8�e'�dc��m+1V*OML>��(r�;{�T��ٓ��������wH�8=A9r
 �>�T��@��lie2�&�&�bm`���{w{�_��@�6��������csՃ=���8��ʉ�1u0=7���ف�QH]�}D7$����/I�J�S��d~y�uJ�T�����|	���<��)'�O�T��е�=KD��E�p���rD]`��mj��6�?n�Fs�����6�޽�����z��݄*��`���� &]�3��0<�v��kk�a	܈����y��Ju_K^�̡+�����lj�R�
�5�
Ш�:y\������D��n8Oļ?��j��?R�r�#�]��c*�o#��v�w��5)��tw��e�q�zC�l��1@~���C��M��3�L�`"��8����)Fx�I��ƾt�Ńʦ�2MD�dRD�e��ŉ��g�&����/���Jje���M�=�b���_B��Mq�?~��cB��Ǳd-%
�g�M�4�C ��?��HyK�t��1�R��7���"�ȧƸB���A��r������p�/�T�4'�c*��22Þ-�b}Z��t��"T����E6�����IE�5�]p=�\8������;x}����hQ6"(�'���M�p�N����x�,�P ۻ{�<?b�5��"i�y��PR؅�Y|v��5���J5���A�l��)^HO[d.]���o���<I
�c;�h#�5���!(	�������³@�(�x�ʱQK����y��]�|6��xY:�hwW���,C�:C�T	!�oָ�$+��n�0�KDW�#����T�J%ڢb��=M�7n@�Ւzuu�QB�g�2��"��|���ݮ�q��	�w�l����°���"qz�s������d��W�-���7��O>����-�2�q���]�<5���J,���v�0<���mJ��li|�
ZJo��$����V��T�#H\���7[u���h��4%�H��8���M�ϴ��g���`ȇ�0Ϟ=�������z'O.u��)�0D�O~9�D,�a�~+5� ���p���7�_���V���X4����,2iϲ��jח�emm�7\�z�i!J1m�֨�ؕ�tx)b@G�A�Fw��V� f���a�>����D�>�0G��6��PB<X2sPI�}��:݉��(Y
�X�?��Y�S�|�_	p?�� �N$d1��y[�m��Jj//[�S�^��L�dR��L��ץ�n�N���zx��r��
_;99��k��,`�h�O?�z,��6�����X
B��$��C��T6������t��X��Ӛe�]�]?T���Η�N�L�d\̉��"�Ц�m�$V�����>�e�Վ�D�XP+h����O�ԅl�C�%��>��l�@9D����W/�D-���Z�����k��H\E�8�BZ� 	�|avv'��z-4��H~Kq�%�ల��$]8î' �8�R b�񹵿��ٓXW?�ѫ׊�t����$6;-���'xx��B~S�>�]R���������������_8��!�"�jx>�T�;�n����~�z8b���P�Kn٣����1�o���X	�q+���pR(�
�!Gf��Ì����{"e[�=q�ݸ�O�.V3�oF�,	�%���0`n��I,��!q���TO'S����&��ȫ�ЉJ{`#nz���i���3�<s�y�����x�F�~еk�:�����$\��s��	�ԩSP�/��2^ l��؜3�@��iћ�裏�"~��
�����O2[�h8� m�E�2lVMp�Źy�������{���_�!���o��>�����Å(t��?"څ�t�j����9%0#T��JZ��n��`"FB���Z���P4�`�q��2�R�$U�2+�~(s��%�E�`� '�	��p#͓��`��=G-�Pйl��fF����^���n�<�66q�)�9�BAZ��JE�I��'�6��1�>d@Rۜ׍E8"�/a�:.�5Gz�A�yM)�Ȕe-ð���%t�z �H_�R�����ʁL��w���\ �C��c�D,���������� �BIj����$����3���E���syu�C��ف���!�1G� ��:$T2���_lI_��g��s�כ������	s�|o�Zcs8.�WF��j����e{�s}��C�K6�3fQ7>"�7�A .<��[��ӛI�t*{<�TR�Y�a�%o�ZL����p�� B
�l�<y1�_
�	nzRR��F��F��r+�C�g�J~�VK����O��������0n���%�YEm!Z�4�4b'�$e�H�[W�������흹�\����*ɦ����/}b�T+2w��.��~�s��yؒ�W����wqm���>�����'�1)B7R^RsY���v6���MC�,;��[��X��z�U�gG�N�Jo_�k���Z1�X����2-�T������$ܤ����C#W/�ɦ�^��oۂ��ַ^���p9K���$ⶲpUm�GqP(L��IX��R������ى�	/��n���+���B3抅��*�����8a�:{�ݫ�Fl;?�����;���
�v]�V��f�&�������������d�V���v,<Iv���l[��؂v�B��3n��­�nuz5i��a��^�셋f`t����Ai�`��&�rh�� �J�K%a�J�p�J�Z������2N�d�8a�����iZ>a��z���L\6��-�;�Oe������"&�¡����V��n���`��ٶ�5ZM?���$_�u���ѓc�XK�VS��h7k����։�JK'O����}������*�r��im���rѭ;��hnll�@�F���/k鴔�.���b&'k��������B�ݪ�
����p_�#[I��eґ!��l2���H��~h����ȫ�(Hq�4ܤ���L�څnw:=����L2���l�$M�ې�Cc:��8��J;N������� ��CJ���P�''�I�͜������xk�$���"�����;Y�8�gӁ��t��;q��o
ʈR�x�����=�2��~2�^��y��v���A�s,8�V���S�H�:�#%nM�8��Q���,�1L�m�ٙ���_s�t��/�_��lcsc�� a;��F���6I�b!X��x�|<Z�N�H��.c|�Ji6[�d�0w������]������m��^�%\8�?��μ��8�}�	� #�%����++�όb��}iN6JD��|����鴋�&�>��i�T(`{^x�ι�1�G�,,Wr�J]D3{��ĉ��,3������;�x�¬�זM~�aI�K�����f�[ȦtPҐ�*WK��[�Ť�6�Z�ˠ�Ν;���w�Հ��>�78;�h��, �W���t���#I���*���۷	���9��'?��0̛�;＃#pl��!.8)84���8�T!d�[sܲ����W�,�q�f8ʉ����c����m-���~"����
FH)�dƸ6mp0 �W&m�24�j7P�	�"�2$OX̔�C}��/�rDB�p���$3�ʸ}i��Pc��W��+�C�\*\~����
��Z܍�1FZ�O�+��{t�8�rԧM�Ѭ�qX�M�S�ݱ�$m -�Mi{��]{��;���z��f�����/�ܔ��W�P�G�:#���O=��n��~l��v��H��'��!:��I1^�t�]��rO��ǙW �� AC�-KJ^#Bjf��������e��ȯT*c� �Z�uMƝ2Lz��ת$c�CF:�^�I+����|$�l��hwq/l�Al���Z��uU!~��e�!���tRz���#�w�W<�2u|5BOq�7o�|��!�r1�+�r�e'�Y|Q�rA��Gc�666 B�U�щ�x ZSh�Qn�ht�6��@:��M�HJa�Ǒ���6q��*��ܽp�����ok�<&�m�[5��YZZ���oJ�VO����,t(�V*-����2�[�n�L�wP�a.X�u�0��NPǄkh�B�4^�s�&d��hvj:���h�B��g�D��	�]�~���0�y��n�0�+����wމ���6[=8��|��j�L�K�j\�xq�T�+�_�i�;s�zpP�V���/�dv�F«�[�32���u<��.��Z�T�(��N'�H;�V�u
Y���I%����9u�ԫ���%m+^��m7���yǕ5۝B���Y������23�Vf�T�c^�``XZB�{�0� ��*�A�ri[ިiE�|�a �	�����p�r�A�$�|A`ܟܽ;�-qo�D��Ims|buXk�x��q)����^��kw򙬛�]��VP�g~:3�������C�k:+
�N:�Ke���� �ᰏM�k5C���y�xzm���dT���<}jamk�Y?Ľ�>}^��?hw%�ˤy*�A	'zzzV��7o�[*c
Ps��!,�@:��v���#��A�=�z鬃�c����.-�����1R����������Re&JLoʩ5���.�?q��z��ǋ����~����'6�L����~XowzX����X��v��ǐ��� �A���Bݟ�*�/��L ��/�i�3</�}iī�!9{B��>X�޿����۷Μ9s�ܹZ�β711&};;�z!R�N���667�s����//1�Ju7���4�z��\|�+��w�kD���pu~v�JZ2�"ᚿ�������w��������3���O��(�`�f����5ΰ�1����P�(�g����C�x� �Νy��7q횧�"�ëq�Ĉ���l�����մ�m��FQ���	%sX�M)b{}Sf��ɔc�� �,.�r>��nJ��n~�ĵ���8�� �E�k�?5�����v�V��,�������A`!����{;`*v�����:�}���1�����Þkk�L�-T�U!�D��݁�drKd)+�c5~�X�2z�%�}��q���d�2�ws.p�*k �xP�y��+W�t�s���+P�J�n�/��~u�Gꀽ�|;$���[p -itu	��)�I�-%�y�`G���38BY����ջ�p�����[GXK�˗�s�BM���gt�����lrJ��?�-E:>?i��W1����@-�xH����!ҝ�o�Eq52^!� 䜼:�`�r��]0�����%�K���L_[�\(S�"Z�.����ʥK�p��/q����(�����i���7>NB$_�S�J�ww$8�z�
��K����Hz�S+{�0���Ly����e4e�G�A�˨I�?��r��L����р6�F�W�e�m�M�
�!�?�c��d��Tp/�@��	k82O�RK��M�ǉ� R�P9I�'���q
����n���f���l��5�a��8���ܝ�
\�=])���_dm���FdSp���� h@V�hM�G0?ǲY�W�Z����_�F�+���0YQ�L-�`h%�l:�������C<���yy
.�Qwۗ����y�l�����7�x�������>Љ�2刔̃^��@�c�̴�j8��,�/��%s�%̐nfvI�ų����1>�5U�Fg��I
�QU�&a�֥E�$-Ћ��e(@�;�5a�U�%ԍ���!�8�$ҩnW2TИ�BQ�j+��P�5<�v��i��5̄N���8�C����vȘe�8~�#�FT$�z��/�_�E�d�vo�ۮ���;���_kߺu��"�ǎ�/,�M^���ef�t������z>�y�G?<����W����~(�6v��=�0+����?96���[�z�9�}&)��ݝ��d�ħ@P���^M��׵رy�����ޏ�� ��K���)B���zP��������]�]ޥ�y���WV�0(=H�f 5U�'�����Y{���o}��Ϟ<y"���j�Fd��[＇����:�1�A�C�#��G}$lk6���OF����'�{X�����H�s�Z�2(������A���D">�J�OF��.j��ￏe ^�Ec#�8<8����N���G'O��n�Du�n�;�j6粥Z�rv쏆�5��{�s6���W�6��9�K�噰�Fј�������E0=9N�V���_�´�Qmǳg/^Z�8b���)�)<��� ���mӉ��.z�T*5��k�Y�8��V�Y]n��{X�y��d����{���+W����nI��^''"�	��p<�����*ΒJ!��O������׍�{;�� v7��0/%L91fIy��\�b�79/�b��bme�M!�Z�A���#A�Fs��2��X�\��7s�K�Yl�\]!�o޼	����+�D,'�$��O�����oQ���˗xs�T�Y�'�Z��/�QȞP���(���xය)cN<n�=s�5gag���$N�);�/��r�m~����A�W��T��������B�+�	��Q��wyk�� >��#�q����e�;�#���'1w�	��t����\��:��~G���;�L�>v�?�$s�<a�K�����8>}:�Բ$F�&)�lB��"9Bz֊,�*Ѽ4�5�lJ[%�\��bl�lyJXc��M�TIW�f�x	�vZ��5w��5��ܗ,����������r���V>y��O����1�-B9m����]=���V�R)e�"FS�P��t�n�R&�*#�����Y��leh2��CP7["�5ql�#<�8�~i�\�0v���>�����ψT�'�~�-Ѝ7�8�Y���oț�\���@��&�u��I���촭=��GY�4���4�&���:19�p!&OO��Pl�-�M�GC+�e���B��Z��.���(���i@)�%�3u����5�v\���ڌ�����r���;Ϳ�d��/��~s�����GOԱ�Q�Ϋiw�pL���v~�+�\��Z��`���S�lĆͭ�M��yv�/}W����֨Sb�^�t(;%v)*�YK�c�R��>8b�q|�J��*:���Gw&؆HRL_X��aχx��uo,��M���k1�"9���/�CFY%�̂8*j\4Y�ߢ�CNLz��G0����h�q��ÿ�_S�
A������EԚ
���M�8xFA��V���d�͜�&͠J��W��~�9�Yx�{��"�l|������!���޹����0`������\쟦o�
�)L��`:T�����'J#W��<p���&�.���֗��R�Z/"*�b<U�֖Yu�J��L��&}ƚ��䀙v(�*��鰫�n/Po��8.Nޛ��3�N&���,7�n߾�d�1Nr�H���!�*��x2<������o�$AB�:��a*F�xmm�t7I��^�x�m�S+޼}���FK�`�uN���t��L�O���8opn�\���/�~��������~F�Z���n��;=:~�@�V��ܔ��d4^^iT�ų�������͇�?:bv�|}u���W�2
m:���*%�_*���A5�y6M�T������c��Q5y/
@5�W�&i�@�4�d186��#��R�G������G�Y���b�Lڰ��l*�1���il�B=YX�H":�#&�F���G��Z�ՃqF ��� F>muX�$�t؟�(
���>eʗ�Z����W�e��z�)���q���SBM�`>c �T�y^[�����l���b}�o�%���`8<G�S��p+��qp<��0�,<X[,0l�_��AB��`(�í<�Q��z�~&�ع�2KK����7�f�9�}��(3�����pjԍ<��#dˠ%"�$�����m#�9.B�r.e�t:9�'i L{>25�	� l�dlL�C,2g\+�$쓏�Afn���oP�PM��C
@%ө��4�1���qaL/r9��>���$�@���t-�卧ѽ���L�����ɐZ�}��*Lb�a1�j�ĵp��w�}�����z��-���x(nƱB���5��|���ͷ��H	�����W��ۧ�t�C������6A@����H���/7y�4.e�c)-fB��K�gGX��X�<e�>�Q��b���&au(�<��b�(ʨ�V`�`H?���.N�oB�b)_(ba0��[sq�tV�9����� 0&�Q�����0��k�)���`r����jwz8W��ݪ\�L/�_�߁�8>m���vuJ�:��"��i�����C?�Aw������WO,���,�3%V���~���2�����������{�ϣ�̗/_�p���:%���kW�2#��b�o>]ci�����������1X�K�7IE5���9Q'K孖��w،Y)��YçZT�ŰB�����o���j\�Kĕ�u�3�@�M,���մ��@A�L���7�O����<o[g��������GP(D�h�k,�<U�d!�����X�DX�����񉸐�'8�&q�;�ү�S�xS�1�~X� ��Y�����<Y��+��a?�?��Ĕ��c�%T_�\0�5E�,�q����5��/`�8����&cmєb#`�IB�f�s�����J\K���E/�:�������,��T/(�j?���)G�[���l����`�d.q0�تt��H���^�����Y���1!H�E�؋x����&w�E'�+e�s6���!�,̲���ĮY���~���G\��?ƣ�T�������G�mm�3[n�kׯHB�+ĂT9�3ßt:4)p�vrS�4ML���e�H�;�hG�Xc������F�L������V�Edw�i��*�s)Z�ʉM�R!5�,-L(\���c�!�5G$Ϟ�/�����SĠ)��K�b@`ɕu$�Z��������G8�R��~�xH�C�����J�F0��n5��j	�f�̆�lu����l�ˍ�Q�^߸z��������ߪ:�aX.,�������+OΚ������ۘ-\�޽{��������q<�Z��B��C��>yWYJ)3�ώ���N��]Y]�����sR���q���&�΄͙U�IǔZ�M��пG�����_~�x����a!~���l��Lɇ6Kv���;o������ʕ+��ʾ<�$���Qe��0�c<S6�gG�?ݮ.עJ=5Xa��(7֙��������g6/-������~o�����dޜo�����+O��r�\4&�T�������U�5��m]�dߙ%V��Ǉ⫁	t.D��g5+���Bn4��g�a�ĉJ�s�eU�>��7���)��i�2�O�ix���KI�]�kZ/��t�^�O��s��f��N#�0w6�䲁u}gW�탇x��2�a.��r�-�f;u�(�?<8�󾾱U(1��o'��TH��������(����������Of��_�q���:�l�G���l�����tc4`W�l:q3m����N����<�j�ܺq��u�}1���0V�밃�>π������9�hTle�n��2�lB��Tt���H��x������n�ז���S�z<����w�$v�^�x��bge�l���:��� �<7�i��{���o���"���9I�:$������hV.�����iT�8a��\*�?��M�/�˒�a;&��O]`?H��w�}�W�[���i���W�^������p��|�տ���~��F}�x�,�Y�i���QA$�����gj��v�%�S�ŋWJ����0�[��˽�����«JW7.��j�;"�_Ej�n�5M��h��YX������\!��5
qu�\�� u��ڢ��c�<���`\������i��_�?X�m}5f�	n���g}f��i
[���dL'^2�Ӹ�:Ű�{�n�ﰲ���E��w�6W*�:�j�D�|#�/�YZ,TVW��I}\��.j�U�Ѹ�O��X2�5��$��u����y��u�3qJF�����l-հ��20"i�<�����+��@ ���!�����}WJU^-f��`D��gU(nH��F���o���.Ό�r�r��������zrʔ3*��T��$���!
}�$s!��(��$OF��` gG���%"�iV&?�,-���O��Șv[6��5�4/_����0�Q(������
��0�϶�K��z�)f���9���k��TJ�2�1�>}��\����E���Sך\�n�쑈l�:W�a�p����Q)��b�l�,�(G#��F�� ��>�	�2,<a��|jy���XQ����ûL�}�����H���[���p��]�Y��c˰�3N��6P��h�es$J�������Sjbe_���v��񱸍�VV1�R�L�p���Q h��Tih��`,�cC�ke#�uk$rF3v�J���<�B�T��ͩ��*e�ʐ���7j�;L�ZB-Z�S�F��K9��G��DD#���5�j��3s�,�qr����~��ׯ�W���1)FN����=VX+���J�C
$��QouU����3*~��O�oeW>���c9��yˎ�;�R�裏���}�駏�=�.C�n�^��_|�~��P�ܚ뇟��u��_^�g8�	̳H�詥�)=3���ygo��:�����M��z��7���Y%,��w�f��V�|�$�3BoL�c�ho��G���]�^���������{����~3�����^�%�HP�=,"�,�N�̝�3��\j,Վ�؂����ny���;���DI�1�����Q_*�Km���Y~�y��>YK�ÎG���A������<|R�7����y�i���3�f�j+�a6LXM�lme����� S��*��G��j�+���KL�.5�˥:��aҶ��d<�x�X�F��/ć�Ǔ���2��dN�f�޼�m7q���FR4�����]Y[����{�|���[׮��߼x���.svrQ^�K��� �^�nO��b�Vo��=׸Ll�R��N�~&�)΋U7��!�M��(q�L&Y����2��`�촇㑘T�%��DwCʿk�a2�52-� ��LF�0�5j����P0Ǫ�����5���>%#a9�QpF��gyj����~�F�K�gF����� ���ݻ;��`k���s|4���0��%��c�����[0�/��� ���dtt8
xr�<�	�w��+(����������f�H[�~�M�\���h��k�,wc��0>9��)pc���Y����݁�k<�~}pt�X�i�hw<D����an$�T��1ǰg۴�nJBפj'5�ό�(I\x:>|w� ���6�����G��ӓl�`Ԗ�~���E�Л��L�u��w��s�B�p�"��n\��x���p���L����w�lJ�_�6�J��Y����6ۅ��o$��P���1�iS⻶��(m������o�{P(��	��B�ܩu\�
�M����_��L�����p�Nf�I�f6�N�`jk�Ic�K��9��f0	:A=7�e�4љAdl.Z]]�?;������-��RP��h��^G����Қ����t6Ľ�5���Ʈ�ί������jY݃X���X���$э7��ڥ�3\��d�s�Ew���ڜ2�������^�띷hȯ�'L�ýų����0y8/�~��ؚ���c(v�6�*8S�F���E��Sv{:�,��Z-�=�c�7M�M���޷o�T%ߘ˄Xٛ[��m���S�X������1�ӣ�êS�H\fJ���/^��]��h�"���%Y���;����VZ��z.[��^Y���~sn5��\��#`$�b��h�ep�,@��'����Ԝ��X��]l�r�j�?v��,S��իW�<��^��S���p=�TVW9�>>(E<�[�:'�5�
�v��K�@���p���c����%6���Y�6�xn�R=��9��~�h�X��uսoX�Dm��A&�wu�2�U˸ǅFB�O�w�,_��<��D�Xz^�!�_���0���;V76�D\��XJ����	�xr����.��)�R��զ�5�.��ǧ3��H�q�{��&���T���S��x��p�
��<N,W�)^*��S��Q�e,��I�G��:�5T���w�)��Z"�\��<8ػs�N�����o��q�c��������_�b�an��k}.���OZgU��ك�x-m]�J�ښ$m+��F����H�Tլ+W���'��3|;n�ѣG9;D��̒���r1+S�-��i�y�Vƥ�X6��h^����4�)���4^�kk����~'V�~x�:}��I���U�z�θ3�,΢��8�k���0&ef��/�Z��&�m�NOO�l�3��Ԏ��b�P)��T�l@R�ϼ��i{��O��e�-����s���ǳ$�ÈF����ؚ7�λF�'��˽Bd���/g
I�������%��������������s�k��;)���ry	~�<͜4I�w�Z?iu��W��n�P�r���ƫk��دJ&̋A���+׮]C�+��� Ǉ����K����5(�ɬ�+�/�m��g3Q;]4�?czل��Lĳ�u|]f���Mc
��ԧ�ԪaZ��s	�K\�bϫt�RvѱN
[���Z��G�q<��<�Wk�8�����n�<�0�Y��V� ޛ�a�I�(�L�vA�j��M�؄�f����xJY�󸷷��?�����Y�;��i�X߃C�b�$?'G�kJfq�T�P���K�Z_Kl���h"�k[:���l�ؙ峣l�4
j˫�-���԰gL�nnb�\��V���I14���#���W{�'��͇��g�� "��%��,�q�4;����3TqR�Qև~�d���pztdum4T*���/=��P9]/���R`n�y�C2������x��}f��K��'_�!j]]'[�`8f|���g����k,|ET(�H��"zls'�I���`-~%?")K���I*�3q܉�h���4�T� ��ZͧO�a�ݸ}�����U�����g�:s�B6���[,��ղD�RR�P�̽�?r�<
�r�T(K�������Wv��b�C'�d��p:��Il��9i������<�\�uT0���9��q/M�j���i��\X�!�u���r�˛$)I�n��V����7���G��6����,#��}�[�o�d>��!6 ~������FӃS/+~�t�%�_��d�J��A��xѥ�I��~_6����{�,E��1�'x:�ϙLV�kyv�������y��6-��s���I��`2�6q�))��)D͒�/���[��Ȑс�]��8>�����_�x��)�׹l���j}��퇃�����W|��Ç��$����.1�b$�P!�"B���[� |��Ȃ�ɂ?J�� �E��]��i��+{_  ��IDAT��e?�E5Ś�2
�1�G��g�!p;��U;��� 6��y�Wd
��8,��%,0�+|d}|�	�6��f��>����E=Wbj�M��*h���6n��ݻ�Hr��p��|�(�� ڨ����zt�'L��&���kC]��{°ay�Ar:](���gJ$�D�vW é��3#L�3��^:�D,FƧ�@����K�-��x��A�8ڋ�޽��'I�Z%��.�{D�pA�R��zS�d�I%"��Q���Ss�hN,�baX���b�&��~��'TH����o����o&�
Vj�L�����#9���+�,z��H֖jk��_�N["S;�v���2��1x-�380n|�F �\C�ò��6Ǵ͒�l���������*����L���{������帏�=dK[,�Wu|�o��Y#��(�$�؞��K�6���ӾO!h�!�h������3���o��ܚ�5�3E챈�PU6��������Ը�,��=�%a������<�+���a���5N[di%��(���/e�g����V�zqi�$�aϸ�a=٣�s_��W���A����ʷ]�5~8M�k=L�����W�����yJr��K�Q#� �kө��:޼ySEγ�Ö����}�uvzvz���t�&�,�|���yj�rq0��2gg��L�L)��*��e�d�TO�H*�!���gX�<%��3w�h��U7�Β7o�I�R_���믾�z�=������,˷���"�OYN=��D:m�M��P�Մ�,��s�24SD���VU%|ly�R� ��괻���	K�ܬٝ��q��̮�4��V9�U�ْ1�Yù�[�����^o`�;?%%����#L6U���{�^�tݱ>�5��%�Bo��V���*�V�a�ޞ�2"�b=� �E�V���$��Sf ��&�\^c̍�3b�PgO�iw�elcc1���ƣ)ߝc�y>$q8v}����6[���$u��#��u�U*U�S�Z���z�/���0B��P���$i���!�BL,�IL�)�E�|>c�ؙa������R*�9qSZr��rυ��?4��5;�sx�JJO��O_��Ϲ��KQ�����y]�F��f��d8�ɁE;5>��M�� ���/1�A�'+��������0�<^�,�Df��>�l�Zc� ���,��̣�a�b�jzoi��M=z�|�=ե�W��_�����ٿ|���s��IZ*O�dzl�"'p~���u!�wt�z�F<�d��h��KF~~F�~:�����s�'6!�����*B�|�u�f��r��^��/�:���Ttdq�],�����K�:�Ʃ91�n�/خ�+r������c�T�`4s*?'!��++L˘Q�Y�>����h �	'�pi�����C:3}i���m�]L��'���_^�b'�}�f����?���_~��矗KD埵�{�w������ϋ�1�<�vG=2rTڋL�p!͓�X�4�D�I���P��� ��o��E''�*̜]$s���?��?���u����믿���d�a�i=�꘎����>��w�75~Gd�p֜�f���ib��0���Ǟ���Q,B�׹c��XVL�&�_o�6N�
S"�=n<�u��gj��0�Rؒ�u�m�I�w����{76��{|ʬ���/��v?4�$�P!��ϨE6���kCj�X�ߑ�1��D�[�QNpȏփ�6�{��s[�Bv��)�ak�Y�7�Ϯ&�'fs��}XC�>S ����аj��EbH(J6{�eRHD��je!�aU컳!�i䋌ϒo�9皌���Ah*�˒�i�E#C���c2ɘ��
-~�P��<n�Pi��9�1�t8�ErR�H�����o����Ej��W/��Yn�h֒&m�4�M���PȉmI5B�G����Tǉ(���B�Q�>�Á�A!�����3�{�N�/_�K�����#�_����\�� � ����?�2�i�SX3ՍK�o���?�w,Z�^\�ֱ�mq������b&J�äJ*r�� �(��9vu�8%���#B�ј[F�m��n��G�����d�|��agg��R�R�p���Yn������u�y��[o=�~�7�H�1�=��O��l�ˉ���47ʸ�N�k�T��
y<[�H�˳���h���],y?��� {�����2�N����wfNf�[W����rc髯��y���r��1EK&=�*e|����x�����1S.�$
�0�<u���(D07Mb��x��x�^3M
LPN^3�<���&����W�.���(K��x�P{:���ð����5>k�`q����GO���`?����6�7=����v����yK	,�Eߩ��b�Y�W N�7`�3�ʛM����&c�����$����E�Tr�VR��$��G�\�����z�������0w����O��G�N���56!i��:�Χ�7o��Vs�"�O�"�f�NN�~�%e;��N�z�p'Xlx�K�-L{.�F��xeZa��#���ቂo�wLM��R^����e٩
'Q���I1��
VޯVk���'��yDhv��m��_�N��}���ѣ��e0�S8�ِ�T���p�xϬ��BC��ҕ+���g�ߚͮmn����T�Ҹ�$�pD#�`z!��n��4q��9&!e<��\���f�Y�b��V;����{�I��
w�/d���/�7�����׸?�c�L�T(f#��{��il�B�ID�#���_�j�L���x6���Uj�m���Qa�����(��w�8	3j��a���a*�G}qLvh���v]p���9�lb���X�7߾��߾������|p|����r����.Vlj\�g���+��{P�X+�����^֖X`~��i�ׁ''qٓ��s�K�+,
dB�۝;��������``><[XDù\wLA�Zm	���;|�S��`��w�����/�Ĝ碰x�Rx'�S�I����Tҫ�؈rl�����$.)B�?=�h�6��9�ص!=ĭ(w���UN
�6�i�H45o['J��=�$��&i�^�@
�3ĳ"��ru�׿����7���w�~�ǁ啸j{{�1 �^�(���t�7H7=���s�k9M�1z	Ă�4��!��P\��$�&���"�A�:���1�< 704���)͌{�\����R#��j3j���gi;����ʆ'CZ���X��V�(>{�I�[���r�[�uM�5��B5��M���M������U���X�W1�_,���r�#y��5�&�VGQ��و��P]е�)+����?6M\�������b~S�YU\�z�	�,�P�p�}�!\f\A�P�lf��R�g�A��>�e
�>����5����ϲ�����.K+k��D&E��f{v�)p9#�����w1D�ɩ_���N�{��	��ܐ�Mz0�%��D���G\u�I�]��9�tƛ����=
Gv�<K���&��lA���>4N��h/d���C����1 ��-l�)��sCTΌ_�����\9�ZU����"�\�N�HTM?���c/�N�)n��YehfU�ز:�1ԓ)c�����z�R�Rm�<e��[�6p5=�����_j���쪠q|��"�,�B>w�ƍV����j4�r6Q�
��\*�Z�i:����$��Pnx6���c��t(�AR�*E�=k����������$�	�8��$�%��{ӄj?��l.Y�L�L�e*p~���Ԫ�o:���Y���oh)|J�)�~��b�a���'�n0���Ǳ5��Ϛǭ��)�5�Z$�^Y�V*��[W�������������o$B0�F}��T���+����&cߙ9��خ��(xg�<��]`Q���1:Rߋݞ�Nr��r�}�{v��^�b1���"�Z߬��O'gG��s�S|F���n޹�~��1U���݃�1݂ׯӖ��s��z\SlU��8�<�`���ꂔ��n��Qhhjn��)!��.=8�u!�z��>�?8;m�
\�^�i�Z;���b^®L��h��.Q��N/�^Y]]�rG���̈́������4y��$�c�r���O�\����Y�����teR'q/��p��
�>��!�����ڧ�U���̂Lb/RmBT����Z�����;7��iKHJ�{A{�q×<=>4�_*�L^&�����[��Ɯ �ga�._&���Is�n�U�*@�8vs��-$b^0���c��
K<��qa��3AhD�c�H�JEx������"� }Ĕoq����2�hxF���a��i����s6<�h��p?�2-����w"?
w8a@��'I&<T&�Q�3�Y�����o�Ȓ�$+t*�>϶��5�`i�խ+F~CA���l���)��ͣL�R����v�����;w�`h._���B�����;� _*Vke�C�utR�ŏl�R�YQ!
&b�)Kc���l>WH��{ɸ��T��t)OP"v���Qy�z����8�z�!��@�u
F��J���\P�V�4G�<����WNx�%�I�vge�ٻ�tjye~E�Z.����W/+�[m�5j���'�)��a�|�W)�l���H5�Vנ���իW�u��@������?��U�Z+�4O.�O�b��?����bÚa���홶�Ώİ@r�fS!#��Q��W�.�s�f,_A�2�Z!g\A��)�Fpl�?��rH�6#fS�_�ҥ�x|pp��~���ΉB���Ǐ�:|�����ʍĥ8O�/��7���j�6�jQ?̆_ ?d.����;�%�sk��E���h�(���w��<Pa��,�sa%�]!�.<�[M����������Ne�a�5�&+����+ą�tՈ����D�~��B���b�"�̎�.�N�I*�
�J8ֵ�U�_Ӫd�UB)#��G�<x�+h���Q�Kt �}B��]�T�ZE\~�C��e�s���wQ8�ٜZ:��[��_���V�Yj�2��S���*Z4jm�-�Zt���-�J]����<mՉmq�g�ZG n����fu��
*ƦF��cI�&2a�����NG�Fj��.�Zs���;�O��K$�c�Y��AH'h6fR���E����>��,,�H���upx��%1k��Pt~Б����n#��O���k ,s>"��7e@6�IW0�3��i/<��.	�j&+!yAB�	ў8��x7|]`�5r�VK��U�I��
]�+,�Jj�c�ezc&���*Ϥ>�j�ڢ��J"y4IQ>��es���ݱ"���f��]�W�;;n��Y���=`7VH\F�R�A`P�b~�C�^�w�9���)�����dYv{��Ak����������'�
.�K$�>�*�II}
G���^��S�f�G�~3?W�t�USI����v�'8��$h4ئpvF�jv��F1��Kz�xg��,M�ձI-�K�N;����󳾼�dJ8s>���K��Z����_w��}݌�D52u\��<��y;�3ƼB�f��D�};?�/�/�;� �%��CWgbҥz�"����
[�X�G�g�y��K�E�� ��#��Q�e}m�����t2��+U|'܎��n���=<"�`�$L����ʤ��(����E��z�ͼ��$�-�_�5˰'����|�j�381��X/�����6��L�8�����a+���s��o��������W^Q�+*/�\?S�d�.��p)�Eٷ��v:l;�z[__�R���(yyuew��ol�D���9u7�������5?��Z�){��S�s��i:|�0O���&��Wch�s��0nc�M��]��.�Q��`ػ�6	��T_�7��sy��\�+/��
�\��Bq��dd
Y�Q�,q�t�����aPʖB�P�`��j��hq��K~��dm���>�(v��?s�j3��,����V�OY�/Gek������UJe<�֕��^l��O()��������S�/�ݟ���@^)Ӫ0�4����C��9����5c�嶚M�g3��e^��:�8�z�4N���	N��Y�Kɀ��s?k�*1��@�e��Pӿ0�V��u�>s�Ы�kl�=\.�Vh��#Q,�ʋX��(�6�Cp��Q��pZO�2\M�X0����JC1��`�V ˕�d�~ޑ����6	ɟ<�=ߺ�.�Dܪ���Ø�x��8�eRcRN�K�o�"�m�޺T.)n���s�M����Z���6mj�g'ǆS�Y0�QI�Ncz[bs&�ߍfz>��3��
z����-��6�'��yz*�p���w���y� mjy3�ٚir5u��i���<�����.�6 �,���2'|m+�P@�#�!eg<�ظ�u�[�a�T�7g�#��U�r�<���xd��
?ga.�ƪZ�8	�"� k2�z����b����mQ��.��ܽ�o����R�C5���-<�T�P++˄ϵ�V1*�����P��Ŷ�U۠+`��%/���ױ�p�⯃��n�I��1��Y�9��HWFğ1b( +:u�´��q5�/{6W0ឋ^�å��4�����N�WZ�ks�;훳�p/ҹ[��ZT�MB<Y8av$É����{{z��K'��E��p�K,tȨ�G�S���q�Ό� alΒflM�7:\
�#ܰ
��z��TV$��d.��W�f#��pFF�z�*nn^��[KVc�P�R�1�fG`�s5�<��z{�r�H�e4��8�9�ys�9qL��d�C&zlABdQE��E&��O��4��Īg�"�N�
��nk���`����2re�E6緎�_=��i��L=��r��{�?�-Y�����Ft���=K4���!9݆�~)>�����zH�p��X���e"
k0���z��BL����y���G��;07~��Z��=?<i���y�~�Jp�'f�m&��XWX^]�
�o��W��fJ"������RʃQ���B������am�R���`^1�b3T�?�q&ޮӞN'��Z�9��7ooo_�~�t�m�������v�����~��8ұh�TC�u�����6�'mS>�ZTT����I��iX g𛘽)Ҕ$j�HXj���t4�;��i2fl����GI�R��j����v�jĆ_[]'0d8�'�Y˼O�_m��
��o��C"�K��a���\�^�j��@*�~�vz�ڠ��7�Er�X���՟x���j�����rH�A&(7��j����q��w� ��2kk̢�i�G08�y�>ΌɄȥL���c�7����� �n[��O��8�x�T	��F�u����@�T��z\Q�� X�vg�c$~j�N�;?3���Ib&x���xXf�3xb�5�GՐd���G;�{h �t�΃�ɇҪ�����}ք����IL	�a��_����4�,��,�+<��u�Zw,���S��a��n��d]��(��=����5��.�A���E2%;d�
\���ݾ!���~�x<�	iî��N���:�����(*�Pm���~|.<2ڐ�X�7jU_����ݡ�f�f��-����au	���m>BO��6��(*c�S����#l��&�^�\^fc�]\iH8��;�}\ȫƩ��sQ��3,&7L�����8��z������9"�Δ����@-��^��[�r���j�ҙ�F h]0��뇞�I3g�t!��x��u_*W�SMiP,�L<Wh��Ɍ>��"�ZRB��Yi��F�8�s�R�R�\<%�ɣ����G�#���S�y�x����~��֍Mu���b�[�-u�����ݮp;
���������#ir(Ӳ����?�I���!d:=u P�k.')`�C����"�S��dHu�7�1��g�d�J��R�@	r��e��d�^���^ÿl�X]��><zr;{��)Y[���w� �L�� ��:>��x}��7B���E98�"�C1�8Zq?�?!�crxx�]S ��7�,l�+d��Bc��t��kR�,�\$�i��n�x�����Mf0K$�x�������:
,?�7Z�;��c�b:���Nbm�%b�U�*e=��˗//�j�px�S�M<�	;	k�N�o�T��D}�����<N�`��R��8��7��<���>;6�D_|��_|�'��3�du��=�T��w$4jn\Y#�Y����*]hJb��k*?,�DEr��?H��+�>tvz,�*��,ҴΚ,���XZ8�q���
~�4nD�9�ju���_~��e&Č��c�������?�Ӳل�,X��=ۤ)sI�7X�-/�zR�䞊'F��P�E�`��M昲�W���#�<�=8��W+�}k�vke�(�ej�'�0L��,Nc��S�y2�����n�ό;g��z!S|��>}Z(/������&	�"�)�P4�\q�]�r-۾��hw����Z����S'��lT�2I��<.����A�31��?�D̓�/�9�cǛ��$����A�X	�b�WϷ���K�P�ve��wb�OݔX�Ѹ'��hl]^��*�bBX�3��`<�Lp�ьNcf�K�T��M9=;db'p���GH~����!������֝�V�$�I���Y!Ȱ~�Ly�ݗ;�ͽB��s|?M�%���u�Q.*�k��%�K+�sp������`��vw$�l�ݥ^����2��P�P����&B� WT�Y�,ド}'�|`�K�+�s�!(-&݊)�%'�q5���y.bK�i��o�r~@5�r1�O��
�`���NO���\�5��;3?��rl=<�B��B�['�N�h�3��{�!��<����[��^Z-�|s4���p������(�4x�Y\�T1/�� �r�ׯ�ԛ=l�N��Ѩ1�Z���-�ٞP��M��̉�B~�����?<!�m�:O�w:�j�!�wW66��u;���R#Ȅ�"�Z���	Ӎ�Kd16K�� �yVa&;��Fl��.���6����'�W�_N��	�5fFy`]y���ָc�1pa��	\ߘ�`�p��!�[��N�4�/���`ʋ���������[a���9#?k�fZG�9^��N	��֗;�n��;>>y����\�|��q��(��b>S��!ظ�.�d�7yVR��[#-~k�<��+.�N����d�0�����捈�n`�!���0B��x�+����Z���Fs�2Y�������:;!U�W(�N�ƥ|؏'~!�ؼ��ŋZ�w���'_�,�\Z>>�]]��҆/��ֆ�02�_N�)ua,�`�f�\/9%�ix�b����d����o���dV�73�?��VW����Q�J�5r:��NPjB���7$#�+���u���Q>~���<Fl}��}|{)��+�L��CoA�:��!<���LBg�$|="�3����c��g��4�{Ǉ�6��� �����z�DRY�#���X������"|��(��?��7�O�/��K���V�����@��|���l�s�����I�ƆAQY���%l<�+���͂��V�7"���XhN���_Q<� �݁���	�(�4��+`1SlM/��;}�_���w�1:�G�~�]��"d��^ok���ՁfA�nq�c��8V]��|�u��T,�Ԃ�X�]�9��>"X�EʂW�OrIk��e�M!a�Wq6$����-�[a#�׏Mo\K��i#V\ߢu�-J`}&d?�l�[O82�ZQT������E#�A
w;H��F������ĸ�K?&,�{��i��4Eg���\ݏ@�B��S�X����������@��x'�>7��(*`�lGc�6�K�O�o.�Q�*7�Ⳃ�,"�iW�9R�؁��(�ǋNY0-?׳3dy,J܎5m`�a�(L�J�DU�b#�m��NtM���=���k��5�Nd��t�gwE�&�XR�)��%R���q�x'lS�����B�(3�J�ڊ	��p������n:Nw�/�e�:�n[��+�R�a�`^�~�g\�3ߕ�u�_����4Y���ϟo�_�ћN�H[4����`��_�P�w��L�>�J����ʟ��c���,J3f��e�:T��'`��[zm��%&�Pc�1�]��d5E��c�|���W+U��ܷ�Z5���G_~�0�mU������*K3C@��j�"�{����<�M�W��Yl�;�|$�J�S�g�~�Mte�j7��e��B(��@��	2f<6>pv-$���j���L����v��G�?������o�i��_gz-!r��F�6.3m2��S��5�f1N�Y:��=��1�k�/:;�Ot�#�S+�Sc���t�þ�{&(�*'����p2��������7^�$�bo2��{�X�8
�<~�����K\��|�̏ � �\�����>2e4��|�C ��w|&�=��2�L'\�x��7��C���3s���~�'��]'�t�n<�-2�yz|�Jť��K����1�`�/�*�jq�����)1l�499# ����"� 
H�C���۞���7����g�9�JL�Ѭ\,m����n��Z�&Ҟ˗�J��w�y�ٳg͓����D�C�sEuފa�x�X��a�n2��ΥK���ƣa��$��n�^���(��KE�����=�y�J5��0��%����]��u@�@�\.�`�?_0�&��LdVJLY�����*NS���1��:���b�T�T���U2�W���s�M���B�g4��a4�h���3��l=Ig�d#����8��'��JD׮]�	S� �Z��P�|#���� ���_YYj6ۺm	���-9O��H�"�(���$!�K�B�p����������?���W�>zz�gWJU	�!��k8��sඩbT��K	%��dy�e�-P3��~���6���#��z'�7?��_�S��D����d)�)WQ��,Qj�6ٟ�0�X�8�K��{��F�K�9��(Y��,w$Z�V{�FY��k��.�~��K[7骏�8�q-x�f�驐��q��:$�'��MucJ��L;Q*�� :�*0�A���/�1(�Hшؚ���spdϺ��3
K3���m�ϻw�`I���W�����?�t+=ǥ`bTt��N::�QV���<��7���!J��E_���������v�.��E�OL�m>����eM$���߼y���aW\޺��S#D�U�-���&g�rb4��,��="�t��=t��M�smi>�����g��JIµJ�x2U)��W���n�;w��(�Q���o�F{<UM�ZL��䓩��X|���[N�N��~G��ؔ1;;0;�}��9����i�ǤrB4@��9+�[�����7r�3���HOE�>+M'����I�L�\�x�mȄa��WYQ�jE8'��&�$H�x,���LHC2gd?�έ�4�z��(G1��S�u������ݻw��	|a����pj�'�={ųب_Y��h��}� ��6���^-q4���F�E�F|�~X5]
��4Ül����-��q!b�_�O��0��0�
������sN�ˊ�9^�2���j�Q�5/�<9ly;.#�b�|A�⇁�""�He���.�/>�#vJ�e�wH�+W(�4����	����v�\b��RRޏ��a�	�»��*�1<�Ѽ�.���J���Tr��q��0��$�(B��Ya�VW&c�jqJ��Z�В�h<���^f����f�
�=��2�O['ر�n��%�S�7p"v^�0��#��|4a����Sšؖ�g���,�4X��x:��ٲ�&i&��?3�r�ecx
p�\o��W{��1�L�AM�r�Vv���:��&�_��O�1b%u:-������/�1)?�I�D�\�B TQ8E�e 9N��آB^���@�,.X��}��AI�њ��ڨ��,$~Ⱦk���<�\_�泘��/pxn�ֽ��J����R�o2�}N��.������=:<�?{R��f����Y�Ş�lA0��xST|�>G��v�L'�$�XO� C�؅+nj`���\I�|��øR��v�����7$�i�� �������� �y�K�V�g����$}��ʕ*�X.q��y�Zy<�^|b��l(�lx�����"��&!�W�\'��Ig����X@����� x�;a�T�ų� ��?�_�1b�1!:Ilj �=��� ):$8�(4b�$�x��.F���7�u�N�ݻ���}�t�p��m�yJ+vrr6O��>��]���˗o���������˗_��пiq�P��`�ΓB.O'ƶ�,e�a����9�K�U���1b/Uy�I��1�Hz�����V����^��(����dJ�e���7`'Av��d�c�������QF�A���>;��H�K����,�ʔ�Wת�ǔ���Jn���nu��f40V����gR��`�0G9s�����_�����/���ճ��Ӱ������/?���?�]������7/��.��K��F�],�_�Ѧ���jB.-գ����<{]R��-Wq|Ji7�cT�W�4��̥����0��k�㝂�./׬s>o}-����l(��ʐ]Áb@�馦�L��'����|�������-�C��`{6�$@�I���c"��4����$/���=j��|��x�Ku�:t71]�-�N'�,W�fl���ļ���Sc��n̪U�"�K����3�BF+c��`��B�iOj&�������Om�ĥH�q'&�;3M�Z���cCH�2FurL�%������?�[\'�g�J�DDӄ�B>�������(���!`#�v�̒�Y���4��gR��J;'2�C���-�(���N}j���D\+��Φc���΂C��M���8a"�fd ���d=���xL�EG���O�D���8G8r��8�D��Zː�\R�`;W���R.P:�L��YZ^� ��3�G�P�͘�$c���F��\D�����-��hv`X�B�s�?(��`װ�
��G�?���X�Cl���$���S>�}l�]����e!���\9L�6���*%8��� �D��N�h?r���J��E��8Bȑ��&�/��/^m���Ep��cC����{,��������h��C��(H(j4�`b�ީl���tl8� ���Y�ͱ���(�0��@+�o���~����Ê%�#i}`�CX�٘keql8?��'?�����TCr8��z,�� �6�v�z�N�,8��hl��E_��d4TI�B��U���9�ق�`B�����q�9g0sΛ�R1}u;��O�b�i/�q�Z-��g�'MrKQ*$Bt��w߲ܔ+�6����:�Rg6"����<��������c��z�+]�z�u���\oXaf�,��t��\�aN
_3��A�t�0y����w>��듓��~�W�n��o�;8:��@������7�J������/�˷��#��ц�M �h��sf���v&�U1�\J���B�͎hy] tV����+��m�(o����ĝ����Lt���J�N�l4�W+��_~���G{���V�bC^�}����h�"cs���Oa�6o^S���~�Ru��s����T�N��91��*�R�Qp*�o#]Z�(n��e��v;��L@3��cj¥�A��p3��jօ��;�ܹ��c���es7���� ��l]��tV2�,t��lwQ�%�����ق��X=�Æ58�u�r��n�������������(�70�qB+°�~�\y��F�I|��چ��((�=wh4쥚u�w� ������q��z[w�����gե��S�;��[��B���Ϸ_���f�?�`r'�����ׄ�3e�5�7cJQS|i�����`�K���ɾH*^4[�1����p�:>I��А�xOb�&i�QrNm~�Q�x�I�r���V�XA`�"`�bX�"�0s(�~��'�v�*O�wVQ����V;$�R�q�<#ҤH��x�mBx��W��؋pS�(9�8�<;բL��-�F�aw��V�����sN�m|��������NN���"�ܾw������Q��eM5�IFI�$�',�Ii�šf�x����t4������v��Q�9,���,vpx���KE
���ו4@�Pƌ��1��Nu���#���R$	6���tK���ӳc�ig1���c8wy�}A��R�ĺE��)�T���X"�u�K=��G��/�	1����~1�}�6���矷[�Jږf�]����Ч?�HJ����ihbD"���b���Ĕ<��ţ���h�A0p�Y>2�T�҈X�B(o.������&"����^ �y�Q����eU+��jY6:O������Ċ���2̢K�~��CXOu)�x�J�w���˰��=��:�i��a�� ���Ƙ\���L_d�z)HR�� v&����^�.�6��3�m���dLY�f��N]�g�|��g�r,��~��OH����ի��5�r�s�Z��U-�e8�"���!�$e�J����3
�':�4_t]��R�2b8��b/V����6eҩRc܌�4�5�BQ��+q�΄����V���X��cx"��&	���#�ge]�Z�j[� �'�.�E4��a�(2����|����+�7���BU\���^��`�֕���t�w��m-����'=�jo<R[�kM��!d>�Db0�9\��b�T��b2MJ�\����:�vu}C*�
/..�Z�oј�����c9dH ���/kZ���y�g�6��^ϓǍ�Q�>�-7���f�Q؊ߤ�N�Mm���K��Y����]|�.���O�3�U��g|�q.b��T�jq�'���qb*�.�O1��1x[��q<(4	;��*1+x:��XiOqK�_�.|����t\l~1 ��{�H���X�_�o�B��8�2�K^��8����,����/"��R5�����L�R�+��\�t���!.�
�/������Ǹ�;w߾z�곧�''�	�S]�~mss��o���v��챩"q~�������P9X� 3%N�|�¨�wF���xvtt��[o_�r���~.
?����F݉gyn�<m����T�C8A�:��c`W��UCVdM��V	���G�����u䨩Ji
����}Vu��b�Е�G0�Q�~��^��pl��LlN��R���ex8�1wW�\��?���*���vI@m��;�tS�¼�$�$ω}����B����)8FtJk�^-���� >�J�،��l�뷮1�/d3Q�,���xA�?�ن�����3?�)a���g�ԅ9�V�涎.�A���%�ׯw��0���*o߿��y��9���B�#����{�q�6>�������ad�;�K,������q����p��O�2���p���܍�2�ib�������>ª�x@��x�[�Ջ�<�7���y��
�Lj�v�Po^�s0�	T*U�e�����a��F��$IT!�,)A�*+<���s9��j7x�U[�Ŗ;E��Ø~�/WT�3�ۭΥ�4g�'�ZndJ%�xZ$j�plĂ��*��ǧ�V�m�'TƜ����[�7CsR�}{�~�;P�^����%�B��������⯽� ����s�R�����H�:���EX��#R�O��qi� ���<G�^X�A��yb���х�1��;n<�sl=/���f��եR���a�i����_�6��~�˯�oĩ%�}*N�6�ft~x��Éj�������|dTDh�h�<��,,K�0T���?�����l�|Y�H�Q��П|#�y�&fGP����l����J#�`�#Jĥ���;�`�o���Q\%�$�V6a�@���Ν;�}��g4R�n�� �����B�uo����{�=|���įNZ��b��	��d�'+U����؈w�}��_|!�mo��3¶�<���L !��09��� �r 7�:�kN�@�9�Rj ��3UJu��a��('��X�1�E��\��	��+��ϕ�סa쇿��o�O��߼���d�%�lx�ޔc�ER�(NKb���f�b��nX����b��F�U��(�*���J���{�=/��3��bT�@eeF�x���w�����>�h��|��ţo������c!���b���+�5Y��G��H'��l^�e#U^ qY���/���Y&Ӣ9��1�F�N�$0�m�Q@�^�Nll�:�&A	be/�pC��tP�3��eϪ��zO�8�s�D�ys����+�1	��"U讨5ķ��p�Z�"X ^/�������#7Xۗ�_i����c�^ru����5v8�����(l8lUB3B�qRTv�����Z�:>��4K�	_��޼�����fX�M&H���?Y����eYQ�|kHѮ�VE)�SW�:�^aY���k<�����8���沨�弭�>�c�Q�Q\?�aga��c5��w�ɠ;s+h;ʜh��.M�����p�x�l�D��Ō���z�!)����N5�e+d�Zz����x4��_�擱��@@T}����t7�˳�7���o�&�4wcw<7�rm����d���j��U5rB��|����y}�� lL��K�Q�E���GD�gg'�?*!Z3�-��h\�G?�u�ll�Y���K�P	3��
b1��=�RP�1�z��A��;{����M�V�9���h��X�)9��R9�ߞmlm.�ew<�XT�58�ϟ1�k�[��s�&Ӌ���?�}��_��+차Nl�}�O��_�aU#>�n FB�l�!y������Q�{�n޿���}�b�eo�.f��{_��+Ro�Z�X�f�^��m]D�KaZ�lP*�3�,.Y�QF� ���b���6yJ�V���x�o�4���^߉���&|y2O4���0�wo��{�|;���o����4H����l�:�h���2?3���Rs�M,D�����&\3��]�^��D�,usW��L �j������Ώ>|7�lvE	���&� Юp��8S:�Û,�Jd��x����d�C�Dt���U©�̬}�.��vA�*�礌���$��i�u��}�|ws��^������!(�e2�K�z	�Y,B,��u���t�"(�^�?��b��1��LӔO�/:�U�-�W�=��FN[8�-�3/&K6L����f���.�q{��z����f%�8�*,����g����T�:�0���沛�p�
�k��LOY�àp��5jх��k���oӧ�d����/XO*�L|��s5f���m����7���v�M��̓C����Ç��T���$^(k��n�ql������Ƌ
3 �y�M_*aF=���|:���5|��ݝ��QR��O��M_T��- d�!�pg���	�/�
���ד+�O�q��������l��9yZ�Ae��Á̆^�w[���V4�J�[���C�,�>k���9�El�&I&�h��nwN�+lS���bG�𒑖�M�!'-J�=�BRy��7�((Ș�,�gY
r�ttt��?9��}��x���T:h9e�����%�I\���R�10j�h���8�U��i������]�"��m��$��T$�C��;?��"��!����~�<��"w��aW�-�cxp��p��6pa��6O��Yڷ)�"�Q ;�EPVd�F�Z��Ք$
�&���f}�"� q�&Z��YDz��F]h�F�ew��']*�Z-���Y�LE*��̾З�oP�rn�轠��
�^jI!6����/�%<��7�m����ڶ�t�L����b��?�B��`�w�C�>>~��W_!�{�.n�\c����<��&\jb����I�����ٔ�������#	��63[5��W���K"�7n�6��x��׫�@js5�W�</
�8�ђ�ɹQ�{~@R�8S$Av��7���K��&���y��j�x���i)�Ty"��^ǣi���8�8�2�8^I��c+�R�A���牛Z��`5-F�����@NΛ-)��;{
p�X6�y�b;ɓv�<ǎ����Z^SRTX�ੴ���W5�y
��Ⱥi_7E0zF�;�wU-[#�S��j���e#anCp׭W6����{�>�W��_Mc_��	-�[�t����*`)c8!�*���5����LE)�`�Q4��"��ŭ��b��J��Ѫ�,`���o��t9��	83�7H2���"��â�{��F����g�>�q�����������[��������wv��uN�朵	�fŐT�P�p�dTx4�|�jgw���ؿgϞ������'xϰ=��pԉ��3���g �|�uo�w�p�94�|<��>�{�����EF�岍��!YZq¤���H�=5�I����L�9#�DX�x����t2���!p�do`�j���X'"~�i�Z#�5�p����-W��qL���4���&��iT��f�d0�fs�A\��?��Av'��o~Y���]v#2�KvLAG�yf<�����́6\f�u���D�y�մ���с��rOD�Pr.��|9whv����ۻ�����?�Ih4;�n��S�&ӛ��c$z�f8oolsĂy�:'��gg����xv]Mш��	"U:	҃����z"Wr����`:Kr�w�w#d���*�{ap�c�s�M^4�AV����R^���`/�l��S/�D�ٔ��$��zq����v��T���]]]�+��F�7�c�!�,�g��|<�.�&Ď�q}�ls0A�d�ړ���{X�z�]&���U�U���岳���@}$�u���u)����l)�r��
�E��5k@���n7�J ��b}�>�1�g-.��f࿳�w=89�����W�^���88l��y<�;�Vs>��2C����<e�o3xIs3m�S,S/�P[���[
9�p\E�0(����N)^K6�*^�4	轀3bKa�'V.��#,�"r�$�p��R3��Ce�m{�w6wO�4T�X�$����tbM���^RS�;dOVt���\À�ø�<U�Ͳ��å@��j�,�C����H�Zgȡ���Q��'8o�Cܹ�.��dn�2Z3s��8b������Y���~m�	�|���������h�E�ƴIrqq�-/�ŰH8��ق�u�`c�l� g�Q�ʪt>���������/8�{�������v��[4ǲ�D�Lp�q�����^?����~2��㏠t���>�Ej^62��z�5O׆;���RxR?,�p�#+�8���d�pei�,�E�f#{u�KC�Z�A�
�L���S0����u2t�o�Q�~���wo����ok�E�R��RȢ�oΙ�
�cf�ݚHQ���	Z7�z<�1���p`M��#j/ǠDFQ7e*�ʌ�
�R, �|�	}"Y^���sqhv�t¥��59��S����!E �k�{�S�Q)ɫ�'�Z�V��K.�}�^EN�(v�Yf��w�`���Ę��?��i*4�:錌`$"�u�3l����Ep�8t��t���/!�O�
j�R]J[�co���H���7m 7o�y�U��E��O*4*@TFh8��|��gd,M硿��g��}G�B��_�=^�'Η�7E��G}Ԯ�H8a���m]]D׫�>��%�����5�i(�c���]*U�+�厇t`����8��L����ώ�n"4[�81e8X_!4i�,�\�s�ĈMɅ�DC���������C8�3�����l̸2ް�$Ǜ��u-:d8R{����uń�u:lrL��o��`3���L��M����!���#��X�Q�9�4�cW�h�m�S�F�p���������,�tZO�~�\αI�N����rg{����R~��gt��3,��|�����4b�i�')�%+8Q&����OPX����2�0��Ɠ���}��Ij����e�g?�tٗ_~y�ƍ���q�
�������/T�^�L���6�q�y��՛������@���2&�z4��/�����pi� ^�&����ͤ��r52վl(��, g���[b/�37u��0�Uoċ�؂q<4T����;7n`�O�Ύ޼�lsB}ș�1� 1��Y<S
+�2����ǀ�9=�P�i��*O���PU?���◳�bh�KM����˫����z�yy��V��|F_92x���<t���p��s�LK~�n����9����r�e���G}bs1�&x�G�� �^��c�����
|F��Z����-�]�K_��2���%[d��K�bl�D\�H�rE#:h����$��#��<�-��M�\���6�",O����W�]�՞?#��፛8L�)��W����Bl��9��%�m:<��b���r��	��5�O�z,}˺[V���")T�
�a�6^�c��}���D�E�aG���V	����yT6�e�����֭}��hKp��x�6�G��&E�op�'~.�
��C���Uk�2�Q�=�z�`$�B6���=#�QWin�-�b �	�0��j"lm��J-)/��jX*�	�p:!h�٬ï8�썧�n��{��?���Db���?��O���J&w�
���U[�GQ|j��ʨ\��:$���˨��2*a+2���L�/�DE�f����:�i&���6=妸�Vt��f�~O��6�i�u�U���F��ߜp�٠����]Ꮰ#�����$8ܽ�'�S58��k��9e1�Hg���e0���{��CL�i�*#����������ûw)j�֧�~
����l����y͉˭-���Jq�#�W)���	}d6c��jd���D���6Y���$�r�L X�0�
~7N2��܂]A{��l���'GP.��7өR4��n�`3+k�q

�i\�_'�q{\̓|U�L8����]hm\�|�u4YΕ��`��'USK_�C��Vy���b �N��W�^Ag����f���1¢��2!��-����tm���O�l�-M$@�+���#T֛�����ǅ�C�J}bTe㞍,������[�����C�)����-e!��^�ȽS��|q%��(~��"
<p�g��련Hn��ٕ2R剕�rc{�Y[Fjw�/!��Zj����q����Z�����e��A�r]G�8<��O�a�T�̶���Z��c��M	�
=�uvC5����i�%�,���_��	��,���|B�R�kz-�� 0U �IL�$�Do��+f��tI��{冮9uf%��I�����Ճ�I�U�W�t`��}!����)��C���M��%i���j��/*O��QNB28$�<n�xdK��P$y�1i�YŔ�bt��ٷ�E*�1�xD�;d SՄ������g��&E���;g���O���F��w��z���Φ6`����s8Y�n݌���o~~~fe%�\�����|:䰸�]XMu8����ϝ�ѷO��Ç#*'qj��p�8���2��F3p���^e~%�6ƣY��;��|>�T����?,�jt>;(��K�J	YUOrV̧
��j�c��eV���P!��$�mmlt�d�#x�mT[ݭٸ���|�	H$�0#���mwdEpH��FC�T�5�7��#�Z%[��:��8����F�"��[�*�;G�ǽ� �E��h6��V
�.鱼�x��q��Y�xy�����k�@��&��`�&Q�I<�h8�A[Dt;:A������ƌU���Yy�E�/o��ݽ1|<�yL����1�[�O_��I�9���n�Y�v9ڨA2���3��k�f�c �ٝ:�2Q��>i��?؅��+��,��?m���Z�	�nwc6�]��g�y�׆������'��u��b�#8tQ��ҩ�k����jR&s�='��q(�����;��Ō\U����Q���H���DaYX�n��Y���R�gV�������A�Zk�7$1s�Vo��ݓ�a�-��߿��j��=���řw�_��f�T�?��E���T�\/��0��Q� EI@~�R�Q���Y�f�����
3npm��V��Qb���B��E
Y_D=a�Gg�%�$g�����V�m��6^,��f����h<]��Oo܂�e�)�dʸ��{�p�Q���9_��3"��Z��"�+I��m"^#Z
�M�������\�mo{
Pbs_��m��E�D�z��i	��R���Kh�e�lU� k����h�*nT]����f���9럗���Epz�N��|����J)�<�8P�k���|�����23ЈS7�N��̙���ɔ#*zW����'�y�g��A��n���O�d����h�.h&����=/����Rgk� ��X�z�)�f��j������z�Tn�H�uú�~Z��\6�
Y�_�aW��j�SC�8j����O�^ݶ��ç�<y"zL�5��N������w}��|F���Z�/��f���qN-�M'��Ç!v8-��~��	��-cr��c���W,��M5�dD�Ԑ����
�栤ҺR�r%T0W���HGIA�ƪk~��)�ŕ�qV��6-�����Ń`; ^B��^p"7� �c�X}&6�3��>�e��l��H}Rr��1}a�ݲU%6�-,���rꖔ��u^�x�&3�g���Y�O�l�3������&��\r=�>(�)�<nL�N�NEx�jE�.�>&���W���6�"���*���:?��hp�'!�����TI%%��2*���'W;1d�Q�-O�����o�=*�׫-Q�#���ȯ�?�\Ok�� �����&uK�V�Q�o���G�+����n(Ba�rW|���2�[��zf����|C1
������j�@���n��eK��U/�/*���X�Y\?�X��,i��7�[���L�q���Q�Q���x'Y�,)(�4��V�^�e����ށ5U��TJ��n\�}]�p�OS�.��,4�M��i6��i�fe�<4#�=p`�T0��<s`IgS��ݑ$i�����f�%�q�4v�����gu��t�6x���F�K*��L�=1t�hH3�j&u�Xd9a�b2�H���U�|�7���g@c&񃡀�;�5z_\�m��;-��t����E�FQ�gx���rɺ����]F�)�Wp0]kƦL$FXƉf�[r�{�r�Ƿ!w�a�����"�ys|T)�޻s�������b��l>�2K������fu���3���1���te�����
z!������������� �Jt(�ɜ�:����T�WD��b�����}3��68q3xp��S��"Ď���=\�Qk4����c�W[�;�,�&�����2c|j/��7�����q`�W;A1�;�8�!���'�ydaƗ�Q��^����m����s��ME\f�]�|�,�w�{Y��٪�t<~��-�(���ܬTfmc��Fc|����kx��l^6c.ӫL�t:>=}s��@Aj�xn$zʿI`H��n�ɥ��&o�zu�S*��eOS�LN޽sZ���	���@���N8��jE�h�X}�+~&��8�j��i��'��3��
Ή�pyn),���Y)hߜ��P:�e%�܃{-�^�ͫZ������U�/Bdϼ(&���S�����P��>7�[�vwE[hI>Z���	�6�/f381�R�W���͍V�fgg��D���"9�zҘt���QT;��B��q�׆J-�[[�_��$̉�8,Y��N�d����R�l�l�+r�4��?X��xJ��R)b`3�x����N�zjx���c�k:1��}��%�����t��h<�����(5���l6�#��Al<`�`�W4jk{O~ttD��U����\��%�8*�q��l�������1@����qB|)����Ҳ��̕X����4�O��:�;I\
�������Q=F�|"͝oT��[�ݏ�:5�U
�M�%�G���Z�E�gK�Lֻ���m��mB�67���4�Ⱥ�K5g��q�gq�_pS�1R;-�L/ �������A��,���/��ƍ7���kժ$(��a߬(E�P�&�b�����*��l�J���Hn*I�:t���SK�_`�b&E��P�n�Ϧ*3X�8=�D���w��`'ư�
�zM�13���P+��A������O���f���!NH�$�������2O�>�b
��ⶳ§������-o�T����vL�Q-Ɖ��q�|�	vyؿ�u�{�w޹s���x�f���N���5������Ù���K3S=�T�̳A��lw�fč�j�Y��]Qa[6�깦�]�2C���$���n�+r
��5�RZ�Dp���y��(iS)�^������1-.�l:�nL�U,��*Z֥�[�*��Z���p��85��؜nwŭ��̃c�p��kH�jW��%��򌜶����Șв�ۃ���Xa����x��>��t�Bfߍ쭸��s��T�ǚ�bs`�ɉ�G/���इ��3��T��}'I�ؚA��g�`����KT58�Ϊ�'�Zu@xF��D���sZ�:��4�Id�.��6'��<S��+�o�,��0ms�z�2�Yu��#B�6k�V��8�.R����W�XM"���
��y�\l��k�_��A��ڭ�P!$\(��aM*v�l0���(�u�b>�<� � ?cȢ�&):��+n�9��_��M뒹"F�I`�Jcƕ��W�2�A?a:a��(�7w���^/���|��۱ �ɩFq�9T�̀��r�E)��u ��8N�cɌD�{�{!��2�eF6p�KL�57s��f�%y���#���Bn�����f]������܍�#�U���ٕX�0��E�'����UA2Y�A��� ���j�N�iN�f�	�3[��"`��ٶ9Q��=x?��=)�������$�ݺ���<��H�g�ús����!q����,M�3�=���z��3pjg�-`ooj��]r*I�"pa�&�L#ׯ����(]��?���D\�Ǐ���	5�<�\�NsQQ������Ա#��:�K�TÅ-�VY�Bw;+�2k�������6w8UxF(t�~{��2�)Y�J�[�ԩ��$�W�K����3�̗��(�������iq���U����R�C�Vj�L����\.�I��d�v��,��0t0 ��4�'=ion�6���y`x��@i�\�!��ןs(��q�2�xR�V�3q��rUp�Zːo�37o��:#��M#�&���C��i�=z��1��ܸq���z�2�gixy�֬�ɲT	�z4�,b �Ng;߽��+����xJ%���ij^���H�7�7D��������޵\�üx+ �[ ܪ���}�z�@!RX}!e�o߾�����E2.�i�iÄ~S�8Zs{�P�����fc~#w��RnA�U|����G�Z�Lc���M�"� +����8Zȴ�� �Vm�+76H;hY)�!����;�2X��#��{�7{c��v�lt��X(��(��;�����C#]����2dȍ@�{X��屩HݤK4e,A����p:�8|��7oT;��h~��f�Nr��2a��F�+�D���K
���
_͟�`ȹu�.��>y���wc��[�IV��o��;lo���^UCj.���+���q��J���s�>����Gjk��*��̷�~�Ku;],�����@�]e�����&޺u�4$�S�	�_\dv���ޠ�<G��)�B�h�C��g�Z���}fP���d�T�}��9�#�#d_��n)V
�V���I�K���Nq�Sq<͛Q���5�U��S���x��P�%���z�%����d�4)���[3��x�S�X�pC�aW�&A
��Vߘ��<��{�Qp�X�o-b�>V�a90�b����Eא�u*��p|�v[[	.�2UK�Rd���� M6Շ��n�O�Z�P>�%T� >7�=�b���.j�}�S�R����Ν���'�L�JQ�!6�޽{�v��ߎ,�h�H�wqy��6�J�����/�v�lVm�C�3��ف��\��b��:v[�WY`�k7'0�� �r����O���X�-Ǧ6	GAp�(�V���w�7_�z��4z5�M��1��!'d�[u�������1��:E��u�dɕ����Dl�N�����ӓ]�n���8���0\�e������YjQpL&p�U�(͛��+,϶�X�J�ls��d+2�E����Sv�=����t�|FO��6���*\&���S�%3B�[[��Re8���s~�f�徵�a]���r�cxp�wu�;::��-��u���Gb��Ն��X�sj��K*9d��hZzwa���`��<��r�)�����9p��*Vf�����d�>Xdb�Eփ|K�r�
��~�O�(p�\���W��vX���
r�*=_��'�ot~EMGa�I���|��aET�/�ǎ�>A�T��J�f��lQ�M�'��/��@�3��<y�Srȭ5��|G4���ʝ*ˌG��^1>��?�9O|�E|]�U.�yr�Z����dE��u�m�j U{Z��Q�͵�e� 7.��S��Ŝ$��t��a�w�`e���QہҌ1+ϡl�ڞ��Bg��7O�̝��n�T�{l)m�K��9|~kg�?������U���T=��%�)>��B���OYO���++��CKl3�r<�C��6_-m���Z|&�����y��8 �
�̧�o�,i5j�ۘ:�v�T���]n�@���=�u�fQe�����,wڸ?����Ű��i�Md�Vm(m-��!U�!~��/_�9!����P���8�K-Z���5�w���Eh
�ɥ۸�^�b$1��]$�W��_���x�Y3*k��H0*�[����E�g��5qu5��q}EC��Ђ�Ȏ
[�����:��{Q�A�vW���bj�[X_��f.�ĭ���./D]l�{�. &;��5�[��B�ϫ��j�R`��V�β�kF�[ s���C$xҳ�+Y5�<Y�ï�C@xK<���i.�̓۸[!5zdC��r����Ǜq�_~�%n�ٳg*xꚊ�R��V��=�i��HhuTLI�Z�"�L.�[MY��lʱE���#!N ����[�h6�I#-��6�����Ϊĥj������G���^n���rU��5�i{�ř�g�x'DfC�Ҫ%lT���X�VR��f�Wb\W��Dsb�ˬ���4�w����,ٰ!=KH�I�����j =c��9�h�p2s�Nn��J����c��B`ć!�њ�+�55ꋌ@Z%$5�NyHs�<��3���d�,��W#%��N�&?��v<^�}�����L#�� a�û6dp>_����c��b_TB��ݰ�,G��[K%��J��c����2&��b�s6�/oƳq����t:_WG��h(�o~�Kz{��喈����>�y2��2j)�����	� �d�CY�`?�RX�ߕ��۬�#���[P�X���g�Q�g����H|������,����O�{o�$ޣ~A`�k����vM�Η^������8�{�f}s���Ѯ��4J�q�^;8�?��ɼ�g�,�S�� ���؉%���,a�ax�\�L岠���	K����چ��T"�+������3�Ćh��6���ܵ�F��7�O�Y{����k,D��j�2�Y���KU>����E�zE}Ξo�ڐهŜ;3��lo$��c�����F��p��ti��l]xT�KE��>�ƴ[o8H�!�˩|�K�5�����l�z���kj�����u�`��0��zMZ 2	Y�@[iʖ��P���!�-"1s�6Z��4�Ĭ�O}� ���%�*À�J���"��;�RĠ!��kxS%{���	��-/Wkv�s�=����S8t}�g�ٺ/�^�ؿy��o����]�庶�H���\%I-� B���J;+o��j�9"J[��շ3�ߺ�R�>�b������}�;��V��JP\`�r�Aʡt����+�-�Z��(h� �{`�ڹ�KR�n���a;p@$3XX9*u���W�U�@%[8^�D�ƕb��S����eMʢ���Yt'6~�d���J(oק��}��|:�k��a��++���/�f�K�j��-j+f�t�;G�^Ù�W�xP�
a�7�|�����_ ư����g�/�-�h��WI|*X
�s��1��ጌ�8e�e6	��\�f�68����ir��5��z�1~-s����s��t|��=N�<���uV3�/.Ϡ�|7P#��{{U�e�D�������%ͦ�x�7 ��L��WJ�X�w:�LXY�RM���:3� *p�KZ�n�D�qVU8�_��ʭU�k�R�r���HM�e������؂/�A���3�+aY'ֳv<0��bMP�j�t{�I���'�V�+oTErI�߾�wvr&�w�����D�Z&²����cN��`c�}i� �5N�ȭk׷�P2=]!p�.8m5B��Hl0[����jۉ�xze�|	 	��5�� 
&H�W_}�j-7�z�6�#N���n��~qz�X�����gϞ
ň�߿���۷��^)=����駟r̢�p��%][�*=4�h���9�nna!m�_���޽{�ٳ'�ML�X�:O��bq(�(M���RjU�5%����/�ʩ�r�{��"*��E)�y\T��5�ͼU����cwgC� �Z�!����R6�M�!�Y�@(,��y�B��|yʃ�7�9����2,YG�[�7�5��h<�إAJ�Uח�<�Zc�d�R[gr˔�]+ee<���g�k*E�Xpw5AG����p"�Q�v�w:�Z���gE3�u�w�n�?|<F���&�n3 �Q�Z�b*n>��+�bY_'2Y��*(�y�j˯R����%�)'�ڭ�e�VZK~�e݅���F��_���F��f�ju��I� AIz�`�7o�א>�0�K���W�T�lϿ�����mۭ�7����%�N��V��*��ߝM��bYow�r)�sܭ��, %�O��#$�a���^����7�˕�P�Ȇ�Og�$Su�2KС���:�W�\��N������N����$�S^�j��S-���:�+��gG^NZ�"'������x��t��^O>��fV*/��i\"��?VV��Aϗ� �L�`4z}|�r:t�d�j�]���rǖұ�zc8�� �uu�a����:�W@��>���������~&�l��8�,���ϱO�<��[B�=;�ω�����l��ѧ��P���A�����+��!ܙL�͎�-Iu>y�����g���`�"y�M�T.��CT?ݭ�Nw#������k�6���A��Rh�������~�����VM�/-+d�%�z����2���Sw㳏[ݎ2v��X���� B���^����~!�XFMZ�f��R:J����Foy����tىU�1KKԪ� HO���eI�����CUC��,��:���_�{*D�)�Clܴg�jā��ٍ�|���
n�T���C�Y�ڄ+�gbs9���V�&:26���0s��#0z��[��<?]r^�Fj��Sc�]IWh��Q<����6��Q3��2��R.�w�>�F]����Ck� �cg�����]�}��j� vaӖ�N��e'b
�!2h<:iVP�f���-b��d�6�8�l)�l�������;AbѕRW���jq�S!mk��+s���Ľ��pm���^��ޕ#��{���(.�V_��묎�j8�V	���^�LP$��@vI���zЄ�/γ}�~㬐is�
cŮ�ɕ�b充P߸�Etļ�]��"�h
�"�S'�]�j�D���Q�xi�ʼ�䍗P�}pomKd�4� u��E���*"�Wd}�J�&����*��[i5Uݒ1���zj�����3:���n)W�:۠܈@޵j_������7��pA-&~`��J��`T���g\G^$3�aI_a���&�h�y��,@���<}������������h��1�K�
�^5x���U�.9%.��(�����F�(q'e;�"Ԓ�Y����5�|�8���]����Ǯ�Y-�r�6fŔl��X�<᠀���u��N����7�$N��+R4�&Z*��cB9L_�Rz	t�s����ʬHTm(����!Mg�uBIa�T�jU6KV0t�8*ZӭyP	����k6���	����u%T�Y��93$<C���C�*u�r�ldN*W����Y�'-Y�X��29f\56�w[�H�3YD)n��~��R�. ᶛ]*�1���m6�f	)<+��!��x8ЩI�r
;y5�R�g�S�U�T��Q����b��R�VJ����7o����'~"�rgg�_SkTj�O>��k��R�F��^���7oބL�#��H��<�U5��䶋8�韄8}��8���*�z�����p���2J�Q�͉͋�0�\�'�uVM�ђ83�6�q�L�,�x*�9J%�N������I�����l�ѫ��ԭ���8��=جZ_Ě���hZ�X,�Ѵj���0N�g}C�V����s�#Vٴ�EZF�)yC��C1
o-y�����}5�I���ݪ/7�HZ�;(��~�"^�6�7.�D&�΃��������n�-f��F��f�.e5�
�A����qf8��:��?���>����cS�ݻi����{}2A(5���szrqq�݄S��%�NO���I��Y�5l8���\go����O�s�1��Çx��\ª6Ȫ�
(�X|jy�;����
��v|���c�MyK���I	2<�RN�� �����z<4���O<ob�Q�`#^�x!�YM�;���ja��z��@��a��C8�7bj��?��
RA�O9�k2R���Hѭ�2���hrlP��$���w}q��ͫAت7��g(��I�s%�p[*�P�J�n�]#t�bnyY&g9=���Q��]�.[�NM�ĺm�7��##����m�:̲ި5[�wgF�D��%��J	����Wj�0/<HE�r��x ��I�7'~��Q�n{yq���G:��U��9J�����)���t����ӗB'c������Z��#���ap���i�q�i!l����$vNޜQ9�+�{�!�P8I�Ea����6ܷ��	� d��SQ���?�s�WGg�����Y�6CBjW-o��`���#�~=~��1��ap���\��������}�Cxu�L��g3������>�h�~���&�\�dj�XXṴ
{�L(�@B;|Ak�=��3!�,2o�,5�F���
,)���^�P��m��ʭ�[�jZ@n�?ʷ
�R� Xe���}��!��0g~q�yy��6��v1�K��X���7�TQ=w�3�_%��.jZIY}:{<ũ��ʙ�U�#���s��*��W�?[��jp���<�QFJ"ݹsGԙr�\�9��o���իW���?������7oagŏ$�H�� ,c�}��
�c�;)n8�W/����0N�&�_��ݿ_i��5m�jI�$M���Ò��<w����c�Pm�'opq�f����O�NY�J������~�;!�g6�BƗ!�&�YXI��,X�5Yي�.�q:2�D��;��٪�v���c�X�r^4��ؗ+��e��e��l%�$\�fhu����:8�*������-�v���^���*�^�@Y@5��Xd-�J#g�mJil��d-��PI��"xwՉEQq���P�7��z�)u(�i9g5lje ��w��;�`���,�3, 4��ϩ%\O%4-,MJ�1ٺ��ۜhyzz�Ș`9�}�(&}�%'D!,�k�6�f95� �v���"
�߁��������=z4�%<��Q�s5Eu o���vC�}�aG"o�>���o���	��V��Ҋr��/N��g�qn�teT�Ym�?�P�ˀ�c�ɪ�JzI99sV9G�d�U����1(5E|JF9�P�Y�hR�x
5���[s�rXnj4U�U�3��xf��
|����+(�F3��RѮ!�!�A�����I���5
q!�ٝ�]lӛ'O�
��ꬪ>>�/�ʄO�2t�8�63���ZN���0,'��je��4�ϼT~J����{���\�v�����[������GA�����T��5�9=;!a���?�1!��z�����dN�<??��x͎SԻb��ݻwq?�_��b�� �l�ڕ��1�B�Y1����E��Ӎ.s���A@T�\���)/������A�-�SgFO��ؘS6s� U���wIBuq�x�8��<QaB������O��ggp(�1`�\[��nf���ե���\����%��q�͆�5yv�T9&���
K�Eۯ�X�����$�X���]rr�p�ʕ�M��a�Y��D����)�1��9/L"��k)�dZ*V[�sl��̅�ܿ�#��p���@����m����b��oYF]����P��p�s�,c�g�0�Hb|.5�z������M<^���[�V�s�:U��J�%'/Fb���?�E�oHy����4�rp��T���?j6�}��?�!�U�	,)ͅ�si��6�y�6��S�s�ux,K����"��oK��ܼu����`�F�H��|��7`�z��-k!I��:�k�:���W��--+b5M%�uB�$�]��	Q'�P��7o��Sx�Ѳ\�	��R&]�ȱ����ʒb���l��:�J�\h��Rg��x�.��ގՈ��˷>�ed��,ꏉ��� 0ȦZ�����`�8
U}as!Sء�B�3�H�}�%�.]�����B��$K��n���ׯ���n�&����k-�����T-��<[6� �!tJ"o�s��Gp-��bL�A!��ǖ��+�e������m�ƠpM���]���/��S��/~�AN�w�I�
�O+y�޽J���W��c>�j�����ׄAolB/O���>��#|���9�� ��^a������~�;����_�ί��HCY����I����7�)W
��N�'O���a��G������?�69}b�5/_�[\��7[;{�%9����;Ij��{p��#c7H�R��ä:�
g۹��ڛ#��Bʩ��{Q*�y�;���!%AɟL��D�yI�$�B:����J~	�<���D�@�h)�/�r�;�C�B(� �"�D��{j�Wb�I���2 뤖��N��Ui��JI���kДO�qi��ԥ�����Iw4�E�����K�IP
�-�ʜ�"e#.��E�QsNF���fl�I�hذnLz���h���݇�b���á�����]M�tV,G��a2�*�(G��]��5p�����ڝm�ۂ峧��yAɥ�����\	V���ʵj�Z��$9���gu=������=O77��(�V�A�:os1J�������������ˍ��]睕����|�"2u����g_��`a&#(���Xfd^��*�AB�r���8�<ZV+���mF��i��ry4�"��Q�W�\N�9-�O�Idd�K��5Nʂ�)�JaL�d�d@�NĴ��$�fK�jI[f~�Q���P�<W8RnU=#�X�W�JX��I��Rg:�MI-n���"y۪��K6Z��]�i玛�q�GK�X!��T�i�⌘c6��^��l����$��H�kZ��l��F��~��_D�۔�ެ�D4󫋒AD���p�Y'��7t�����7�|����lt7�f��P�������?��Ð��^��yyp\�����/����/I�nB��C�����xכ�F	�8�8T?��/q{��˰vi����0(/��Vm]_���N���f�l��Pv8,X{�����%5EI��t
��U/��"��wo>{u�.�f�l�ys�������ao4>�կq�yXIò_����E��wVl�ONN:[� �n���U�\3��>��I�L�����v���lyx(�W���0����#h��������<!z.t#&�y^LF2D4�h�J]n��E�ZYΗ.�Z��SZ|�'8RĦ�)>��T罛����&�^q���5o�x��hs��X5���#�z��ա���ܾ}�A��U$�f��z�.���5��8����T��� ��Wt��5o߸��1�
�E�>a�6�g�|�+�q�d��.c��^ā��G$�_/;[��r�Z:���)�j&#����Q���.��'��`1�_��^���=��l	�
��t��~�)e70~eZ��v�!1rdu����V�f�_{c�f�%g����r1�ssg)]�Vb�8�p�52b���])P�WwH��|�f�%NP,���9�֝C�8�4FsZ.��l����$���٨9OF�m��RE��]����\J�@]���+OA��JC���/&)��-�"�x�U�Z	}9�r�C��ĂP����L��wW�\"]P��cda�Z��5�E"��r�J�*#������ �ɊnD�l~/D��f�*�2D֛7g�t
9�]��v�e�1K����E��^���������FT���D��rQ&}��J���~��'?�я ?oNNlFM�(�u[�o�����?�1�,�A;�jKX#z��SHb(�4�����K���ja0+���?��o��5g@m���jNW���ݿ�7_|��_��_B�q��]{��;������`�&QIO��?F� �4Tw��7�7x��~��eZѢa/ȩnA�uJ1(o���c�S[?�>+ьW=��?�#êႝV[LV�ĭ���/��/���g�x�I*+�l�m]����ӂ<�S�,?�г�j�{x��²��VD[	��YП4������sd��9'���hu2kDe-�'V�/W4P]5-=�y*�C7b1��,gse��'`&�u�b}�fؐ����m�"z{kY��W��T�5�咅?�(���	�>=�K�ہ]̦
��*�.��0�^Z/��^
4u�]i-��֝����_���
+�}AE��zw���61;�q J��l���Z�Fƀ��!>��}����V�l��K���UϬ��(-��P��l:cgv�k��s��_�B�˫�S�_��jG����Y�k/��"f*��	��}g�A��Rg�沴��}����@ 拚��&��!Jn�8U�֝%�?n��o}�*W`P�U��14�c���⛤�jĐ ��ԑ��RQNF��ڻ�/j�e�.3ܕ:���r}oMЦ,۬,yM��ĵ����Z�`Z^�2#Ynf2�q��S,Qb��%TG��I�b��+�A�޹�A� |{Z
��� �����K,����'��/z�9����]DD���z����8��Y��-eY��/��# �d6_}���>�M5�	��B�������W�!����>y��=x_z~yʹR���8Z������)삘�T������ը����7:m�������|���-����5m�Q�ԣ%�l\�N;e��իW8���d4�[2�S�̩��ݽm��./�Ñ����r����8a�o9�GF;�mu���|?{��?G�yl �C'θ�`kbs��WA��̌�(9�gITf���m+�ٳD��!eu�_�Q�z���A)�V��29���l,X��/���㼜1}Հ㧧�"��}��k��|���V�S�ʣ�~ܢ�N3�s�u�09ur`����y8��r5�v�� ���ac��Y��¼��S$���(���8��4[ʃy��'q��Pq)�����.��S/w�I��\k��iB~�Lfc1�Vw��0ٓ�gb�j6۰�v�|��02������is�-U �n��^3��9�<��JOg����S,��	xG�!���ѣ�%
q>W�44_��y�����jȪ�o㊳��������Y<�`4������7V��V�w��GM���Ui�u�WqF��ߏ��b,�'���K,�T��NU>��/��C�dV�Cw"s-��>&V56�J�ꖰ�l�e����	��d�.t���;f����kB���l��������Μ;����h�x���x~�����x�B�\
tT��o��YZ�V-�˿�{�ώ�Ծ��������}zck��K�M~vt��
$���)vC∴7�c�F�|Pz��`xL<,���1>�w��W_}���~�)��I�j�.��]��V�������������f���W/���/�[\�w_�FHyŗ(b������۷o;��_iL�Tk���j���'����G|���^�
����A����dɈ<'���II��� �z�#�Ӯ���4~K�f ���k�"�zY�l-jn��������%Nl�5k�?��(�[s@'��QAQ\pN�Bڪ�q~�a5�4�xt�eQr-T��$�[U2���+�RM�*I����`/f�q��^ߨ3�Ԇ6¨����v�ŰF��������fwkc	�,�����%,��ǃ@̘��F�g�XM'4'��0u��5ٌϵ2DW�`=�U���a89��A�a�G�N�t���^#��"�l����B����]����׽	nۉKh��"Pg�)���FwKB��{w�#3�XQ���ث�$Bfj��|=!�����t1ܴ����1��Ɠ�XB��;C:�H�\
\ʮ���ɜ��+JY]��%Ӵ�1�X�y���^ͮ�>�P�DU�A���T��yv����wĬ+(��o�#*�	��U2���s�N��dѫ����X�lKc��=����,'��,=�Z���`<��LMd���NQ�qG+�%#(�ɂ�V�N��LI��������ѳ��?����c�a��B�*��bg��;����&n{6w\���c|�~��.�����t2���+4L$���?؛\�ހ�����o���>����'ЧP��<�����aO�����F�	�$�^pN�6s��d׋8RU�,8��jl��FG��^ã�Ǎ&D�4�7���[8�q�R����<]�42��)�%�c���Z���>���m��h	����e��<�y�(;H��g�Beǌ�9��o]�8!�.#^�J������n�"W*f���Z=�&����{+\�}�ׁ���1'\����!�ͥǲYoݰO��n�Q�yTֆ�V�����W�W�oyv�5a�9>�l9Q�X���:��Z/��e��S.�,84���H���	c|p�#��!Dx_X��r��VL��OwA1@�`������K�Y��t�w�ƃ�x:�~��^-W(H��YݞV<Ogӱ��!���������`n>D��57Y�Z�+�p(e�=|������2I�Z��L
��!��4|B{�$��x�y��{�I�D��7�������Љ�0ݘ7�ƛ��$Q�"��
��n�T�h��N߆�<���F.[�S��^A��=�x�r4��i�%+2*�j��	"��a�d�d!���9\���P1�_��E��uթ)��w%�!�/Oy�M7Eo��1u��%9�jP��	yu|
e��l>�q��f���|��yv�'mįm��k~�e�q�=�4x���ӕ"�&�������_~	���B�D6�M��Bm������r�F�����R���c2��'Bi��p`��)��I�mǧ`�`,�޼��__�V!..��12�r,Dk��r���a�fரh���-|�\��Cח0�0	j��O��ub�Mǹ2Ze�փ�h�����窕�/�7Zg�Z~�����2�|l���[9L%Z�X�V������$����X�1OB�`m��V�iC|�i�tYʡ����M�H��h�9<^���s��P����ͬyt�  M�F=�*��k�X˫,��g��[�	p8+-�0i�UR�#\�kE�{L�Nڈ�d*x��2$�:\���c;�%u/� �EZ����!>p��蠀c���:�Q�����k�������a���&����ݲ�XA�T�L��(��sE[�*�2�E��&c�ΎȊ�q�;����44�+~�����	�}��f�݄��Q��v��}�R�����؈��,aMr1��γ����}��x����٪�~�H$��]C�d�{�6���I�n�M�@�G" ���ZG��0��U���D�'sYp�����VYfJ'�l1�6��z�q+���ѣ�d�����j�Q��7+�SvuMS�f.N�����T\Q���R���֚���^cc�������P�+�0h�,�cN���S�SC��r���~��y᭨��X�xW~N��۴������k�L&d���#X���<z���	I�juf��V�{�!Nc�����&�v8ya-s��1�������T�h�db9�K!��=|���u;�.nc*��W�W?��q����0c?� �yyz��l�[Mܩ�ha��,�uxca�J!Ѵ꧃����B��c<hy�7���+��#x4�Z��Њ���g�!�a�~����~�Q�4Z]��a��"���LOG[>����ݹu�md��e��9?�z*�K�h�1���A�̹���&��i�X3s�P�,Oq�j��0�,-J}���0"U�b�Wt�z�	�#s�E��ڼ�b5��b��
��9�p���:u��T�B��ҳz��*��2J�,(s�'��!�֔*���kf�Z��i�]�J�t77��2��lr��/�?~ջΜ�e*+(�^� �SB��θ�5S�`.�c9|�ջn[6K_�0���t�d�G���jS�-��G�lt΃,�]n~U '����}����@%��難W��bj��T|�n,�3E'a���k�=].�U#J��;�PnX���R2թ%!�pH��k���.ˉg�җi�o*e_�9����E�lzU68ӳaڳ��_�H�p,W��j0�a�@8z�Ӊ8���ﮋ���qx���66l��hO�8@YN�T�6�Z>#��cצ����� ���Y�����a9��"{�:~�%��z���&���ѡI��G+EcA9j������>w�����P3dĚͭ�9�˖�j��_�z��c�}���̪��E��ÚKh�G�~��~��_B�Ǔ)��YtuvBZr�i��&c+b`g��Z(��X��?$h��0%�u���=������mX"!<��q"�����_��O�ӏ?�w�.>|/��x�vW�_���ӏ>�H�<��Jy����o�E�"Ls��Ue$�|�f̹��L�2$� [sF��em��RAQ�nPX��U�-5%���S�:n�����Mm����bJ��L#��Q*Y\�t�خV�Jr�Y1��茒ur�,5�:�M� �J�J��u�Ja��%ي9ʳ���r	p�KCR<�e�(N50T�6yKxChqy������e��\TH+J�$^��r4@^�_����	�gCS\����^쯫8Z����o=-"�Rʌ�OI3�^I`�Br��A��+8?��el���/���\ �s/sc�R�(8Ƽ@�k�E�o-�p�P�r)��R������J��o~�F�]ۗ��ԃ�Nv��������L7��|�����}�����"q��F�������qG3�B�B|4a�L���)"8���xw�ܙO�/�Wa� l�k�V�����]S$GC��ݻw���d>�Xyߧܔ+�|d�g�*��in��`��t��F��ܑ2r�.뵪��3��J��nL]�a���{�LI�X�l`��W�I��$Ԭo�$�|7t��ޕ�6� A�Ʀv��Y��4�u�Ͱ;/h:x�;ۯ�����j�j����<�Ӿ�#�Wx: �6_d5Z���ƽ�!�c;���h���t�C��A���8�e�/���r��8���g8�o��[?��V'usJ<x�(01%����$$�v}����	GM�a�z�(<,3lnF��g�5v�Œkm��
�������aAp?,�.��5��]'k49�d:���׸y��WƠ�0 E����h.<��6(ˊc//)!��X9,\a�x9�A�Ź�V�6� ΅�&���R`��=��KE���WUbs�N	<��^w>�wpp�|8�ӇȞ�o(���>֕ͳx2X̖ҕv:��P��^�t�㢎bz!� a�zqS��䕠ʌm�3�$���t�`���>��م�*� ݂dM"2xH{=�#Pv��.'�}��U������B�]�%oŸ%�+;��L��n�����zM�O�Ԅ}.f��ݿ{��n�6s�0�vK�N�X���9)�H��^���K-���\��d;l��Ű�;�z�b�L�K9!�Z�9\�&CN��oquINh.{]&1�%� 6fK��������A�Z����2^L5��.�=]9��Y�W��a��^(��P��e҉��#q�d��ZoZ-*�
VVZP�,��`��[*v���!)����9��Hd�wG��c�"�����q�U���&{����J��dQ^0(d����ۆ��*����CI�Y�r��I[U��G㋔�J���Fu2��ߎ�Y�)�@�J�V h��f�(l�ןpʞ��N����(r��f�29[�������c�.V�<Vz^�����X<�	�R��xpՐ�N���o���/A,����x��[�|�A��[ұ��h3�H��-ǥԟ��A/�đP�O�_����}�/���DV
�
g�ٳg�|ά�Sy�V�詳�,D��R��_(�:�2��v�F�_�Ld����^�Μ�q��l2�pW�a�t��u�v�`l�|᭛F.�HD��|/��[}���'����7�|#��x�����ώ�ٕ`&2�=<o�{���l�[!�6v�c4R̟:�_���Hӣ��نd�]d�e_����G"ݞs rF�ec�F�d��g�=�\��{ơ��f*��:��MU��Ʒ&�k$?sD��V(l����ۃ+3�͍�e���Y�KB��Y���_(MR�ۼI�@ܹ� =$���˹
��X����T�a�`���s9�Ke �C�;yr�eLȍ`���);"�g��7�t"p�+�/f��k\[�]JU�E�"*c.Y4I����9Z�c�����j�fI�����7�e2+w.دυ�_���e6e��bA]��ׇk��^����眯�𓉁�*5Ee��(X�W��v���\�Ep�H�v��	T�Gq4fD�ޤ�{x|T'S�Z�9�U��W�,�W�'EJ�����~!gH����E��y���Iyh����׶�����/��AG0��W�0�+�pm��ӥHf���QȳV)ONɊ�f�L6�;rA�]�"d��t6Z��h,�(���6\v�5cR ���ʐ6�����b���~���lpի��kk\�Qopvq~5�I�>��CW��B��K����N�N������&�"��S>��#M�����9�ÙS�G����/���[���?��o��{������~���s��V�o!c�9{������o�B;i�C�4	����߽��i�W�#��Y Uo��$�\�O��ނ���e���9xs������_B9}��/!��v���c.ӱ��}wm��/OpMsIK����v�_�WWi��ys��j6[Kb"1��0c08؃~�Յ��V���� ��S��i�f<<<�i���t����jU9�(fxa6�!��'Y���mk�����o���˛GpXe5U��FdRˢ8�o�c�֢�E�i쨰��ٓyJ|�U�yI`.ĚΑ��T�~�_^MS 'l�.m���v}���z#�C���ĵz��wݢY<���>�/:5*]+ ����c�p-�%�;y`v�r�8u:�!���}���|c��n>�Q��y�m4�r�F�D�֏�-����3x��rS�Ww�9���K ��}Q_й�hx��br�Y���w�g�������b<'����Gp���V�Ҵb|;�i�a��b�
�`��q�8@N���=$?^��K����������\�<!+���Ē6i�&�DeF2�g��j���#f����7�7��ن�c���E��;y؆/�>�!Wz �Y�l�r��4,��c�,��5��+�Dj�䐫��4���6JR��̪�������P�8��7�Dv� Lв��V�XJ�C/'\MF��=,{��n{*P+��3^<���D���2@��i�hc����S&$o�ͩ��ij�ȋA:�,�d�U�U����rm{��?>z�B,�ϟ?���ΡĬ���[R���zQ��Jم�Ǘկ	߄V���,"��b�������O
�R$�г0]���w���	L3�UN�6o���A{i��~��P7V�%��f1�+U�?��|c�`�B4���ŭJۺ����.��!�uAE���!k��o����|����"�_��D���0�`բKD:֏z��K��yՆ��VK5Y�b�%��N����܆cl}K$�v��1��Ֆ�<<�U��WL�.ʶ��'�j���U}b��*T���U��P�bK�}���
�t.��$S�U����RSę5	�e�P<�RV�(�hY'�����!�<]�i4T`J23�����^b�zA�b����\{ ���a�i���o���pJ��v����mie�wvv���[|kg���5�a�((���5qI�*׷���f�V~�ې���XT@PRfm��Ey������vT���ƽKh�v��9|���C(gXX�nܕ�,���h<R>���8�,A�?�k�6�|q{gw�&��.�
���`���ثr�&�qO I7A�M�ET�U9��O�=|��L]�?�sO�=~��t��5a��0� �k�d����8���Y'Cd�*�u�$ã�"�=�Z��h͒�ڨ�\�#u�C�*��t4�M�8���4[��E/(é`�K5�H��̐cfE�NV,1��i�ͪ5\*O���W_=�j�/�+MvL*�h�����Z���{�����K�$.��I��|���._�W07�l �y�Lzq���|/��x4L�ho�M+��?vL�c�Z�Mg�����?��������~�k�ư^�,� �v{��I���S�'�Ū�E:�n��ld��Gu���Ƶ�ׯ�Q��%|�iس^嫕J�V��u�bl���BqܺuK{W3���Q0��a\�^���2c�=owҜNǇ�|���������|��^็�g����rx	8���3�N��	�1)5#OZ-}�aT*gd=fU#18����P+%/�܃��]����)xҎ�x7vvq���Q!�k��HD)-T�*vF�uՐ���Z����@����l�!�F�1�s3W��ٓB��9&��]��݆1�M09�	��K#�@s
��<B��/(աa��U���,�+�[ޯ��a�C�T,A���ǃq�/l�m�|��r�U�,&YZo6���$�*պ`�L�\�Z.�����a2���z��뷊�z��'��DY(�a�_a&���X�7���:̵�mjU�:��8&��S1ǌ��ߤ�e⛷�݄��V��&��8?
U��`U�	�#Y,� �{P���N�G�[��C�(BI�d�Э +��yq�m5�ח��*
���΋k$a���ԧoԼRH�(ԥtld2(�"�a!����خ<�W'�-}�[�%�,�� ZPO+/�Fs0��1��(/�3�����o��6�V�����f�}6N�\F0�u�~����7�1ӄt��B����O�˳�YE�X�d�nE��,�<�1�h��˥�8���ؔFB���V�� ����ʉ]77!��������͛7��_����H��>� �'��Bok$2�Ow�Tjm���:�b��V�����}�]HC�?�&ݜS�As��b���U�+G8�R8�+������������?�裏����C�ɶ�ǧK�Z[E�`bgM��U��̍lc8�J�n�>��tS� [�#;Nk����Q����;�Y��ѫ�2�EE�c!H!!�<#}R�^��!��Ӯ���(��Ya���:��S,c7q�
%X�'���Q	SDg�'�,�c;���fK��Y�zAӗ�`r�gf�i��}jR0�j�+5�sX9�f�b�~����Qv�[�(Á���a���MsL�cTϾe�._`��Ƕ}=.N3O�"ɖ��*��*\%!���kT6�B[�t�G�˭�����"��뒤XxYR�lDLV41�J����Z�2�=��_�\���?���ӵͭ���le����c>���ՄCY)���[$��/�[VX�tr&�/��������_X�%~��^*�����YC
�,�(�&8J�������v�=�D&�nךL󲺭�P�O��e�)�AѢ��.�ߨ�v4(�*�N�Ǹ��ß�dt~2	�0K�hc�4[P����3<X�Z�\��U�.��\�JH(��	ǡ�O,�a�g�J���jk�gZ�>"L7�����R�0��q��3;9z��\:I�����7nB�%	ű�t�r�b:a(� ��t�JEP�Z=srɂ��S�5V�$�]u;FT���t�..;�,n�S�Z�T��y�b�������ޝM×���:j��(�BCD�ڴ(o.c�5n��(Z�OMX�a ����/�7�� ��ި6W�_}������$�n߾ݿ��,��k��P�v�̇sp|����n�ь8���vbo�����3|���p��T��/�>�<-�����W��Bs�&���Tk'g7KTP���\��L%�G�H�=^i0�FF`c9��H�:���?���,�l�|�j�b��:]�����8'd��d���M2���={��Ө�'*ڄIo3�8��$�{�_�����=���_�x!��=B6O�@���'���&��S���.T���2�q��X��o}�ގ��$i�f���9_�i_�l3��V+�`����"<���!��ZF�K2�l]��(YמkA��ꂩ3+6�o��a��K���5!L��hrp d�������J�����&��X9t�Q�9vqL/�Th\����z��am�TI63�V��s̏�٣s�%��G}	t�ƍa(��9eרn����b�"����T�}v�(V���rBs�9��!�¯,i+�A�ΙC6��T8����^2��	t̤3����Y����g��RH�5��
V�e
� ���*���o%���-H(�b��$ˑ�Y�3gQ8�y���Ԝ-Z=��WW6��@�I����c�@l0���L�9G޷uɁ�Vɑ��j1�Q�uk˄O�z{~���K�g����������r�}�Ѵ�=6�

LV{9֬s�o���_��_�on����0@�`�0$�/3^kk���� �ؽ��� 
~�����X=?����}9�𴰋T?{�����NՓ'O>��,�`T�\�U1�
����\��@�)��^��uL̱��0	T�[��	g�E��4���(�qt����m<3�k5_��>%��a�e��J�2r��!�`&��:�+շ�֜������"/�>�Q���m�.�B�*fFَ���J���W|�O��M�&�G�)��x9ql��`4	�ⷩ��e\�`)�p��>��{�����M�<;�D��eɽ�;h�ɏ��:�i�AI��e9�Z�cS侘�(%��MW��ׯ_oo���S���a������`E/�A^9��O���͂��h�"�2��Y����P��,bK�m]��;M�޾=�cN�lw.�?��4v�l������_�=�Z�Z-u�tlk���'���0���7�6�C?	ˁ[���N:yn�Th�u�g���7��Tj��1�Z�%�O�v^2��Њ�C���l�/�7�6��{�����|�Y(�b�;����{��ǐ��6��I<S|gVceՕ)��z�22l\`�T�{��s����X?z<pP(Ƴh��()�K�h�1�ċ��o��,��9>q󾅒i톖N���n1jd氆J��b'�{��?��V,X��d��S?�N�����l�Tk��^�Y�G�hF<��pR�FQ�fN�l!�,����U{�ˢ\�d9��v��x�i��YyN.6$��<=����VJegD����O�j-bUݠ����]<װ�%{M�Pn����?��3��:x�\��i��&R�}�5<�Z�%ԛ�p<���,��W���xk�/���76��nyA!L��x�jA�8q�9|���7�0�={�Z�H������o�\�]�m��6�Kh>�+����)���7X�p��E���f�����w?x�����������7^�zszp�x���z�v��������V9ρ�'�U��~^�R�	!V-�%� �(�h�j�rl쒟�f� ��i)�>c��r��r7z�S����O�a���3�r�>	�q�D ~i4��(��4�Q�p2�5��k��oWʁ_+�%�4_�1ہ���d�ȣr�����M�g��"Kg�oކnw�[�0�덕��l6���I�9%cno�a�p�1����f��MgE{��h��#�ҵF�/�ꯞ?��g��_�>|�]#)�˽n�:�ہ��F��*W���L"yߋf�F�r��u�,�Ǥ���ؔ�n��	ʂ܍#O��Ӑ4��J6��=�X_�֛�o-�R�_�߽��Y�id%�Z� �y+r,�ҹةU#7K<��׃�j��:�ڷ(�j�QoԒ4���
�n� �8jml�֭�/I.��F�Z.:�G���Z��P,޸y3���Zukw����1,$�<��wc�1��\<�3�1<`�F����%�lu{�O/ϰvv�p�ӓ5�%M��v������u��22�Von܀sr���c�n֙�vL���V��.yջq�3/��i�����݅8��9��f��C������R�������"Ør樟g��,���5� �g2UL�R�mݜ���1J>7�
�ń��nÕf�W�	#c�4T�L��_�9���G14��fU�q��6��S��A%(�E���L%
�M"&�k%���X�\J�9v���=�%�%��j�ƴ��)i+H�j@A#8ʟ\t�8[ka"~]��zu+���A'Ot��"KO�~bq��;�)�l� a��=�ʅ[S��d�p*`���X�����������c,,���W�X� `����۬9pXF��_�w,W������@�k�+���z�L��^Cd�B�`�xj�3T���6��ɒ|˺_��me��h�fLL\�A+��`Nn�@�N���`J����)�?�����	)kC�:�g^'Ġ���S0��Ζ>��V��\Ga%�-��]�A�S�)fx�N���:=H��8�fC	 �K?��!����b����lѢ�h�0��s�|}�
�s>X����{������6���z�2s�h�p.��xH���G��z{sK~�$$Udo�JY��J��y��S/N��q!C���n�;oUg�EPo�b��\\��\e����e��S���{�.q~*���d�V+#�	�,x@�y�v������`�3�ؑ����D��_��@��o'�YH��v��9�[{6qE!�q�qFj��h���1n�ز�k�+�?RT���c^@Xa��/8Q���ݻ��_=�,�湷����!!"o�j�[��n�����䀧�����0,G�jY���!��F��C�2�E�
~���s�wQI�[P�Ab2�F�eF�!�
�̒��r���˾��쒞�#c�~Q!"ek���8�2����iȚ��tvpx(�OkfQ�X�Tj��
���#��r�dU*� ��J��/�Ho&���9��.^٢C�B
�B�t�ڧ�猧�3��4��Є�Z*�C���*���l*D�
�,mARX1��HÔ���,^�Rf�l0����xu����?H�6�g��Z��6�*t�d2�tz���g���/���������-~zz�su6��BP�}��w��`e�ꗿ�e�����$+Pi�(��N��zcsc��ߺ	+H�����ﾓ8vu���S���"��˃#V>;��%�����kk��%�Az����.f���qj1}�_�����\�yc&�qy��R�>�Z�o�b`���(��"�RvFc��gW �Ɏi�E������/>�����Yǵ�i
� �&��[ԇ+E���ZD%�B�G����J�}ٹb���l��ݻw�Pgg�X=�c���uҮ�"��j7�N[�p<�S&�EL��)�f�&
*�\aG�(�'��r�*5M�ŉ�7���Y�l��&eq�,��%k�T��b"�	D�c�)*>��4�jp�ܣ����>���tLǔ�n�&��Y�K���U˔Bp�Hq�A�O���f\n�b>��Дt~��C�J.�-^��TpL�����*���PԘ8�(V_t�
 �L���wO3�Q�V5M��A"L&L��<��|�3t�
�s{{��o�������������x���o��S؀->��<Ã_�e24�XwΫ@esa��i咀���P)2�Lm�9���a��Rm�T�z�ZJБ�ʫQ_���)��d�c^d$��މ�M04�*��U/�k��q�Um���;���隒�����%=�Ԫ���8�'�RK�1��g��5mD�V���rY��l麾�?�	�a9^��Ӂ_:)Cp3�<�3�/��v�'�6Vd4"�X�s�������no��.Yp��HIՓS�g|�B��8'��LFl�J��Ç�`�oჾ��=E�1X&�۸?��E
�ya�o��Zs�1/3�Zi�W�63�]�e����_��r-F���*e٧��%έ7$7�G�/�zvt���^�s����iI�8�h2���0c���X��Z&ƣ�!�Vо�8��DG0�7���a����n<bs�шe��">�>15*wUX|y�d4`{�X�ȫ=5���U�zuRQ��6�h�)�g��)ӣ͉9���&_n��H ~�a����)_��c�t��5�jj�kmפ3㺇����u0$����������L��y�Q�9����w����p̉x���X�.���{{[�/g�l�-�}��(�<̏�V����|AȽ`mG��̓1Tf��U!ܔ����鏫��-,��w�w�ܩ��7c�T�)��tDe���6�KBm�&��8�'=e����%�ߐ��n���
;+Xȏ>��c������|�F�ڼU��y�,	fn���x�?V��Ҿ�;ϰ��3m�&��2���۽���d]�7a�E��F��ExX������~�NBۚ�y�X� �/��\H8�,ݚ�

15Ix耽+�Jt�4R�@J�=E��	���
�y���R�p�5%(�d^�+��`8:<:��Zr}/��gC��(��{��6[��[>�0*���R�����R��_,`��'l�(�������!� @:���( $Jb��(�T�J�)���|����Lcc
��	i��"��(��܌��@s:	��1�Þ���9�Sq>/�J�j	,���\1K��|7��k�a=&�j����srx�s�\��α3����,���'c?���'��&����s��W��[gɾ�;�Ƅ�۞��� ����!(O����*��	��D��UA�H���P�b�`�lloË��Y8Y_eO�n�;#�4��*�U�K�^��"��ε.�����zd-ˀ�T���p�5ᕯ:��ʂb	Z��h8G.���\��M�
�����	�������n����kۛ�j�����������g�ڗ��;;�G�
���É�GC����d��P*��`8(I�ٶR��9���h]���^�%��`�W�J������p��V�OR��.T�*�޸9l��1�G�\}���g|��q��,{W�6a��
E8�E[ l0�L��|��uG8G��̋�;L�FA!��W�6e�3��4_ & [t���Q�TK��3 S���&C����p��� �Č�{�SY�mo�z�����;إ&�
��e��I���FU2&\d��pRlHLL�J���,��2N��i�ĸ�츕F���1�*��p� F�Ϙ·(F'��?~��x�����2""+~<��|�I�#!�?��S��������W|͇�b�K֣�ʈ��0'W]B�1�P*�<�"�.�'�8]��I�P.ɐ�c�r��e�� ��ᰏ�իU٪,�Y_S̈́n��J@ǔ��Ň��b�l�c/wn/}fE��El��(Ȁ�dB��&Җ�ʛ��$�hA��c�^�5��1�͒,�Q0��Q�Dl N�����ի
RC��������7�fˎl$�-��4n�1��`�|!�0�6G��Y1b�L���NYKY�_~���{��n}��;%���|���?���������O~��pX�⯥���3��Q�_�R8j�!�!���okqh/�믟`f��'.;Z��oFN�*��O��Jk��Aup��Ə�)J��N��gg��O�opSތG�����K�OY'�%��1��r���/��jj@�zM�M6��
����?�� utlD{��<����O����v��P*���#W��j 1W2i��UM���<(*b�!��Ģ?o���T,�O��U �[x*Lf���G�Z9alI`�R1�ŋ�_�Y��#2��ڻv O��O���X�r鼇�2�~oKde�>3ņAbnq����F���!��7�2	����/-�L�Q��p4 b1�s\6����`5�e� 6���Oc�WQӨ�2�7�΃�0�~��+K��\�I�0Y�J=�%��q�M�Mu�l�|~z��4ṣi�Md1�+�>fF�~x|[�d������}��٢�cR*�����/�U��b�bl��>To��/>k������;Ｓ��eo8����H���j� %@�����M|2�ҙusMx�����rM�����U�5��0�G�:l�c�Q�85K�  �y~eĢ-B1�,�:H�q��3�ȗ|�pxr�݋����ƺ�����N�HG�ɬј�LQs�SH �q1P\&´Z�]^�eiۀ�;�7e\=���UH-Ѣ��9Y�����8�ƃZd�qmk�T.�-X}�������+���*����W���&O#�L1��}�x<�'!����D�0O._�Ԓp������?��ق��+���-�
>����������������/�@�Wk��`sk=u�>d��/�F)ȶf���x5덽��x
v�4(��9�r��C5�|Y��,�^�ف�dX�mc0�VJ-Z}�V�[%�0E������/����ܪ�䧾,+5użk1F%�)��֨��l���;~!2�
iT,+3��Z��
���pjM<�^\�1��&o��ܻ{���{��ӹd���0Kb�Ƒ�9�t����)T^0�4>�KeSc�������]�������狻+���N�/��`�֊'X	KV�E&[��h�P�͚�
?���I����%&[;������>�gR��vԼ �C��%k�f��[+>s�n�ed�z��߽27w�3��tkw���K��
�ʨw��uYP����Y.`�2<�t4.��i�����Ё::zcPj:��0�X�T��6�,�7<� �}J\D��
��䃃�y95l�r�l�#��C���4R�"�������<��~[��2o�@�gk�S�u/E3�0I�6g��R~���1M;;;8����u�_�xn'nS�Ec>�>�-",�T(-G[��RaY:
�2�X�7g�KA���
hD�֋v�蝉���bA����`N�XV���.���,��H�d��ȹ�X���	\:�O��l������(��Ȩ��hl\���$^��Qm�i!�Y.�wʜg�=�p�����䔻�����"�$���v�_���</���7��$N�4�'�LV�C�Y��f�Q�(U����74%� �+�角Z4���'�>�1���[�+���׿�ۿ�����ǯb�r�����`'X✇���mw:�bI癎����`�����up���K8���{����{�!�g1�<k��W]\�ѣGb�Unl�O�_�z��
�j�1:'�!�����e�t��{��}��4����ZPZ��� wyx�6V}����j2�a���
�C���Sk����3`��`����ْO�id���@5}��ok6�,�"<��DY$K�1H(c�~#��i�a��߇FSRw�ӆ�	&���2:�ee�����`+A3�#ф�-:�o��t;�1x2��������%���|e����̪�06S��x���j�R�z�ׯ_c�a�a5����p�W,7.���X�j�t�]f���n�ؖ�Q]*�.m[jP�n��AkF4�6�U�8�Ե��&Ý�L�)Ui�dOe0����,��Vs�������׏?�8ur'g��J����:�Nm�G=����N��{�,`�꫅��t�qk�U�r�ѬAd|�m���~��g}�у��Qp��E��DQd�_ӆ�t�Xs��"nr�]�x̬i�~���_�1�9<o�Y�Ŭ����T���D���Rm:�H%3�?��+'I�C�(�����������0����j�y��3/���^K���%�d��{�`���׻�
G#���B�+Dn�� �j-n�cF�H�����y�,|��$$Ў͈�*-K�N��e�R�#ع=<%����&ݵ�{���d@���{I�B�i�E�����ZWjU��.I0�5lb襹���'EEJ�n�Ӿ$O�Mn�ZŁ����)��T�ʲ2EH�_��W������������o �U�^�o��F����޺�g�C��(J�y���E\����xt�V�م����W�rY�HHm<ΦLp��
���
�Ą2�f�W�%�;�R��hv�捋���xIdt�	|�r)�N����o4�4]��c�c(���
A���G+U�4q�iT�r�m,$�%y�N�LIj������
g�"Yiqvqy����b��`��_K�t6�B0����b.P�B����8��Dk(U*i�_�u��}�&Ll̀ ��Z`�)��{u�=�=�'�P3�����xB��,pØ=��X���z���_��N�`!^u�G�63���M��dfe���
��x~��Y�O���t�9���ꍕr�>�Y���)h��"�|�����N����J�2�qʰ�M�G�H,�EJ(^Y!��Z$�z{����~��|��1�^*�i�?��=Sm*v��:��ئg˭��c�=klrwa��G��Ó=<z�t�@q��r������ M��95�o-'���D�c٪���������E�Z<i��T�����Y4�q�ƭ�ױ6�}�݇~ج�VϜ�P�I�Y��&���,ܚFL&dTeL_��=u&��RkIw��&Z�7���^�����2[���?2+��Xm���RA��w`�+�8�`-
�Q�]�.Ê����2�'di�a�t25~��@���D��,0��t���]�:�5�tQR.�ʦ�W\aww7� Iqq��@X��pZ+D�7*��U�ʅù���_#)0�=�
O���ZsQ5��<>"���x�t����U2.h�������C���1�����^�b�bm�wH4̘Pv"w���D�;p/4W��d!���Y��Z�'�����xS�~ͻ{1��N�̜-mQ�mw�F,a0П�T	d��{]uY�� ���-j)s�'�G	��&���r����ln�y�Ra6F;������b�U
�ȋ�s�PE�Nb6���w���-��0lL������ݕ�N���:sn�~�C(֍1���c����{J���|��|D�;������仆��G�e�LP��[�E�5�����6���������د���k�u�t��1D��J�Z ��B����a}��'��)ac@0�Rg��}��v�
F1��q�`lJ��y�9Q>�7�������q��B�xKV|�S4w���B�̳�������ɹ(���O>QpٱzL7���������駟v�:ЃC��G��w<��&|��}�`��o����bL�a�U�d�Ԛ�;����5�*v*��ݭm�x���Ϟ�x��]Ne�P�V<�UoSr�g�
?Lil�x�����U�7����}�p7EK�XoW�i0���@q�%��Ꚇ��W�u�}D0�1A�v��"���k��˯����j��(I�����.����m5W+�v�Z+�s�B(�L�i��`��b|�?�"��8�{Q��悠��d]��=��#8&���7	 ���U�Sh�����}v�����q����<��d����s#�&D��+IR�c�C�#Ԭ���d����jc���J��0�!�0�w�ͼU�� ��76f�3&�i�)��kN1��n4w۝�����?������#9?;���{;�[��'o�޽���
�4�� �o� +�by��S$~V˦N�i��J2��s,,�C��ƣw�*ؽ��v���6���O�J�Q�P���
Fձyv��ᓃ�S�2���!CmQ䒖y�Xt�j�Ń%�Ǝf�ԭU�Fi��j��GM�K3E���"��=��,�C�@k_.�q��P*?|��p4}���w�^ܾ~������/.�ׯ��I�sT���M�y��&H�0)��^�a{�4�jF���.�]Q�DG����x��?�RJBb���Jc{��v��^�~���E��f���B��J��Y�b!��a����C�Y�ܬ�7� ����<��p��Jucw�����_���3�8�OeS����s6�&�14"��B῝����m@fµ��A�X�ܨ�|�JL?~�'����DI�����x��yw{�}v��<'s!Y���� KzǓ�p�K"��V��K��Icp<x��\D�7���Y(]Ȃ����`�wz��RTV��.��x�k�'�����;��|�ǣX!?8�W��9�$���f�>�ͨ���o���������6g�p&���)X���� �՞����g����;00a4�M���I�j�xѡD�y ��Ԫa���`:������Z�.�j��s^Ac'6!�V+0��p5\�L��� ��h�,��Hwqp�+�Wi,C3�Xd2y��A@�ٺ��aA=k}C����^���,0��;ơrb��eT��I"(�$��㊞;�5�-ʼP��*����뎭�I�ʦhf�FIQ4%�ݕӎp��2����D{�:t<~�+�)AI�u;c���Asr�Q r�0c��Ye�Y�dw�u�L��ZP����Hspzj�J�Ό��a�qS��[/�/*aa70i��
|ߗd�q�����۷�#rY��~gg��J^��J`�$Gܔy�E���`2VQ�����n4��R�
O�*���W�t���l5s�]�"��akU <��\j3K'�*�<2S��0��}�#�����9��͢+��?��OO�>}�w��Zp:9;W�Ba �6�P���b���Z|��jE�4/9��X*���5��Ǘ��W�ьX�x���AW�3�'UC��vww�{1��ghz��E	�.V\��L�e#g��m�1�;o��4���Y�I3b1�qb�&����ӳ3Y�8J�l��r��V�ǿR�ɫ,jV�/�C̒�$k��"�Fʭ2�g�Np$�nYo����L�/��"�|�� ,�@/�F�c��'C! ������;4߆<�;;88�\�cEU��a���p���Z��/|����ڵ=��B1(���%���z�3�ޣ�����?}���'��ݫ¸s}3�I�Pn`�R�N�=~i�TI-��ߒ5���PGF9�Ō�AP����.X�$���+0�A��y�͡����d��9a�64isj�o�#����{�}Ek5L�z�9����>�]|��-b�˴��v2eJ>�Y�Pr��]UV��|��T�z�q4���П�����;���&�ل���'���&���
� v"R����c,C�L�A�{�j/���٥��]4�,:cc����#-�<C#*%���c�{�3�_^I��,ɉ��g`	��8?�R��I��~Ш����?(�X4��}�#����������>�V.�Y��w��d8��˗j&��5�U��:���f�꠿����c䥯09�j�t��,�RU�|����ۅ�7�Ѯ�4-��u��*,Op���1\4�^��U�OA X�`L6�b�"�T�;ųȮ6R�/��a�C����zU[V�i5%���fr�n�8�P���e��	q��j������%�J�Riw�O��(��9`�<{�_}��GFډ[�Y�~V�e��Fb(H���x4��c�Tƞ�`!OhH�lt�E�;�@�j�}qt@櫵�U~R�ݻuks�_���ӹ�*,�Ґµ�-�0�ے94�i\�6[�֭i<�rcfh0U��NNqS�`g�����7����5#�_"spx���?���\�����/�۬�`��.^�8��;��F}����B>����w�z�,t[//�u�0,\��H�f%��^�h7r��q�@�lN�,S�b���#�T���x}h������)¶*Ujuc ��ғ0S�����no޼��Y�
OKN�
V�n�M���4Gv��G{	�>�Np� P5�S-��y��6�_2.����c�K��j�oC`��uY��Z�8�����ٜ�0���Z�d\L��պ�?���U��B|
�
gBk��%}�rR$�&�fp���������U;==�s������!
p�۷wNO�����(K�M4��}@�9f�Gq�_�p�_��d@6o�fE�yt(R�A:I�d��әK�<	�q���_�b���i����xmX�R�����/�bG,S��U1 ��
�莤����=(�/�c�Ծ[�G�;ݫ6<N��"/���6c���N�2x�k��/c���(�PXP�.��tx���h��gl��
�Peꉉ�r���>Y|6�ܰ��Weվx�:Xq50Xr�I���홄�E�ĉ�Jƶ	u,GDY�̻4�r�Z��!�,�y+S�����-���D��/_��2b�R؍�󳳳uuտ�����UG�jS��r9*M����PO{֮�atzz�� �1��6U%��^�Ep^�,=z���:��f
�����%`�ܸ}k�m��Nl(a��E���{�ǜo�*��{[2ڶc�_or��"����:
�ΐ��ض��T�v��z_�yUtY3Q�O�RǪ���A���֠| �^�"F���,޾v�1q�������$q&�M�Jj���
<?}��!FF;q82�5���I��L�jj���e��Ht��~��¡B�t�6Cņ����%D�w�R>�5	߼���{���������a�3�S���&�Q���,�Ǿ�1	�`�*u�D�+���{L��[��ǟ'6$G0V�Y�^T:�=K����#�Bop)%�����ؽu���:9e�_�ʥ��;�V��h:��ϟ�lѣZ��������C�ełD'c%� ��i��7��s�gdn�=3s��ټ Ѻ�.t廛[���{��˒how�����m��+���:��e�!�񙊵`��C*��c��&������1ϛ��ʺ+کVc�V8��l2~�I�c�1,Z�3�ÂeFq\e�d����x���������LlN\�W�����?�.������0���..
�V�)��f֒����7�&W�3g����� h84H�Gs8X������N�����)��R愳x{goh�t��2�!�77�u������mgѬb�&��_Πx�B1vP�Y&L�|�:t-���bYO�M��k �0C��sF�
�4���1�Fdk>	ċ��+���&��R&9/(t:�8��yc�9����k�/���3k�%��D�T��n`��Xׄ%!/�ͭk���l^�Fn4X_]yp�CLfN����|������/G�dh4߼	'���o���"�#k%\����tLn���<ukuu`���х�f�4�bc��N"��̅��2��l�s!kU�cVD&	�����6���d�݇�gysx���j�ѣG�_��P�M��04�X,/�-�l�^�Mi���j͍-�ۢ���~���������n�^�ca���K���~���m*���W��9a�ku�e}f�W�B9����Ϊ:v_
��G�xZ�>b��ꩠBel#H
B�'�>�󳳳Z��#2���?����ׯ�:]a�UK8�P�OG��T��1~UY"�E��Tm<�5�`��QY���l���z�S�ݚ����m_��_V�`�_���;C�;3��:޳B�ի۷�A���0#&ʀ�	ԏ�@p�$W2Ke>��r洲��̌�?�+�H�ԙ?�Z!����l�nQ_���c���gD�(ڞƤ`jԘ�l�6��(�eRG?MB�+����ؑ�#�K&{Jt{z�"C������,�B��)(�k׬/fG�S�*��8g�Ƣ���d�0�K6�7*s�[,
;��GJ��@_k4��8�x4��{�:�Cy� N%ʡ�C��0ð����XT{~&�V�"��4Y�
�g �`�gR�k'�4��VW�r�s�[h��4"�7T�Y:g$�%�)�l�d�ɥs��HyF�I�+d�,(�EB���!
;��=�M5	���V�㒸�wO�d�mSk�W;�4���$w����^bF*��vL������G�LaC�����%��7�|��̳��I��I�Ro�'-�./M����t����`�߭-N/�sK-ř1Z�9�x�����]�Y`�wў�Q�]sǭN�J�1�3jE��*���
�n����F*�(��� ~��5ڻ7oC�t�z��Rn��y�a��G�����?�G��>��鐥��Z��%'�t.�κ�+k�t6m_u�Ev��Js���Y���%�s?&�v�_�|.9'+�F��{y��ƭZ���[>���z��f��������r�^(�ֶ6�cOO��ϟ|�I���汿,NgW	$�Z��G�w(n����.�	�±J�j�a���|q��XA�^Ӫ���p�r�
����>�?|���4��ڝW��c%�Dd�ɿ{�N�R�����&���x�ϟ<��ڝ;�H5/+拳� �{4M�0���Tp�0���+�V�Ϲ�J������r�%ñ� 
0��$s��s�i!����+�i8g�|isc{c����,t�r�J{���kw��Jk�>�@�����Nc����J�o�Œ�Tqf0	Ps�Y��h5��E�"���Vww���8�g�l�T*��]̼K)�ӼS/3�;<���LX?�P(� 'ga}}=�hK���Ei������䪃�z�����w��{�λ,7IR,K%�"�2�4=z�*�b 7u�X�[	�nm��I�f�~�Y�m���3v4����nB6��+ƓaΫn�n����}~�����F��ET���w��J#�[�k���ѥ�)^]A��Z��\���b���R�K"
������&��?0��$q�\�װ��d��gc���V4���/�7e:�).Ѳf�7�ek�V�	��c���+�ɤP��S�]�:͈ԙ�����{�Q��6���ַط��l�ju^	񧯟L&m�[�>HL�,���	
�x��tk}�lt�#^�-TX��@���MMo\�a�Cq�&f��u�w�������z������ɓ'�B�������`���ja������9|�Z�:�Ј���7�gQ�����ۅ�ĉ����Ùs.ώAy�������s8�4W���5(�ˮ��u
��)�{�����}�Rw�ݍ©��N�gV�5�I���X�Es��kk������GW�
߰�sK�TY�b�3P��5A�HYG���UU�
�e��k5 �ڝ�wq��>���$^��M�a�`p��=�ǌ(l,�;���L�C�tNF�J���<�*}o��^��!`���a:�{�����ꫯ�66���D�nhksS<��
q��Y�d�8J�����
}~�I\���;��c�I8��Q���$eoK��XL9[;��&.ur~�"�4Q�Q |�+H_*%���:��=�
C%�>�%��hF$���2/�NY�]a9�o9K���#k%b�H�0�������l1QB�������Kj#c�.`؇��x.,��03�+dZ�����/K�̪���2�Xi��d�\SAQc:�^�x�����NX��Fl^,U9�b)]p���F�4�E`@U����w���X}}M�%"�Ė�:$Rf��R�>�0�5�XS�Pd�ܽEO�g�z�Hu0��Qh4,��4"㵅oA<�J�(H�ME�&Y��0{e�欞 ��)SR*�d\u��V,����X~��M�ў��Ux��^�ٿi��~!��fp�1�o��#�'�w���9K8�+����D	����`÷�̒�-X���Q�;ʧY�ٷf:���*7��c`��Zj������b�`���Z��]o������â�4^�f����[H�Ke18��~k�B�ϻo����c��b�nl�����Hyc4I��s`� x^zTy�B�={��t,W*,�@�@�D6�1#�gww�&�1d��4�?8�7����U����D��`b�@gj�V��m�Dt���pW�� 㰡al��7񬐍@I�kF�����͍Nw��Z�)�����?|o�ٓ�e5~d��H>>+�/���Ŵ��{��������r��r����s�wVD�(�on���}놽CvO�Vq�j�r94�/�� 7�˥i>�|i
�g�&uK5�W	��U?�/�ۗ�5#�Äc	V_��� �`�r�)rE���_�\y�z�=���$Ǎ�F j5��z��>調�y���[N�B:9Oź�e�yrth��,(�i��J��伬	LD�U�f.�oE���F�z��	�@��n߾�n
�����Xln�=���g`�!G�o@
@E��ِ�8.u�@T��3��t:I���+���k�SH���r	|�n�Z�޹&�Sqj\��Y�����x$����wo��Z���7��}�K��5�I�u��]����bW[���iՊ�8 ��Օ�(�]��{ｇ���b/P��Q*)/x~z�g�٩+-Xw#k=���ãa۟U�T>�@���5z�\<X���(	�0�������k���˼�#��j F-5�s��\9�G���,1g�p,���ֈ�G�6
�_�Ό�p���7��\�^�nmm\\��0;�%����-��~�#�W*L|�ʹ<+1��ȴ(�n�¥�5}�}�v
a�v��p2�]�#Y��`���#6(���ڃ��>&o�8-lԇq��ͷ�v��	�*�����0�C�2�)3(�[d��61r���Z��$�[<�.�I�P"M'�Ha�j�qP�:�f+��
�՝�h��xL:*�J��1�'�o3��]�ڹY��
-p$	�j~�۠u\d����R�W,@� ��j���W#���(�i�Q9��>ʼc(�}��0�8ۯ_�vo�kO��g:����d<�b����׿��\QW�z:{�x��K�Y��,d�GV/B,ɻﾋQ�	d��#�s�=N;�"[	1�3oM��L�F�4i��GH��NgX$��.�8��#������}����$-&���Ǥ�<?_][��^�2N��T� CB@3p/U ��dDB%)[���'�`��\����Ui��`KL���V�@�X�EF.�Y��UJZ���h/���4�2����2� oo��I>m+�d��1$̼(+��w3:R�t��:�3�.`f�"J�.��Fq�j�ф��4|��T��~�;Z��U�w)����ۣw}���X���)��A�El�K�!�;,5�����MÓ{�Y�ԅ�YD1z-�jq0{x�K�H���Y]]�/v�6��+�i3���A0��p��9<g�ث?P��"�S+t�3��ф����%�����/u|�T@f�9��K�:� ΋:���R|����*si�ԪU+L��Z°�)���K�Q3�6&Pֆ��R�"�r��:��+#�Z�g9�y督c�(w�,�dK͔}�D���*��Y�5����WL�+pi�3���V�!E�-�؄�a��yRKrZޒ�����x��E�y{,�?L�h80��J��n��aJ��+޼yO!�tŘ30�N�y7]�oQ:��Oӿ?�	%;�UɐD5�����r�}k�?c^,'��]�.<6�޵k��)$����f�z���#�.��4����ō7p����hNI���;�ǔowy��9�J��|�(��d�mn���\ġU���R&��\v��bl^�[%�����"|w0 DZ�넽��Ŗ�2��M�?�[pq���'�-ژ7��n���պ��&�<&���8��Fj�ӡ1R��LIH�/iUmn��ml5V�s�L�(�[[-��zҀ��r)��6�����ѱW(z�"~���V�i[Cd>d˰M#�o9sz��2���y~��l�Fë�X�;I>i���AS��a8�4�����͊b�B����sQd��^�F�-/ŉ�uר�� S�VR�'���:@�����-��߃LǊ�>d�-�++�Ԡ���due�S�ol0=��"_,D�����ë�XJ��͛�8��ۛ�����bZ�»s��%���z}NJ>��޿?9==��ʓ)=���3a�3'i��	�,b��,u��׿��WL���u2��`g:�S	j��a"�����Q�a��֭[��g���6ª�zƍ)�sn��s�J�7�b��7F������B�4�
����SsO��tEnj�4������4��[)�"�6Y�.�4v�Ȃ�A!/���"I�7a����Y�����D�ݽ{s�����_��������g/^�����
~���+(�Y�Z��9�m���k(��hZ4샸՞D�y|zf�p��ga\ȳ�;��~Ҩק�{��f��֪ǁ���M�T=?%gX�O&z:�&�e�[̇c��/R�fj��y������^�;�r�v��6����H֏N�cf!�+�ɸO���aUSX�wfI����F�?;�aF����f�Rf��K����\Dk����w�E"��7piq��"r6@wa���;~u�ŋgX����f WT�Y2.Dv3�&��Y�)������'�|̺����:~|���m���j�7��"�!�B��W�K��D8SX4Ͳ��yk���Z=|�6ыg�`_c	U0o>�X\�zV^D|eeU0$�~|�H�]�*^�Rۋf�ݾF��΢W<�e���8�*Dx��yw8ߟpuBUa�īd�f0G7�Ԫ�(A�ui��� �%�����&hf�pՒ�K��bc(rL���.x�]BI��/�wE�h�(��$��Y�B9fg9���=_G���Q��a�z~�R�-uh�[3�W���l2���*4��UQE@�SkmU��g�}v��m���+Q�}�?��s|�e@03�h�"�N�5�`�1L�﷊�9������pY�dUW��[��W-Ȳ�ײ�/A0�Ƣ�4�Ӌ�]�g|�yU�+(A�{�ȃ�L"e�]�>�0CF{��!����`�xYR�v��D�[���.?2�\<~����sT�5��vv��@��/kW��$G98x��c�J��9C���pȢr�����V=q?S�$� ?��Jݽ���P�Ze��	���o��eZ����)�QH\X_��x<�1��J']ס���'���l�����e����ߘ�Nŭ��x���Ӭ��� V�j�,§�GJ��U�Wj�˭&�20�x:8+����Ā�L��Χ���D��A�3�:�CK�����|3��;���|m�������!(y�V
�w5e�R�<�ƶ(خymE�\�5�0�^o�ܜ�8��d�z��؂L�}����v8�{6������U��x��3�{�)\��j��a��2��E��e�Z}o��-��ej�P*���x�����wX�f����vM1%�U
��7�8;�}j�{��鷸��8J�侔��y���a
~�R��������n�f\�z�P*_^���d�k���n����G�#6�u0�ILY !�+�s��������xѵWF%�[�Ҙ6�� ������M�:�������l�,I�Y���Q����Q�!���mon%i�-��5W�"�s�hH�
�{ptf��`4n_vI�R����D!�l����*��3`�ĩ��kJ0��<���V�ͦ�Q�Ѹ�����w�}w������ g�8�@�Q.;�ǋN��~�]�ץ�Uă1f)QIdՐ�O��X��mw�"Ϯ�R�d���	�v����'�PW�i 类:y����i�:9�DPm̦��r��=1L�3��%��jk�D��?�?[h�����;�"�������Fktq~~mw�у��}�;�y-*۴��Π��)A7�  ��IDAT�i8E��h'�P�^�;:92�<aS��V�q��N���+��`*�/�����"����"�	Ma�����ӹ�e�nD�%B^��n5�ʄ'q�s�F!(Fa엊n����������2<���썭���M�7-�
���7;���+�7���|K�9��$8,2de���l��zp5�����"l��ԳR�83=���|Pq�X�C�L3���q�������X��:���.T;K�r;���u�~���狂�[��R2娪����1R�.�	�C�������Ľ�dwv�l����|Uw�v��p�䌖���V�/���u?0�]�Hq�`�p�����+�}vϹ'+�jW�L����򙟹��s�	y��?e����,����$�M�S�e����V�m��V-��c�d�0�l�J����;{b�T����X�l1���ȍ�Ȣ"�ja|(3:�6��(l��"?�,P�~!�Ks��uB����,Ĺ{�~��吔�)��y,'C���9P���`:��X���53�K���ʀ��z#N�_z*�h0M�r��EO��|Ae��%w:�3"o`Ӽ����]E��I�D��I�j������Q��qB���i������_A�%ϯI��T��
Ad���������Hs��Ui�4{�z�z�2p �iB�"�j4�0�y�V͎�.zZ�=Lf7�����/�������K-`�={v�Νu�H���&J������Xʢa@��o��=��w�o�@�:�E��`�佉�)�Ȼ"���ܕ=a����r��՜�0��-æ|�u&\-��2Y�W�8��*բU�u��e(����YNKzź���pc]y�,?��^<y�~Ұz�(���>�d��B���ǳi�hs���[y��DmL��w��$�5��Ǐ;y�N��{�>�e���V��Q�aE��ic��R���g3�n�*�UǤ�J,N�z�d���Մ?����Ҩx.�m;k4��3�e�b݅)�R�SJ"B2���b�amw��Sf�ZQ/�c�F�K��~!F8�r��8]�g|���f�Bs.S11��jB�Ѩ��͕]����S���T�L����z�J�1���0��z��L�{���Zk&�I]�&nnzlT#^����IY����,���r��`z�"��w k���?�����	L�����n�;,sc'�@��lN�m�%�
'�d<!ǭ�z�W䀫��*��&�[�z��:Yjް��R�Z������di������bN<�F�,>��b��ٲ^kFX��C2��[����V*���g���T�;x���1Џ8��s�Mf�4[έs�A�^_�"{�A�]�:$~�^)��шlQ�ɴX�z��V�3ƚ����S?�p���F�^K��<��J�
�Vl3|�0���t��m;�ϰ�9ԇEا���ѲE*����vXL\RK/˯�Ou��r��Z�*�a���򽾢���t�>��ئx6�%ßP���>Ѡ/��%��p2&��l����"���n7 3C����/,�%��k���'o��8F�r��a8�8����ܮ�(���ɞ� �o�)��\��ݹ�r���Y?��h�������J�$���.�7 \"#�X2؈%�k�l��`��g�� (�V	�5	�^�d�x��-��Lkf*�T�^��>Z�'O���\�ķ�Y�t�e���J�Nʁ�-Wj����Ɔ �:�f����玣�b�>x�d�t9)���o߃�;99YL�{��Y����,o�ެ@�ΓY���F�h��"�ژ���&��4�f3�r�1/���l�6�|���7���EW+]����j�߽�[c�M�o;�%���Y�Ge� �ą,!��;＃KAN��N�_Q�d�V�����������0��:QkbV˵yJ�yf�Z{S֓E����Ը�0�y���E٭*���_�)�ZS�x\ ���g�}6[PP*n.Z4�xE���ru�~	�-�1{*8�/�5�dkg�� 3"~����}�]7��;f���,���τK`�M�@����?����ll����K���]"UY��0�����3�2UEcbF��M�aY̍��g�v�蹦�
tK2Q`�0�P=�k�
�!���ߖu�%�&��2��Z5��f� �10��^c�tc�ydk�ܸb��}���HQ&`��
�=������CIb����;v�C��R�L�V��FjD!"��q�8r{w��4Y`�[�O4/�v>�� �&`��u�_������9��G��"$xd=Np��w:��99�Z>��� �>��S8���������	��R</���c�L�JUp�o���4
�d�B��-	��n���-'>�R�3���G�>|3����mv�b�h��P���tY`\!wٳL	>o�X�14�Pu�vWMDLQp���c�O.�?�S��*Q�:j�f�Gᵿ�2xap����<�кJ�|�iө�9�1�svU�N���ޠ�`�i?>}�������	�h��r��FI秣�����6$���Qɱ������b_}���B!Ʊ��$�&6�{�f���^����1%N����LC+������ַ�o��b-��٬[�ׂu�&��g�0�
�f�Xz�����P)8!�1|(�cp�&ҽ%��ڜʊG�����M��ob�D^��Z�f���=������l�Un푇þ�%|�V�p������Ws��YP8����z����[��}Ϡά�~�i�X�CZ�G��������Γ8�Ÿ���M�R=y�27�B��b2]��27I�R�������-�ۻ��Ԛ�U	>������W����gD��#�&��ь�)*:���*Xh����a�OԖ�R�]�������M�PM�Y�ަ�5���^��+E��б
��K�l�+�n�cV44�_IXX���&�"��$-��Z��ma̬�����x�-\j1,����T��($c>���{V�yA�Il�p<$L���˿��V�������	"�Ԩ=U9�R��m���ˡ[8�zC�gV�t.�D1�i!����N<wU��KL�y���Y`t�lts���{�ޙ����������[0/v�08P!��Y�,�i%
��S8E`M���c"���2^x�ˋkM�*�Y�<�o��v_@u��*b/����]� �h�P�z�ίX�|���eu|lb�a��.�)��V�*�(��H�hY�N�_��$��9�ۊ���4��R4WV)�{�w��ū�-�Zq\�Z���`:m�۰C!��a8����*�|*��l��r��3oc w�յ��/�r��y�$fl��Ćd���� \��l
QC3����L�K�����X�qs�gNwc�l2���'����G�������;IF/���*6��������ug�DKo8&�[ ����p7��Y�7.1�ToWD�C��Gou7�$�mԫ�{��n�(�qp֡zy9]�c�Q������&�-�88YN!NGT��ق�T�[o���ٳ���a�\��R�Q�cJp0��H�y٪�������Zx ��R��zf-^���H�](�DF��ÿ�!���-�Khʾ���Og���3֎.("%�eYK��j�r�L�|if��LxD+ ���눳��_���Ƶ��XZ�ek,/�}��<X�F^�=�2�k'T�	^�ZVy �y��r��캀Kw�
�r�$N� �
8�H4���<	�<Š�͕��/ܗ\I9d��ʅ�QL_�`��v.�F�dx��`.���?(�$�灞�L-S^3�z]���0�C�u�0�Y[��7�W�Ȫ����{�=Q����*�>��e�ے"�B���<[[���9��#(��!e����)����jًm������t�՗�%���K�$�]�`A�ݩx���1"=���n�1�%����[mBQ|��Eς������2w`�'fV|;f�ɁeA|�.f��B�si�����7���amX��^�������o�zV�X�[0(J!%+3jF�shAa��s��v�QNB���c7�
�P�>x�@��5r�
�Ȕ:�-�:�k���-T)帬�'�j��IU�((c6��Թ�h�z����ky�Q����ݽ��"�GMoPa8�E%�m�Pm�RSn7n�#����c�!�	KI��%����Dƫ�����U^H7�0,��nZ���{U�8��'�����a]�`����	��O`�-��$ax��N�sp+{;$؀�Ma���p�a<j����ރ�ʕ:[�_Z���wU�M��������_2`��E^�VU\����˽ÃÝ���&�QT�n8U�-Y7fL��]������ؠ��-�����$X��Ft�۝9Kp*�WU�zX����ǟy��n�GC+F��T/?b��&9.����d��4;ݮ�W
A�+�_vKa>6&c��(�D4��X�ԗ���)A�f���8���|��qjX�)���ә��5K����>5h�_m�B�\V�t��b�z�#��ؾ���nMg�$�5��Ep�`��?}F�\�����t7�ї�_��O�����<�V��*y�� �D�o�as�*�Je2�{nZoT��t8��U��b-�'PX��Cgs�7�5d:�.�e�޽O`4�Qޮl�H����D�s��Tk�Z�B8�O� ����gF-��8��"wGÉ�h)ߣ�ćM�˒����pDgj�)l����kU���fW$+"a�[�y9X�Y��p�a��򈍫X�ᆔ�y�K��]N�5��U�~M�����۰p+���/����o���;�pC���N�G����\��*YZh��MO7)��;0��BX8�����#�:�.��".e�J�zh��*�'��MIZ`I/�Y�Ҩ9���f�����)�t�W_>}���Z�W�����7�K�ԍ���-��,��;�����B=�B�����;��]�_t�����o�cj�
 e��g	F�/����a}bF��N�m1XJ�V��s��W��[`�E��wCN�;{�>|���U� ��G�H�7E8�X��a,�ZSؑ�;ݒ�	 aVgHc����)���.3^�ޑ�8jj�������O��xu|�>��TL�v�OnÝ��1���Lq�����m�&�����Oz|50�D�g)����X!����`)3�1���q�1LԊ	�K\�4�B(�ɶ7�O�=52"h*�d����^�t��GS��X���\�2������Z�Kwg<%��i�)*?b�kK�A�;�K�,�D3���+�&�*���&i�X�g���7�'oUX���xzNFY��ι�8ae1�6�aT�S��Ԙ���祽p�O>�7���#�{P�⬆s��{����y�V�H3J����UFi��9�QEk^^�c��Z���3����b]�-?�˿����tgg�`)��$�>fgh�90�J�I�Jaȧj8��0��7�%k@b��S|� �E,[Ƹ*�&�u���*o<uM��hS�3�.��>�jy��a`�nmp�m�,y����S1�u�<����]ȱpo��ֻ
��B�
;:�{z�k%��0xoՊF�`��D�.y���S<�q����,�Fj�`��%�,�]eX	N53(lF"P���4��=L|�A��$3�%��\�-F9�ʊf��B�r��/qۿ��/I�/xf��˽(�?2�$�v�1R�=����͙%c*r�Ր^½��x��dHN��Q���K���T����sٟ��^� 3c[�t��4%��:J��s����ѡ������nn����`����-��#���I��|�;��FW��i����M���/��rwo���_��!�g��8ION��i�� ��r�]�z����m�?���?�|�:��̳*1���ATb{Ψ�{�����a��~�=���W6�l������Y�fj�_3�0��c]��:d�d7
o���hj-����R(��ɴ��6[��$���.���k�:�8����e'ɗi6��i1���nwK���B�a1�
�T������/hْ/R�жO;fK�f��������i����X�9eh4���shJ��;�Ñ�2V��KM�����9�����a�bi�a0�i�wqu�J�0"ݎ�~X�566�2u}�y|B�-ª���/~)�KbkR�B���R�$��G�O����$�,M�l�м�>�����I��TR����_*���\�$�mCc��:P-���>㊡��c2���݁}xt����E�X�.��+�>s�5kᱛd)\�x<�+�d4�X�	�[Z��n�+)!��ˌh-��Wy���ڜ�a�kCA0�ek%���a�1i����������Bm(cK��J�,�SzˢQ�a�_�W�fx��d4=�V[\YTl�w�ְ�E?�h��e=���j��X+`��a��<R�̅f�u3��p���sj�Zv��U�ݽ��{��N�m	Q˧���R�ȱ<������E���G[�|sgS6x���@��_�.nn��|Ng�<z��~��A��g��9���/8Ԯ�G�Oj)'�����ZX��i���0r������vy�wu�޽$N^�|iQjv��VU������Y��V�vDj>�m��q�-�"r_���M�8�����	���ŦS�L����0�r��d]��������;�����*�������%N��$��5���=T!���ɏ�ސq���'`JʕPä�˗_� u��F�������m��(�.¯��z4�c��߈J��V1G���y$�H�j�F�,�aI��꜕6P�@�rrX���IB|�ܓ5�� ZamyX�W� �i�Hd!D1l=�\��s���2(��\u�jޱ���ּb�glV�R��ٍ������Ex�T�z+��Z� �nkK�&������n*��B�d���>e�#�O��OO�?SD�We����~�C!�uf/�j�6j:�Aq�*�����x�����7��J����)�� c���f,�Ǐ��і���!�{C��2|d�����Z�m��tE6�"�3 �Y��fU�Gc���R.�Y�~�)�#��S�z�-�Ðfܰ�J愛46��PX��TgPk�m�GR�,9�s�Ν|�ʞGw���}Y5�-䕯�$�bg��I_�ҟPi��f�~��Y�=�om4f�j�1&@a~�{���
7�1��S@�S��E������h�e)<�1�Y��?J{�KQȈo�j��c�XȒ=8{��~�����6���֕�;��70�za��|�▊J��#�2rP�aU`a���)#��~��4#�8�D�^�^�>��ܭ�����\�
�L��c�M3�q�95�&7,F�1%5�C
���z)�����'�Yއ2ϊ�嗿b���pogwǯߜ�����#a�xQP�7�sb�n���By��Η��5��̄g1ŇW*�*�>�������ܭ���}r����{
�b6���������.�)<�������[� g}�R)��g��ux��7�zo.�[�����N^���%��nlo���������v�E�׳����{;[��FRDI�F���̀X�݃J)/.`̖yi����e�i┊����ژ��aG�����B�Lqk�Z�2Z����/�,ƨp��U�l�-��	�	��kKω]'.�y�TL�$.�lR�V��m&]'3�(���,��<��Zj�g�vn�ga���������W�8O���/��s����L'0?�xaa1m2_�i��1��a�2�n��;�����O>��k��+VS�-�-��������.7�tX��W`}�z{w�|M��|�5�!Jᠿ�M'�����c�=��^_\��xoYy ��A�PDa1�͐��(,�IitӬGE����R��.4	�D�ܻst||�����Ofy���ꞿ9eEq�lg{[:���=��E��'�^\��;do+��p�H��s��c��?|r��ڴ�	����驝��S�~���ǽ7�ru6$	M�L������N���C=E~�ւn��-"�,��77E9\�1\�E����z7��̇������vD�3*g��ky��A6��"�t�0��+�!oÃ��$K���y�,nV⤘���s�퍇g����<��t�s~v�ֽ#�,�R���ݟ|���[�6�5��倠�f�q���ؒPH��5����FI�@�����r�5Dg����g���S&�����)Dd��p<�ū�W�7U�)�`2��8e�����M�{�g��ɢ��F�9q9$�Q#�ü�����g���`��_d>�����p׵̔x�B�bU��W�U�t�ъ�|@gz�νR��Y��nGކ�g_}ۻ�G%�{Y���?0���ax�ՠ��O���ۄ�����h:�F�ޛ�҇P���_|�o���E��X6��bZQ��h�8����O������M+O��;�6}�R��on�<��Xo�(����BE�LzT�8!�4,�������-h雳ZL�'�&xw�(�,Y$�[���d�����H�%�q�:�u����D�Ep{ꥡ�a8��M�۲h�la�)�y����Y�I��(�<s�K�Fj�$�!��6�R(��q�a�h�X�����d�E�U��;)W;��o̦��ǔ����ۣ�8�/U]![��Y�^�ྼ��ɚ�����$�\^	IE��[c��I�7�Oٛ�-�S�̾hk��Nbf}���B�Cl�f��߿��Ê?1�f�7M�;VL�W����|5��b���O�TRքqň���2v�T�nc	H��T��4��(�U-���ׄ?�]����r�`_���k��� �F�����X?��3F��W�lR �uV?���u��}+�H�ş�0��Љ���V���6R��^�����T�4�J>���M�����˜�}g�+;�Z�[��T�fz-�BU�k�������+8#ͭ�j�Q�i����O�����|��������'��d\�LZd��Hs�)1�k�X��*pϺE�����Ƨ�����$O�ʠ��%�A�hTz�x���`��*Z�"*�)��.
VH����_��M�'c�4�����^�x) ���	$�w3`��4�3�}��gW�
K���k:a&u:%����c�O�W�U���d׆ry9c�IPﯿ������ �je�C�:)��<��)�I=�?����Ç��/������r�a���w��H:�KBT���g2�AE%�U4���8�=y����ѽf�cs�z��+Ώ����JƪJ�B�� �X�0���Ĵ|��)�l�eq��X�#�LKY3���!,��\5l���*��Z-K���j�rpľ7��p����i�$�����x�J3�%�ጵoqqs}��ݭj�i1�R�����gRi�+���h�"Ҩ0�IZZ�M�|:��g���|�T׬K7�V[U�x��Be�m��(�f�"}��g+F��E�wX]�#\Ż����&m���q=y�>x�@��>5c\l�� ��>=}c}\�.[5;��<42G��J�:�Τ��I:�/����!���b�X���8f2����rS�t`-XX���)�&s������i�|��Ǹ����w[��z��2��x��V��M�ҌS���4w
�I�_^uh��^�E����������3C^��9�}���$�1V���Jը
ugg�\b'�����d���C����\'C�
�s�Ю��j���8��$
�ba����asG�FE�	.>�-Z���~�rP�d�:���t~��%�a�aU�s���`o�g�|��BH|β����z�@�����b��VȍZ�:[,�HD;����p��2(��x�C+:����ŕ�&�'/�����yl|g�Uwkw��zK���l��`���Jq�f��.��aY#�T:��%׻{p?�<�r�P0ö�P!��)�~���f�%�?C��R�`s��@�Q��1�d��ܫj�  �~�mI	��X 04�e�]J\`����ao<����*��.i�A��2�Ft�UL��pt�>.���B���B��.�)��*g�I�i2d����|����Ĩ�u��|���*�4l9�LUk)��a���~O]�N���N2YP0��{Al釒Xׁ����|���h8�]
�����:�{�)��fc�OUj 1�<�
qqp\d�;�0���vp�;��OF��oX<W��cvZߖD/|��[ 3���2�o�%����:T�<s2�Q�X�>��k�XWA+��X�!,b<v���D@lE"�N��*1��cj%E�KkUMb�g�������ʍ��@<%f�845�)C[$s�?�{��*[��Ш8�� 3�Rf4w��*������4��|o�����Խ<�qD$���O���������K�ᶱUu���u%��[�Y6q{��$�����W��E�RSO�ERe��=p��؊�*�L .l=,���0��V��H��
�%ū� ���E�4rU׌^:Z�%����TwskN�H�Ƹ<q|��*�+�dAXi�d�Ŋl��ys.��J^����l���B�ZӮKu���r�'�Qi��y��ۧO���&ƿ����\)[��N��)��ɓ0�.60Q˨S/�(�4Nؚ�4;�z���~���%����+(!rOXk����'_�k��D�&�H����8��0�T��o�3L��fӊ���?ll2�[)�\�t��-�:�\Tq�Gw7��<>gXcB�;�Z)��l;�5�p��ӢPy�\u�?��;���.��oTkp;0,���|���&���v�x�����2�F���������-7���=Ձ�]^U���N��,WZ�~q�o6��ۭ"7��qgs����x�^�Nu��lg,0د���͈��������O�jӻqqz��s8�n��Ȅiʚlk��[���Y�f�������%)1���T3	Z�	Y#�ؘY��R�����r.#憷�]Z���b�)y&�A�4c��^e��A�D�%��ı�iY�|�������Bبخp��1`�a�����P��~�ũ����)s<"�Y���d44���`��{��r�J�6�I)�s� �5�PV$�������r�����O�ꫯhAWk��N	�A: ���J�T�M����5�;d-e}R�֛��Ś��eO�����/�{Ꭲʪ���!5_Bf��ȣ��+⿭m��g�a��#Z?�.�@��f3C2s(��u�EH;��7�&/R#�a���'C,���Ūт��CYO��pU��}�4J���h�#��D�K�UN5���k�^���r��B#i�������0Lk/��0��A�O��q�8��X�6_���T0\����~�F�o<��A�,Ў4��ڧ+���5\�R�X]9�{Wu�%�OhX�rt`����?����騽4��+�<�-��in��h�[!޶5�>c���.��CZ-�iKA�^�\	\{d��NS�]��#|**�$��լ�a.�A{T`��(@��*�f+oS|�t�.��$����c6���F��ƿX��~X��߇%�?5�o�W�,	�-77�1�Uf 7�l&}Xt?�7���>��Z��V�OM����h2��c�+��>���S�8�J�0O0��D�h���*`$J��v�d�R�a_��\Y$�T��8�&�٭���&
)n`�0��Y�L���0Ξ�V�Ҩc.��$���?3�l�����֚Z<7�V7UBo0׎9Iؿx�ݎ$�b�� ^`(�P�Q*��0BL��1>��`�O?�YD�&b�t���H������!A���8�j��4���T�.��[��y�d[�݆>�`�C�2EԨ�����FFRhPx{��X<(���\4[�`�0�έy��]��7�>�裏��qf5���'��;)ۡ�v�S�ӭ��kc�!���&	��7�-�nJ�DEh��jC@�Y����1��ݺ���z.�3:�Y�2g'�Q��my~��> 7��A��[��e�F*4��wE�����l����̜Am(id��9�ɴ�F��WvG�p<���d���9{c���o�sL[Ψo�R���s��^�jn�"� �	ge~�\��ؒ�K�e�A�c�����	a�J���f.�A_�%��$MT&��SQٓ*�rΎ��D�f	���[
�BRI�H2(ދ?�W��*�TnԹ2J��VX^!���;b�@�lhVy�%S�pg�6��Ӏ}V#W��-G��~��EXǯ��-2N���
��O��{�����Ә���g��5=/�h5����J,i��"����lio\�Wa�{��l>���ƘB�`X��Gxӻ�\�kN��kp'��̅H���{x�.}������ʬ��>�O��p��܎�|sc��
�����U�p�����a �<9b�d%<�ׯ�ă�7Y{8s�8r2��>y��l7������t�����
jIH�w�ш��:8� �*T-K�2g=�c(C�%#o���x�-OEh@�:��]�	k=Vp�+��&�A�5�x����_య�<U�$���C�����h�!�,Zu��`�k�S�������er����c1���fY�XR0r���{{ga1Of�Z�qaPZ[x#�}��<��U-u:�f��Ժj�q?;�$��; �V@�묚oΠƢ�F���Y�f/~FT���C����Sm���^%0G�YT��2�ro@������j�Y/�d�u����'��p�oo��dĚ
 +:�NB�D(��(�6jui�2���Œ�k̂*q�ضx�٨��S)��������j��9l�$�����N\�V�6Ⰹ��]G���`g{�L�D�5�l:=y�z8���c���M���x�80Vv+�@0"�N����|����U���(&G+�����Uӕ1d���l6�.���&K��7�Ju���������x	hxM���VΔ4E����>c.j���֖=ڡ�3��nA���}y���̚ɭIP�M���
���ä\N������x6ف��=�J��%]���#"u���咂�����)�znj�.���LI�b �
��}s�[�_â�����b7��.ȥ6T�1��p�V1ԍ󣽾���Bz@$����Ϗ�cwww�P�Gj�x)��3�t.�QͿH	g%�Q���`\E:*0��'](�4���o���� �٬Z�(��"���}��%�ˇ{lu9\�|D),�-G7Y�ꚕ)�x��>fdf`��3Qe+v|��ɨ63�f��ߜ���R Yqژ���������56o�J�c+���O�Kq�_��W��9d=��ĺ�u
�a�-̈́T� ?7s�P�fACJB�'�?�|��-��������G�1Q�a��1u��`]R�����9��_�h��(d��|�td��S�q+	K�W�*&��V�x�o�����@��5����|�#����� Q�7[��d�n��VM�_��v5�jMt�J_�%�-�m�����<9���A?�Oqm|+>1�f�N���Q6[	�
|���6�t6��`b��J�>@�:j�l�g��s��IVL`�e�*s�ʘL�1�n�?�h��a@���UA�83���U�k�5w2V�K&�I lBOXE�ݻ8�?�^WM��ٟe�����6��,�����-]�y��|U����fz�(�q�b�r*��7Y?�*�7{avv��4����5�y{O*�ӣG�D�e�C���:Fe���'@$��:����3�8�H���ʩpF&�>־Ewk����gϱ1&�4g<��~���;&@hƒ�8mGX�W����~s~\�"x�_�T�IJ��v�y}q���_a�������@�]�K�wߟL�b�nt��x��� �i�����t��Zk�)�&Xk�*y޲����3�C�����) 7���0U''��j�k���(IoN	L��L`x���e�?���n1LA�&�S[�`�j���W_}�ч2nnX�.����AY���P��-�޸�bVؽzͪ~�	2	���$�b�(����r!:JՐ��zy9�C70���ذ�&�W���tzZY���p�Ԓ�`��!�֐(�
���m���rD>�6)�Oha�t���)��JT��ߕ9���t���ǁ����q,F��ٳ�-D�#�
@��"��w7�*話e:#�0��I�>�y��N�aV�R��Nu�x���&�	���ZE��&��G����s<�_��_?x���O?��m7Z�ǏWj�h�3?�Q�y�ˮ��J�[*��2\:ù���Sp�CvK~��I�g��ܨ�U��E#��y�p{4K���`�[�pƫn?�J%���1��l���������L����y��J���ƲWTCj@�T	6�6ިc��>}�%���C�v~�Ɠ!���p$͇�Ż������*JC[a�h[�T���y���2;�9���C�A�����S����}��O���sU� ���+��}�\~�$��=�_ߜ�>���	ŁL��gJ:r?:EFy�x�7��`f�&��4fC��;��{D�Ua�O�<��3�~�?����P8:]�[Z$�m���'���?��%�y-�&v�t[J�|U!^���x�E}I���R��>iks�e�.m�N�f�6��KZ�r����?=��+������ �1��d��;�eqA����L����8>?�N�9�k,��B:���pL��\��,����T�!>\�T��Bվ�)�,$�Onּ�TsK�J�7v6���Ͽ���w�j[;�N������s�ܶ�5
��|��I�UcWƈ��wu� ��`�	�SFj��X���(�[Dm�����N#��?CaV���bR�`�}���]|� �Ý;w�pe��$���v66X�&�i���/�|�wľLdpB�f{{K��L�����H���K��2fd\^�Gￋ#q-M��.����s�w��A�<`��h��q�P��P�H�J���9ys�`4�jYF+�SBA�&��Ypi�'�M�w-6T� #ZA�$f?�SV�rΔ��&/��d�q��
-Pɚ�U���8�m��T�	B��P�&8cr��Ej�K(Z3�F����������k��W�t��_���BW$�jP2B֎�����m���[���1D<F���CW�$bW|>3�
�?�N����):2�)�U��KT*�!��K�5�5QIXXx���&�2N%������bTnnш���HLIa8�Z�9L��.	<�Dm��hh}0kUv;�r�0"�j1��j���x��s���s6���k����?gFh��a�܍໺�Ws������R���14����x�h���v\`��7o�8��[��~�j���gwi�P�}��ԝ�0�KܱgW��P[ۇ�fC&R�])n_���jC9��4
Ň�M�C�c4�?}ƪ��6�<�܊b��T�����":�c�r1_��M��mm�Q�7`���`p�p����Χ�4˹�lH����t��Y�Oa!3�D���S�=P��J5*��S�url�"�+U��E���
�[����Hq�gW7�0��%r�dɕ�;�.h�E��B�2�'�L�ĎR2+r�1�h�;m�Ź�2���	s�����-|���աO�|��?4|lp���!Y��e���P�׌�`{��	�]�!������7of�a�Q{K��CI�7ҩx�/N��T3p-��x:���@�H�t�\�gg�}%3$��8�O�l��st����U�P�EU��,�|w{n��5��ׄ���FӘ4��G������	T���1Z����ۿ{�a^{�L���M,���=�#Ɠ��!�D.5�l!�	�d�3��,ϓ�*�V`��*U*w<׌�^j�(�X�&:g����A�f�p/-bN��|�]�_�-<Ã��z�����X&�F��&��f1�O0��~�°�j#�vg������k�+����	)CVG�M1��1�b~�MB�g���G�kM�͖���9��>�������
ǿ9=a k����>G�ݽT��uZ-60r��1�T���0���(�����wn����q�t;�	��0*a����{�0�O�V�#��9K(�kϬ�F�;�����Rn|�m��ՈW�x{�خtW�<V!�a���Б1�%��I��ɮd�A�?�h���ݿ���q������$�{��a.E��f�Lƚr�+�h|M1��#���/�r�"<�o~�h�b���S����X�x@�ZL�o\��z�`�(�����3R�	^����
Wn&���Bڔ����Q�O�g��Z8�܂�y��n;�M�veP0�8�𜄯�{��]"	���1AC�Ψ ��Q�L	=���^J���[E9t����c�{�.�ꇊ���$ѷ%҅��VԘ
��d��5���=*�Ƒ/_���*�r��/����WWW7�������B����x<�:��H������M���믯�.���l߽{�"+uT��1�CHY�����F�H��P��ȸg�L�u��_�z*A�I��~E�������Qej;!��F�慲�ɂf��5q��d���Zx�TxPŸҭLl��ʻ����+��M+��4�6�����k�ia|7��r��� ���;n�Ĭ��G�F$s�-Y��|{Ji3��6�L�<�� ������zֆ�e��VPW�]Q^�r�8[�f*�WS�U�-�B�bGb	�I�U= ��ٓgg��jn��0s-H]�r"+���y�*91=70⃁!��V��%v	|����j3	]�*��3v�KyZ835�PA�#�ɱFR�|�8ŢC��.ZL�J�nSL	L�Xtg��+��k`�2�/.����}��Ջgla8���lɅ�[N�i�j���c,v6�̌P6���_��.	|�4Ɛ�������x����|4
�J������U8��8q<>��o�������0�8�|:��2��&�JTn���06aߍ�AzYB [�N��`�&�.��d0����{;�{i��k����Qp������rT�37O`���J����N��޽�����6�v�m8�z�
N��˱�b�g�Lx�h��T`4RW�y���-Bq�TU>�s��f1ncM7G�T�X �3���ݼ<��qp:T�q��}ѧ�����g��*�h�W�^`Q�;�:�q�c��Z��6|/v>�ӛ�K&�˕O?��7���byyAR�r�4�� ²�Z� )�;��W���[��honNNO���r�n�Ռ����溴�U����{��F��3*G�������e�n�0��
��	��|J���b�#L�����nˀ���&��t0Rl<�a�&�J:==�#����QE -���-6��	�VҾ�!g(�=��5q�2�g+�j5#Z⮰�הj�LY���$���[�Jk ���¡1C�%e���9�-������v�e,�S%x(�N�5؆S)�Ǡ_5�l�ƣ��O���x��1�P�IƹȰF����ȶ77k�����J�X;����a���Ǫz�J}����A�����BǨ+D3��ѣ��j�)j|�j�X�k,��זg��=K�,��V��z���`�������z����x��:�ޤ9�D?+�Nw+(U��<�-t��e�Mݦ��5�V��y���r-���`H}�ͩ�f� bǪ��x���t�s>V+W���p��&��uXL�[�1�%m�Q�`5ұ�u<�q>�[~��_�k�X>M0������ܸ,Ȥ���[o�C�!$˴�8>>�{�Ĥ�%�����;>�3�~`7FD.A���rl)��Q`T�<�fٺ����.Z���WO��'sa�9�ݶ�7��{-@�ѦK����~�� �"�j6��˞Y��r���=R��>�F΃7x��|}3_�V�:J��U��j$�.��+8�
7 GV�^zK��gǢ(^�X�Q����ꯠ��H�	���QglY6��![^|d���N�m���Fc�
�&d]�:�|��[���6{iD!��5*V2.!�-}�RY�ټ������Cl)rpۏ��5%n�7i1��x�s�h���{v�����aa���C����6��@��a@`�A�c@x~�l�Ē�x1���v��bB�=c?���,d�yh1)��p3����L2�]3T�����9w�Ma���+%��� 5������0*KUh-�jF4kd��~���������3�b���t�&�	�T7S�J%B'&Sv{�(}��7[�{�(T����%o�_���ݎ��gƶ���q1�ȕ�W�����CL����۞���X����:;�����e���g<�L�b�̆�`u���>�����J�";�:A�+��?JڑT�
�	��9�
N���Uv� ��N��!)�ETi�*�v����(=HZ�S��2�pGD!/����/�z����۟/�Ó������0�� ��тU��������T�sX�g��P�+Vڰ|������tT!����z�v��IB��2����?|���
y��uF��JIܖ��C�����!���E�L9�Y��?�	+�R�c���fg��L�~Ud����&��j|�7	��(�0/�ǯ�>ɳ7ǯ�|��V7����:W�9,i���z��>7���2��q�\�[�"r�t��ʝۼ�+u���^K���B�IRz4� �uK�'�)I���6�x�Ν���wD�=��7~��e��d��~2����>��C��X�WW����=a������l:N(���pR8gE����ʴ�ԟY�-�Y���5�h��L�x�
i����'+0���EJůR�@��XGPy
�Z�cQ��5}Tzx�A�Ε�]$p��v,����5�X��&�rT�����mACL�i��0JɊ��So���XK+Vx�-�"|C��Õ�CT&ܵ��+��{�d��ݹ�7���#Ny�w����IGbX&l�hbU����3��[M�D���]��4z��Ç�����:N�7����.�A��|s�Lw7Wם�fw��٨כ:,.-�\J�%�+��c9?}�Jiplr�e �����e��[8ߋʺ?,���,��؏�/��4��c����7�L�����r7��S	-,;��N����GoNN�����"���Cl��s�����1JӬV1��$_�r	�a��<��Y��	��Fw^X��̶G��)��ͳH*R��zlQ��Tk�y�Vg�r
f�3���s+�e�.ـk��O�ސ���]���)L�2Ku��u�x(l �
I:LO渖W n�ŋg�a�E�dO&BM���X��X��Ui��c��Ԫfvt��!~����ۯ���f��k� �9�F�:�7���*pۿ��op�}���ֆb�8ۖ�vX��2��#�#Qm�̜�⩫X�1ʌ�ǳ��X�Z��}P��TB��:��:'ާjg*���,�ovI�:�+D��e�����^�L~%gY�ïNO��3��V7u���K���,�\g��	��[X�*����b�U��*0bCQUTP2�ӧQAq�'���Q@~�l�2�a��k��������;lu7p-�0[��%�3�Ȯhϟ�f�]*F���תׄa��.�r����7eEq�6�l�d�^�,يr�k����]ڮB��:[�V��=�X��:k���
����X,��Ŋ���Ѩn����՚����F[�����	���o� �Q�M3L,}�R�ϋ	���[M�;g���f���N�*��9����F�#jj��2��U鱟Ž{�J����1t�匹|��̅��[��cю3�J��H�`n��1aJb\ƌL@��K�C��J��:0P��<}sB��[����������Or�A�W�w4�Bs�Frg0ga��/޼n67,*�lmm4"h�n�'�l��/_C���:�(-Hr5��A%�M�J���9d_�'O-��˫f��9[.��G�
	���F�U�j��"M`�����딜��?��5oP�"��C�a�/��!��_�v�r���g�䘌X1��ϖ���(ْ}�6���/ǃ~�ќ�'�)k�*�;�i�(�iJA��G�d�ľJe?z��D��-
ZS�8\���������D^w7ۓ�T�KݨT��t���R���,�C�v�ӣ��R~5��l�w6'���5{�n�6���ln��L�&Dkx�oȧא�� �N�Ћ���������E�V�'3�pR8�X���(j��l<��gWX�u_^�F%�Z)�k�f������W_M�ݪ�g%�������3%���-�b2'���s�;��,_$�^��7����۫���{�YvӛVkQOV�͍.��7���sl��F�)�8_Lg�`�/�3��R��?1�K��٨V�,��Y���)x�A��Y�D:Kσ��=��F�D7����V�suv
'e��]��YJ������޻w��q�Ѹ����o���i����_M��"�d�^L�t�m���St_f�Jp���t1���a���$�-�8r�b�����&�Y\���T��^)O�,���z%�͝"��نqJf��(c¬�Q���n+˗0�hF�Ng�`@b��]ur\c�IR�埰"�e*�a�9¢:�A5jz~R�c��[��ٕ�V�M�r3/�~ᄞ�V����B������,7�*��ã��6m�A�/��f�	� (M�z�u���e�nln�x�՗���[ul��b���a�c`�NZ�t���f�/q�5=��'�w�4s�:��&+jt+�wYW�����~��2(��8��=��R"�H�Xi�P����%w��(�	����������U���O����U�~Zҿb��6�dI�R��y��7������j�n;\=?n�>���<��aRܒ�(�ه�E����R����Ƅa�:#�E:VE4ݷ�=���(�U�iS������[�)�nՂ�g�9C�Y�O���yͪ���R�,5�,Uļ�Z+����,��C�}fLcЛ����K�2�׻�d��q��m�u/Wd��!�0g�S��!>��"�U7pn/|us�떼���TQ��.U��+v�`�q��3o�I��I�TW�裏8G���_�-&w�.r&����o�8'�w���3*+=~sJ(g���|ŃK.��(�ܳ��[�#Z���
��Vm�sM��8)����3�=y��Z�����qE��'oL������y�O~�L�֕�B�;f+"�hY*#Ku&o���`�}!�ԏZ�M�+͈{�u�74�9�.
ٯ�؃�h%���4��|�#�~�#�j����]^@�
A(�#�B9�G�ᄐ�2��"���U5��Ŭ�m2�2S�G5�+H�ό�l���2f�`��SD�1G<�JJk��Jr����ŭ
q,���(;���G���+��ǯI���5��A�M�؃yr���J��`���$C"Am����U�D��a�*q��h����T�MXHb��c��P%��]����f��;�5� ��i� t~������gN�z��7�����-f\�arficRS<��R�O� '"�Z�JS��l^2$[�;�df���_������]�kTo��<,%^��dZ�Z�ݭt��ƓF��s���tv��;�
E���?�x�=�q�ᵶ�7f�1�"o<�լ|�{g�������Uox9v�5�U�OԐ���a5�&f�	�XقZΊ���S�,�E:�k�`�}Q�_kH�YmJ:O�9�r��m�0�t���q�����)C��P�mp��4�D�/'Cx��1��i��CN6����x�/�+�����n�E��"ͮ..;=����=nr��i2[�/����!i`�-�y�����y9�5��y���"4���`ַnt�ʬ��g.5Po2��+{�[�uҥƉg<nF��XۿN�3����U�r��k�&�ݻwS��$0�l6a�Yس�(R��.��ѝ��z�D�����m�\��`�x�"5�y1�X{�B��'+��9~l���2�숗D��k��R�_�HH�>�pu}����C\�5�E��@k1W΃B*'�WO'YN<���rDQ�[R�,aڀ�J
Y��4�V�Z��/Ih��4n��$O���
�o,F��؀��.�$���Q_�d���ž�X�Y�V�������q�r�f�P'0�o�:�Ա��4��Kb�*�k����#v��J}iRН�\��n.rKRҸ�'�ě%�E�x��ͭN�=�tkg#
��|���Թc���"�ÞZ�P�4>�6`���n.���vX�Y����J;�dғ�-����Eeg{ø]�$�y}���k� *����@�tw�%L�c��
c0|�O$���)��aA��b�DqH���$���α�0;��|4�`�9WY�l/< ����%��;�>�{��'���sl�	��n5������22'�LsU����ë�7�^W�H_}��"��Qw������ƨ��0h���gg������x��(��ǆ`ҩ�d%�2&F"��d60Kv�W���d[A�@��F�5��_(�xvv�$G��l�4	��D�`���O:���j�����ٌ2�Vm*��r9�DMGv]���P��u�V�J�#ߩ7��f�)H-!�0��dW���J��H��B��Zl�&,Vz�l��~����_��V�"6���z�`}�Čh���Ϛ� 1L<,�a�B�p0�V5��H�Ŧ��w,F/G�̌�������ŭ��c�$�c=�𭜼�8bUl�~Ԫ����������U�����Ҟ�֪
���V��*�	#��g�m����6^aU�8&��[)GĘVGvt�gW�w1����PY��̂V��0P,\�4�2�{6�.ǮҨ����V�P�����|�#�T�u�����vZ"�1���{FCY�>a�qNd� }�D5�Q�<�n��*W+���Ks`~�E����[��R��PܧK�.Qy�N]��2%�q��ݻ��F�X�ͫ``Y�1�l�<4 	��ӧO�z��VÒ�F<U���ݶ�:��2d�i���&o��/�c�<!�����m��>��� =�/˪SE�&���r�^*��n��U<ѳgW���U����wa�*�Ȍ4(!�&���i��D��[y�S�����'2P�3L�+�	��Q��a�����e��Ƥ��O�bcmw������?��7f�[T\?-���,O����JA�G�+�"Y�ǃv��nu�dJb�K�OTI1��I�S��>x�������1�)�^T��?髸�߉�Z��
�;��(A	�����p4�
�Zk����
�e�.�P-�RTm4����F�8L����Q��oQ�B����H�fss����QHp<_@ݶ��l�i6��Lk��b`��x_�8��:4D�A�C��[��%K���&���O>��3�z�e��T��Ȭ`P4ԙ�S1�J���l���p8��fvd�e��5����v/��� ��y�/2#g�a{�F��#�h�7�g�sH�Oh8k����|���g԰��f���"0��d����%IL۝�o��������%��Ƅ/0a{׳mSx.�?ǢR�r�h50�̲���Y�]O,o�uC���j5DR]7�& �tC�EՕ�B"�K5S�$�X��Za� ����K(]�0�C'#�\1h�e�u���Т/�J���ϥ������d�4\��7.�.wa8���IH,��T:+`]��o�ղ�l�g���ʔ�-�#J�tO���>}ؘp4#���\p:*���ja��wVP:h����0�����"��V�/We�^�&��ޚN��-��|���xbQ;������Q���lc.�^�����;��.����~"{xޣɸ��J�<;p���<-�f��KLn��#i4k�[L�8�R�4����e7��Cڵ�;���U^+�=���_��N�S�R��_�*؆V�U[.���V�Z�ZՖ�r�Ɉ�fjh��;�
D��Y�Q��o�ـ%���P	�����Bؙ�֢���#��?��o0vo߹��C^����������7e=�E��j�իW{G,���E���Z��݈�qx��#_�|��:���:ûmZ�噒=���棏>����H���{�'��+;�����m�=�.v�N�II!#$�����e0����cv0� ������]Vz��9�sOVMc�`P�V1Q]��򽟹�k�=w���ӹ!�2kuF�Aڔ����T0F����H�TY��S)�������4�v���h����O��`T�웯��L�f���_�B���co��R�F�����'
vl���G�)/X�#kj<BZBg�D�7�!P����3m��4?S��c�0�wO]c���
}8'��://��n	����$�@�c�n7�d�z<Jok��-!x|������j�O`pj��k5b���XU���+sO����]�a�_Ď=�#�ٌH�u����� Y�5�CJ���;W:%>�;O�q5U�q�R��JX��0K���jP���&��v�2�e�������T> �°R5��$���,`"%ys�8�9�G�ҷƂ;��z�� ױ��̉�"���iZ��h5Nև���wo�f����Z�ᖒWj�&3�%�����㯴U`*gG������f4��t�c��X�����*�OG��o�B������o���K���F(���K���!��w���YYfc��	���I���%,-S�����\���8V�r���ͳT�ZYQ��,<F&���&��>��Y�^�T�����Ɣ�Lɉ�D;v�3��{���������=^�֨	��w�r���D�����իW�t�?�=?w(O��t4eʧD��4�G��x�2���<3X��/���[^���X,�Y�q�&fJ*v��o����F0U����������~��y�m�=�e��p
��uFӉ�_d�Ng�)�ŃA�Ofk;뷷����Nƃ$�!LY[mc��d��4k�v��6�<�}9�X�����~���׾��q2so*jS�1a8��6Bۯ����݇��O�d����oo���L��{��Q����=���
�ފ�qr�._u��MH��6��#
%�D�W�#��Eѫ���l�&�?*#+c�˽~�h|��P�?�a���w��
�5<ǵ��0�9�[���#˽�܉f���g�ʌU�_�����˯~���Mz/0�P��L�k���w[�M��Ʊ1q��o5��q�U��9��3xV���ٳ��Uz�g���}f��$���Bdc�ʻ?��ϣi��t�`�GÚ9��a��R<������w�����	6���V�z��@j*_���O��ķ�g, �f��ADc9+q5b S�b�Q'�}2�I����(d޵`�b�I�(]��Ҫ2�\�Z�U"���4�'���D�:�p����ړS�z� �_*��h2����ٕ�x>��-ܺ
��5�i��h֨�{qѱ�����G�u�ƒ�\�N�{~z&�#c'm�DL<�ȅ������`l������;0ڞ�n�GL�(A�'�"�T��t��5l�p���ܨ
�7au�Ka��v��)bU���E�۱�����I��ч[�œ~�������plL�S%Ēa�'S�ʓcQ�V��Kk��K+���5E���b�����Y�@���
58�9���uYW������Rmoo��ͬ�a2î������ݽ�榔��y</��eѷ�)�0�3��|��7G�}�{�f���/a��1]���=��	R��)��d8�o�%ڈ��C�Xl?xpDf��*��۲�t;ľ_�ܖ��>���,�F��+h������3�ٜxo{qF����/½�x��?�g��P��\�锝e�B"���S�8]�i�O$��[�*�߲����d�2Ww�ɘ�>l���&�v#h��PM�ѫ��B�~��a�>��gx@|���K<5V)���tyy��/�PZ������:���T�a�������;�����^��pQ�*���c�.�����1� �@�y�H%;��)������?��S
F�0:�֫V�7�|�[=3��*��"xi�KLޱ��P��=`4}GG�ͮ/�ԇ���}ofϞ=���T��R��8e�t�� �C�j%>�к����emgƅqr���_��ޮS�r����Ef#�\��eј�Y�r0O��gՍQ0n4=��� u8�0zqB����2��w\�s.peB�w!F�l��S{�ЎC�Q�qttT��U�$�Y2��=f�x�����-���B'����aS�Lm�B����]ZZa���}Z�KS?,�o���5`���pr���;�U�R��k����W����s	��Pf������,�8K��6����؄�|�7�;���������(��trq��4m�P�^vo^�[��/_��������٤��V�uzY�������FAd�Bݣ�#L��U��z'd������}���U�opvL��:�8�3�ky���-�V��ţaV*����bg�N���8;��7��WW������U���$��OO��0�^��7O��E�Qd��f��΅�}V�ڡ��I�^j�a� ��9��:�����7���n���ٰI�����&`�Y~WlK͉�l�����܆�5q�1�ml����a����'�YU�+Uj�?��믞��'�J�sqP�e��?����o�\}���K�l&��o���@��j��7�J
W��/�=ǟ���\|���%e%��ѽ\����J�;w�XՎd��G'����׵f�h���OΛ�F�J����g�nS�gx�|jm*CZ�kۏ����D,�d��]�O��"�x$�C��Ʉ��f�/������=��O�R�/��/`��ſ�[;0Jۭ֒
ݓ�hhj��ckd���"����%�����T�;x:q��蛟�~)'���ӧ����������KD�IJ nQal�ja�%?�MȯD|��fo��s�8����x��qk1lzT6�U<���m�@N�`��T�CD��#fH<CḕJ-��i4�gF��_�c*'&b��H�9�^d�2s�y1_VXs��F0S�{�ǰy|xT��<x��̆���ȯ�La
)��#�1�Tq���y6���i���lW�W>��XQ��E)>w��
�kqhQ^��GXKK�pG�m0nu��d�nd���a�vw�0�&Z�4�Rp��C�Ǹ�A�Q���"��aR��L/--'s2�sNݢ!�t�(�����A��PF�6E&�֖��У��]�1�FY������d iN��%��)a��pL���ypx��;f&۹���hδ-a�a��o����hv���\db��"qB�� �1��i�����C�N����E��=�`no��'���Q"�{� ���{8z����JE�vUbo޼���D{Xj�~�Z�o����O�#�!-Bq%I��+�"�f�U��j1�����x∃�D�$�jt�ݙ>.�$�<�2I^&g�ŷO����J�t6no�����#@�7�ş���U\J=�<�a(��e$�}��Xw��ŁڴT�G����Mn��rfq�^^��B�3����D��z�)\v�=�������a�E�#>�����f���__��ፇ����m�6��2�f���:��"S��q<����Y,Z��.�0!�uo��կ�
h��L���U��j�H�檗�lz��BgY�L���4��f� <7!&���˭�X�5��B7��8a�z4��,��/jf����D���X��UY_]�:=;�q��L�5�=�BI5֧|فR=;��[K�}���~�bv�#r.D�\������X���R��a!av0��0��m.��F	&�h��[d���0�0p����b|�Q,�#4���E����g1��l�9ծ��U���E��7�W�dqW+�s�%g)||���ӽ#�|�ki������{�����&E�%������^n5W��i<�]�XN�.�Y�b�/�{#,�sgFWQ6Y0��Dd5Bv\n#�X{np�������R���(�-���5,�N�����(����ٽu�{�e<̓fF����<©��Q�{'�R�f|��ɫ�;6S�#IgX�AV+U�:Jۍ�R�NS�ќ�Ǿ�޹s�d$���p`[4m7�Ͽ8[][)WJ��f���,�؎��{�l!�.�ƭR� ����L� �ǧTU�����Z&��\�ͣI�c�ÐS?��3����L���$�7­�7�3#����
+�J��:�`<�Hk���`�<$&[fEN�AL�L	<��;Ȅ��|��p ������iN�B1,l�<V�s+÷���c|�<E�έ�2�{����S��9��{8������3nn�W�E�~sqҐ�6���?��={
����u�Z+I<{��țl&j2���VK���/��ᬵ*��pb}XMܧ���z�S����\*����F"`3N�����B��pm������:�g�
�0&"�ñ<K�ps��覹J�

U7"˽���hb%�f��Ǹ>9+]
�ÎY�A�<���?�{~nlD�ʓr��tBOx2^)s����2�.[Wqb�&z�=~�g ����������I�JJM86���O�m4����g��'y!F�,��f�^++o��뛀�d��&_H�Ó��%��*�ai(-��C�$~c��X5��_^ŊŮw�Ffo�c�
�|NJ��Re#���?�
��%������Q�N^�&�~L~<�nm�6�d��w{���ؔ"�xjj�.�jB8>�FV	��E����Y����&�$��q�{|���K���� �p1̉�G�?��?Y�s�$��L ���ef3��O�-;^�!-���?:9Àb�(B�GF _�.�죲7�PF:'&D�����x�88d�H��*P>ay�R-��p��b>2����0�jx!��w�{H����X�#�V���!6�����?����c9���dZ�g8��hG����^��`�^����2A���X�a��׫�H�bx5�v����X�G��#<��<ţ���60zl;Jb�q��0ҨW��?F8�7�$N�4�ș������@�������VJ �Y����]A}02�QķZM��U�t�G#�qJ��Z�.��|m~��J��3|�|�w�O�<M%�ZO8����
�kq,�SaFDm\	y�ڝ8�k(�0\���]������!��4���H��EA�c���ձsgS.�k��aKBv1]f�R
�GT�]H�����c���oO�[�VI�z��c�-�[R�C�w�Аk2��,����g�L��j��Un֓9�1��_��p�23�r{I�!s��e��xgѪMu#�Q�O���F��~2����P/�����|�'�y"��/5���.���%��טjvlGK���W_}�w~�;�q<�B��̧��hP+%OY�q�q�;��&i4�����]X�ɼ{~*�h2�|K�}��	��韖
!ƽ�^P5໅,���x6�N��
��;���&8�T�����=̽\�fZ��=�5�ax7j\��(���\�y�fL�Wq8�kk+����_�ݿuk�S���U��d�kRhacoX��Wl�*�=L�,E�>���&y7�v;q�p/�X�LVth��m��~{L��=#�W(���x:�?�g�4�V����w?������Z������a����/a:�����e�$���	@S-�I��S���U2����e�MB�*Ċ#�C�Vj�;�礣�0��I��ly#�����5��y���g=�_��[[�����s�������̙̦2F:n��SL�!l/���Z��糋�BX:<:��c�G���aմ�tgp9k����6n�p/��aI�WJ�(iޒ�s��h��</H"��5��0�t���iL}�����N37�)�/�*L}/�Q���2��*6шU��E�ٿ$9n�t>��=�������,�^�a���T�0BLKD�KaI�cB��F�XK����y�.�J7Nit}�C�e���md��I��[�@g��ka���u��f���t���2#�C�A>�l���~c;:(������p4*E>�1����Q��q��I�%�����ș�g������d:�\t>|�� _�����C�+�0�>��� �����K�v��^����rc;&�LD���l�c����ti��3��\�K��a�}��:��PT\��7i��O�Rj���\;9!-S��	�z8o��C�l�(��N-`���R�� �N�A䱛//_��/�F \���8�`��I4$/��r���z�Xq�"#)��j&��\XV�E9�8�KX���3�z߳$���o�_��d�Ag$疙���-<_`�n;'jUz��&�N*�*���+�|-�����+3��q"%�(���//{����u��ɓ'�|��T#
z�M\��軭�m�O�<I�mH�Hm�S�xrr���ܠ����0��������B�15�˵g����1��z��GÒ�C���c����w�����ILB�T��Q�ѷ��t���ck�]G�U����u�q#,�|3��e��t��KEQ��Vܪ(l���0��\��3!����2Ӧ��6�b���Mܞ����@^��:�����+�M�����~�ɧj`zw����:�_�5�v�Ν�)L��p)��m���`8����g#���ٗ_���Z$Ϗ�OMHcw˹*i���?�1�O�J�a��\��:�f�}�<�P��y�t#��7M� �xT��lb�����Z�\Rx'l��yG>�V5�P[�}�P���.N��ʳ�`@�<�Y'�i�A�;BŪܐ�a�������y�_K�[,�Z���P�J����\I󰘫��mmy���r6�8��h)�'��{��$7,A����V+����5#��։F@��3���~���q��0��h��F��M7k�D�hѡR�*�j����C�T���z�����7ߔMm�10^��T���կ~�w>x� ��ŋBXĚlLwgց�kX�֒���%ַ딭s0t�r��n5ooo}��c
���S����ec�7�}�n�����fMs��?}�t��NX��7~1�i�tW�ۍ��J����P$��$3���P� )�n,�+�M��qؙ�...Y#b"�h鰵�I�7�yA�L8�d<Hx��wqTʕ�w�5�\8 ö�I���w��7�ĕ���Y�.�����i�X��+-ز^w��L�m�Rt#�Ȋ�!��]�wom��g㉛�q4?;9���O>�r���_|�C�W�&�D9܂��JDp8<��Y���M��M©����pG7	B/�R�w� ��4���x5y�� 5Ϥ	�/����(�����K��܅־��p:ֱ-iq�}��7,�`�Էh���x�'C1��p�����"�(���'�B�^�����6��&+��޼$�B�Ƒi���ǘ��1*�zo8�Q!�à�n�F�q�z15�Af�=7XZgn�q�i�g�{|�N�8�VG)�G�2�QN���0-�"�IT�D�%�t�{ç�<Ǎ� C�o���
��£���������Jӊ�E�=�;/4!�<�!��v���8��
3�@�z��-��N�O����t�RÜg��:Ob'�tc���?�ى+xƊ���h2.�̼՟�}?�Y-�J�8Wݵ��%>���}�^`6��8�.I�g1>2FK, ��^�)U؜h���Yպ�й��B���?c<_�~������6���9���jCf�&k���҆GƖ?9c2��ݢ�G�v4��f��1Đ6�����<}���,-���,�B�{�U	a`���sK��,�:lT)�W��c�\��s(�Z�Vm�f!-�,�qQ�%��:�H1�dF�E��Ɍ�p`������S2Kon�(��K��=���;8���pK�	O�����Ya/�ILw�%T)B�u��-����G+����>L|;��֧�t�3�Ε� �Zt�4��2����d:v_jB��i�h��X}�x.��z�;�q㝤����h�����ʧ��_�K�?\W�G���Յ�{wp��R*��:b��EZʿg�HwkI-Zy�r�q���]��$0Ps�Z!2d4��\Ql�|��.f�9��
\�gϞ��� h��q�D1�_����,f��AHM�p>��� A�p���Ŕ���P��Z!����������co0�f�ʹ)Bް;��ԛ$o�by��W@���N�tR1�7�|<����2���h*MM����s������%��,���%�,��z��1/0UU���J,lb�GU] ��l`�CU�&�ެ�ly�٘�8ͤ����h./..���w��YTZ)���7h�k��E:�Dm���]�/��
]�Q'�x���N�$]�)
�P�Cz��������Tx��>�����������m�D8��+�T�3Y��X
�P�>�R+ۡb���"C�_G�l�y�7Fe���w��](�e���Lܻw��Çx|����[�~�j�?�\���A�V	l00�=��jf��=�S�?�y�r u�*�6瞙� ��w�ПM����ݽ������ѨZ+F�Z��.!k�;�Za���׸��۷�?>I�����x9��NPj.3W����;;[��Bk�:=r���H�����?�����D���,5{}��gF�"VdP݉S��"l�(�c"|��IPzae�r�t��b�]'���_���.L��������7�{B�����͢V6���Aϟ�%Vk{�!s	����/�k��`4��4�ե�Ę�G�~�RYl�G��I륰����ɴ�9mժ|�^4en'K�d<���r�{~�V-s��T��H����&)#������36�y���$p�)N?�K�xڷVy�$1�Q(O'c�i�v�tnm�*;� 8������,�D�?�w:�����.��d*�K�e���{�ч��Vgq��j3͂���b�4l"�����u`��0���_�ӴT��Z.��$8�k~��Y؃�L��������յ�8I/.f�	c�R=v�<,f�Z��cP�v4�A�h`:��.��,
�v{B�$z�uLKM�;v�T��r̢Y�R�T�P1���Z�����q��`�������фu��8
��r�x��Y�0�_.G��M?~�H�?���R*��w��[p������sr��S?Ϧ�t�v�N��9�TKy),e,6�aa���4���C���R���x��Z]�-T'�0C�#��u ��>����1�<N07̹?������1�AV�K�?�S/�Fg^�I)ťFV��,���۶�r:�T��r2+���j�qӱё��ը#�S7��V��<<;�(��2B�j%�8�u/;�W��{���҇�dL��Z��V����[iԙ����bn�R�������e���x6�R4B�a1��F��c��s��K�&�9��׭A�Y�Z5Xm�n�B�EV���,�.�g�o��o6��(��ӷo^���ww����0`E�bD��������'�T�����?�P.��l���gGg���eL}6�RG�lf�b|�F����Ͽ���_��_�M��:�M^(#x��Z�.�*�����3��N�ѱ���<z�|���_am-S��.�R�G��a=�Q`�c��2��ͽ���`�R���_\��O~�9���!m�����Z�X�᫊�	�Z��7b6���к�89qe�d�K;�&VD%��Ҵ[�,��v��{�Z����d�BA�&���ڊ(��s:���+�!�~�Z����s�1[���vUh=Ҏlz�G�ǗWWq�	��X�d�5e�V�J�Jn1�.��5<����D��V�Q��w5�xa��n]�xe�M�Bᗱ��X����.���M'�|�j�b� .e�����PW#g��E��kuh����ծ��JK*��#��3�`���yl��|��ɓ��)lȃ l��>��"ӕ̃|p.ד���;ԜEo#�󊺰�0�B��N������V)V����3�-ߺ�I_�CW����٢dE��h�S<A$t�#Oc�Z�N���5�TU�-�t��	�;�?��׷V?����U��{��y��O?��uG�D�A�<�h�L6�R�D�'%C��p\�͔kB��ຑ�m�-J��ZWW�%1':&f�"m�ݛ�X"5�o83r6\� �����cM-5�����¦I�3�`��/0,�����q��'��痷n�Z]�����K�x!iI�s��i@0���_��+d��!RA����$�����U��0�9,J�"9��Jě��7o�^�|����q�����O?����8+�2����O�o��1�����ؙ�^�%�j[�����+�Fr�������(��^v�֥V���S�������
A���S�A߷�F$�$i�lܢ͍<��[��7�X���$A�qyq6������+��y�j{6�D�֝F�>���$7e�.l�����1�%�"�c�K��)��A�10aqc��0�c�����`<�k_mԫ��t���Ս52�NF!�K���s^C�Ҭ���b��m���Y�U's��~���K��r��魍���;?��O�pʚd�z��RTKE:��|f	�������ti��$��O_�=4���
�����'�����&1l�K� |�y_�X�_Zj��cT$	O����湸���ٸ8I����u2q`n����B6c��l�\�?��MX`���8	��K|�G?�3����78�4︓��x.1`x��D�9�ND	I��LHh4�[X��T-AL!�
Kb%k�j�Y?(x9�18x���[cmnnb��P̺7tOV��'��~�������G�as14�ʎ�T$A��ӑ���NS��I֖�ؚ��t�&Ҹsz, �c��ޠ��4���z�gǡ7��������ʗ_~�a��d[�t�t�Ύ���,�2���#��/N) Y�t�� �~ �a���z:�O���s}��z�P���Pr���+}�8�./{_~�%�ߏ�1�O�&nJ�G+�1O��!�N,Wx٬�E�l��r]��5���x��d��[��+&���e��`�wp��\]'OfJ���HlT��syD#CCж�g�Kl:Y�=���[YY׃��3e��ӾX荈�h䓹2T<6䃨�K�?������T��q�F��>�I�r_���1������.�-� ���RiT�:?�"�J�cC�X��8�Z�&���+t������Ƽ�$b��V��b�ܣ�P�%��S̴v�O��v�.�&8M�I�4�\S�`);w���3ʬ�f�)�;�3W	���N�<%��|��l�H��h�؂������޾}�?�~�e�p~� *hV�<��x�byu3���ih--�|#� U��>;�֔d�=��mz��S{�c����E噲��қ�Xއ#�H[�TW�'�4�<,eܤ��x.~*�������<H�8�_UE���Q���d�:����U�#��fK�g65�Դ��0�ճ��>�����cLS�H��P�f�"ؠ_��X��%)�D�T},�%s��Z��H��U�g���an\I�o��{�f�]Q*�A���4���s�`0;^qW��	<����B{�5�i�4w�UW�A��3O�P,>%����Y`mz�z;�6�����8$��C�́�z^��8�����l�֨�'�_Y_��b&q���t��1�����q���==e`�`F1�_�T�	@a��J#�R�m���ɑ�C$܁5�������grDX��Xw�F��g��Ćė6�Y��T&��;��[�����ՓƖ�#�;�Ԙ�7�fI;_YHf/����[��?x�s7g/"X�;U*��Ǘ��K�./�\Yn�Ʀ��ŵV�ZXT���߹s&�X,�#�@�P��"a�Ґ'��x�tV��(�|_���5����e�h�mYXYŘ�鐪��E��cϤɾ�<���a!��Jbib�/J�w<��U�������{�����M���x:��o�)�͍Ux�0=��NؤV�ԣ)w��{ws�^.Kl�JF�С3K��xnt@lV��3�n���q�^��8n��^�8KRx���3O�=yq���~@��KM���jg��抨�q1zJ3们����k#���k& l����������٠�Ѭ4�M<~��A�(J�i�OM
4f�.�gN�uz�v�z��Ӯk4JؖX9�a4�!$f����ɪH[�4m���JYتz�	���\���]��{���n�ZZ]Y�<�7����=�_�#��!"�G�~6]]&�+y< 6�M�>��x��'_}��_�rd���59��Y����K��k�+ֆF.r!��ꐵ�{�J
# m-/��E!}FK�����ƒ�,��-���y/Ę���&+��_�9�d6o����|���Z����e�x4���<���a0yGk���T͖�VyN4�{R�oi�>;`"�@2�Λ;�1�
U�{�3���șu�pZ/���*�^�_�&�$�b���m/�)DRa�R���i\.��$-��,���1F~F-�P|!XQ+�k���%9�\��[]]�]^L&#<�hؓ�"��o��.3����!��Ju>%�
���oV��	Ip�D�8�[�̔EߥHƥ�m�#kȜl�c���S�Y�x�qB�N,i����¿�YVV�FqTo�d�g���޽;�.�%?�b,V�@j��J�4M�oÞ��i�n�W�Խ�����_�!������?=�T�/~C$T���^����b0�_�o���XsfxW�x^	C"dyʢ�v�H�o��!����z�������P`�*{�FI���g$�[^���Y�n:�=tܶŠ)-�1fxl4Z��i>�k䵑�����I|��h��uuA�B�=�����KeV�xUči�9S�X�d^��Q3���Y���� +���\)�X�>i��$̾��c���� ���\~��߇+z+�X#u2/J#q\���X9�U�qȇ6jو=�ւspj�}��]����iM��O�<�/,e�~�ZH��NWJ�����^�S�w[�U-�`䇰��5�,� ����su�)eN.m���^�z�M�c�4~��J�Ǐc����Ip�����KIP�4,�*ކ�gV*)�W!qE����ؚ���4-Atz�ņ�N�B6; ѽ�+|��Tr"����l�x;�.	�&=ƪF��mb��S��b呁[�e�y'~v�τON�GjR� ��S��g}k�ȋ�@lСI��ո'p�Z�q�JFf��0�Z r�!�q�W�^g�:�UT-�Lo�¯�\�9LbjP$}�������)?OK1�Ԉ��p�x:,�+P���J�.�EC\�hXM{�}f��[5rR`k �jV��#�.UQ��s%a��'���R��\:�?�쳟_^vq뛻ph���#��qrzl��*%z��x�Ew|�л��@R�`I�����
9��|���
���h�.��F�[[�8a�75Q�$��Ir�ذ������<�$�a%�Y4�3��^��eJ~��������I�{�����'�1���7\>�^�9db?���/��}�Ե�s�,�B��I�"a�"� �:�u<�tҰ?PT>�L=�(}�8���,Tw�q�����d83�)o1�0�n4b?�J��F�j�$W4��f������tcf��d������M�ln�wΝ4��y�iS�v�}�A��%ܶ�>�B�+u�u����H�x,ާB������1�Bڴ�ژE�+��B����&���&l�˗Oq�j�rM��g�r�eY�-W�i!���-�Z>�.;�*O��A�����h��R�nڈFbQi`����1�}���1��Ms���q10�[;ۭ���9����159Xj�-|�=vM,�V�����J�v}ܪ�c�qW;T�0���������X��YX+yU7.���BךiظA=ƂQ��x�.�7�[F�'1�Ŏz��deFS#���9v���<��M�F������;g�����;�F�Χ0��1�,�'�&J�[\؈	����+l4���Ɔ���@	v��Z��H�Z� l��x΍�H���\
�^\v�H��-Q�G�|�0�b�����`��ƒT*��J��5�u�>+���Ʉ|q�
9G�g�s�q���Kj�;a��v���/&/֟�~X��A2��L|�C�����zkS�=�%~�ܽa�V,"�vFn�7{G�^gr}}��/&����+�D������nK���G�R���N���E,�=iIR$)}\.�b���eD�+ �c�v�{�Uq�af�.�>�ꠇ;��%����T��L[��!ШR��4��[�R8�{o�R�>��R8G�A���1��?����</5�X�ߚ����lz23t��m��c�%�ï�F�8](]�~(n	&�&$jX�r��ф*�X�^Gq����0�-'�:1��#2�T�W�1��8�9���
��".E���Il�%�bɩV�J	�	"��*��o�"�t��9Q���+�Ȣ�~����J5��0���\�+�6������@�7Xm|��K+�XV�����)&S�rk���̬"BުQ_n��p�f��ݻ�\ǼlT!�5+-IE����_]]�b���V��u�+b��MVdw����vrb?-�{Wl��������K��񠭔��:%[��;\ъX��zd��T�d
Ԃ����t�K	��ߎ9�	I-s_���s�	��x.\�>"01���:�tRc��
�=���5_����K�,Y)���{��^�����{Fqe�仵&��#;��j�*s��)%�.�]'�vSχ�gS�\޸����$yI���s�@6�P��l�,3J��i��ݿ��PD��Nf�9��H����'��D}��j�U���Ȭd�B!`�ˣ�Tq�*YSj�8�K�z����FwȰNXLM�`G�X��m)���Ͳr������\�ꗳ�>�n���Ik��b]���2�{�M�m��Y�c�7�[L�e�$�@��Nʁ�S�Kr*�g��E]GZ��7O+&w��J��p0��&����sp�0��f�x�޴Jk�g'�"����Q)�WM�+K�~S(�����.
�׻<{xg��w	݁3N�Qf��� ��n��X��q�76���e~� ʮ����`�J����0�%ɯ�`0�7&�W���%�ޒ����q@��kVJ�Gc2ݺ&ˣ|`�\�]�����&���-D�5���G�]+����8[b��U�.E`��&%��d�c�W��䰊p�WW��t�����;��0o5�C�~�m�������幥/�m���p�p`e�Խ��5eBp00�[�"��E�0��67����z�捥�����r�:�UKWPƗ��F��XF�ѭ#��q�����gɼQ��ʻ�q3R�#-�JaI���;/���{%�]��&��^k
����i�~O=�t�-SP,�#[X��r1����������8��FŊ���y؟��i��[�*J����Kl40��u����K�n�͍a���.>�駟�f����	�&�����s�Tj֊hIċX~����� 'R�� -�D#�9}�ҍ�����F�=8_s߿��~�JxQ3�?�\pn0,ޘ������jAyE�K��� ;�r�Ba�<I��J�$���ץY��S���(l��3�b���L�6>`X���<����=��^���u�����y���������Р�Rׁ-H76P�8t���,ܸކ��&�Ĝ����'��������l`�ֈV�CTl�̷^��y��~W�����r����]�wB&�N$�L��y4�Y&���~���h'ԢeͺSI�^�s���nnzw�:�,[W�xi#�4������t+\
�h@��;�G��ѓ~8#EC�s�.���͛�^l��([3�`�X��R+S56Bl��%�K��t~�T�
4C�X,,R�v.���x���+���e����[�Y �{�"PU�s=��)�='x�p4��>|�K���\FܙE�S��>��ANQ��JbQzS�[������������j�h�A;���6��V1C�N�q4�F��q~�~�&��|��㫵������ݻ��{�E/3�;�RPzw���MYW��v�4��AkC�ཻ�0�9�c�]$��zsCf�>�<z��9�~��R��f���83�����V����T�I�߳ɚ2_>b`�u�N`
�fWgS\'
,�R��{���u��#��V\0ǳ���ЃW
���x��&^2�"�ߨ�i�AȌ�G�Իw��?����Zi�<{�,��&T���.�Ǔ�L����jsߏ���J����rM1(���F�n��).�t����:�SƏ�Bh9�O�O�6#e�I�+N����޺��j�|�j6��K���^���D��>�E����t��<�����K�zz�{�(�s��Ew:��޽[.�*�rgz٪S݈l�u�v��8������?�����G��W_}E�k���N�ц� ��Rx�������������m��o4�M���A��1̸�ɨ�6y�|���.�.�F�,��SC�2{]ǆ��w���GD�Dc�8U����;�/�C�w|�Y���c�qS�:�e�]��'��qF���hT��-q4��m�����ک�[W�ת��d$fL\m2��ky�I�y�B���Ĥ�
��J���on�[8�������8��.*�i�;�V댒'#7���a�e��^�T�������F�����J�t:]L��!�1x��	B��R��s����N��8�r#5�9[����X����:�Yf"Ig ����Q��;p�NeX��ph�ޥ�s��q�5�~a����c��ZH�&������	I���ꊕ���X�[M�V��$y�"���!Y9E#��\��:Q|{WH~�}�R��d�r^,]�%�q��Sl�*s����l�՗O=z��
�_[YET�9;�X]����ӧ⟏���vU�K�t/��%V��<���SBl���g0��;��HH��vA_���X��{Ὲ_1��B�'ccc�Ϛq�ϒ�DR9�q�#����T�Ͳ���N<#�|�I2�+�h4��	+o= >A��g}�2��Abe�tu����>�I�W���)��0[N��<;������^RBe�X�\�V���7�U{)����Oi��R.þ��C/W\)���頤V&9�&Jlz��|���������|���_���v_(#ސ�)4F��P�q�2�[́Y�x�'EЇ�������<�� sOU��GCeN12�i` ��%6I<�ʁ�w�A\���?hI�����&G�R����d��.���{�����~�)�k��d4��"D���Q*ލ��klY��∾
&�w~^����9��Y��;�~Q�c6��J���W�@�|Ye^���%8bp�g����m�Fmߊ]Q?�c�����ag��9�g�����R��ًaA���B�|]+�G(A|G��i�6�-6s��)=�M1�pr���C_e!�HU;��ՕT����%�F�!y�pV�[�t��a�����v/�w^�g0�(�W1C�l�U���2{���5��������d�9�w��w{�d�s������o��i��Ɨ����<C�d�3��k������G���K-�R��5��쑵3���T;����Jq��=�ݮ��q��-xUm��҆�	���hQ'�;ՐKu����,��f����P����H�B�;N��^���\D���NNZ��[�L~:"A�����SQt}�Rc���?����	�ь���o�qsOg��xR-q2�4�VO�,�MwT��z�ɆŒ��q��A,�ݤlI��6c����j��_!��⸟ǌ.�S�����^�~�\D7[��t�����(]�e����9US&�R����T�WF��hܛ�a��6#1�,��(�ո$�g2�*���E�Yk-/��N*O�~�8%4���B���յ���ƣNh0�3�����߭l�������V@�[S��+�y�n�	J���>H���W�;�B��dms��h���9��W��{�í�"��_{�o�1�@��!s��w��j:ލ?~�ț,��y泙������<�\���8,��[������R� �Nhl&��C���+� kwI�VWaJΎYF@E1vH�\+��$NY�gpR�TjC���f�ˊ��"�0|3��+��bi4���Қ��G�y�:�h�;	
�`4���1��t:�^�����G��Hl��4��ߺ����ի�o�n[R�xO�\)W뗽.��K+\l�3�R7vp��Z�6�J�%�DKxrг\]_��'� ����������by�Lc���<BE.�Fs:Oj����Yw2�U��].�_s~�G��܈<�v-�����sB4��e�嫷�ؽ}�Qke��O?����:]��[���ك��V7�aΪ��<M��9읉��՚�Q�W��R�=��oZjq�QW���h���;�P��9�SX$�L�-��}��y��M��Vd�1�D4t����=o֝e�8%�0m�KQK���\��\���L�Ot�����"1
|����D��&E|ٳR���)''H��������ݻ�1��EͲoI��٩܇��U����~�����-8y��_�x�(��8�C���b�[Z�R�`��������=y�0�?��O��6���U�Y(oX�O/nN%� RX�_�o��� T/�BT����ӱ�>��g�v��w�����8ݮQ���^�'T�����_�����w��?�g�}���v[q�ڗ�L3P"�������O��?�o������Y$�����Զ����^��?������������7�w'KB��$D��빵}��BƲ�G�O][�PhŊQ�4T�^י�.�)�.��	���u�b3�S�kR���`n�Z�"�z�Z^�=Bkn������zD���ҚܬJ#�'f��h��<�z`�aq�>��������ѡ�[�������y+�c�����6��Im}�R��۷ՉB�m:Q]߈3�Z�j�s��q��͊�4�EV:6H�5|�d�>�Pv�y�^X�K�ҵn!z���-���dr]l�8ǹB�;�����o�������zq�EB��Mh�I1U`a��3'+�H��*�m��V�~��� bșm��fC���WҌ�Xۊ� ��S�.v��Ǔ�Phu�au��e����W�mL��޾:�(�lDJV3�w�5W̓�~۱�4fjPo8��������cl��^�����0۳�S�x:�A�{�)�<5I��8�����4%@ɣ��0��*&�۩��W�E����pl���s��4#x|}�mJѸ'^��a)�l;,�~�x�Vu������S�J��2���p۹i ��R���P�"�UM0'�56c?඙�p<AW��`s�K�a�3S���˽����Q����8$������%-���	���!�@���� E�M[Y(�]v?��gGg�����?�%�������W����X�6���g�GǓ�R�;ud\ǽ.��.u�x�ٻ��������,ѵ �D�p�99�|����;�����ɝ�tw޴Tk	�Q6���=m���@� ACg5��]���p���Xr�,�˽����c7j����R���|Ĉ��,�ő��bPT�^᫟u�dՍ�����͍z��*EϷo���y��������B�ф�BH��x�40��eə�*Z2A���5������Ƙ�k�E�D��.KV���ќ�� ��ܜ��2)�3�1j�ل�K�%�<)�W��r+UHXb�?;�B��H�~��O���m�/�s�hX �j��K���kw2U����w�g�o�E-���a��>�~��㓋����å�������_nmlb+ON�OO�=��=��g���w��i�x�g������fh~v�!�s`��9��,F>τ��'�ϴ��D2�W�׷p�^$t�Nz�b�X[S��7�M�h� F���)�K+�[��=
���J���v��^��`�ГrU�r��ѧl�.��+mת���3?pa�a��Z�{���D@Gg��e�Xdw��R!��4�LN%	WẔvc�բ��FQI�3��
�1Ħ�����)��aR�2Ｚ�����rc�Y�3����4Y�J����l��DP������OU����ܙ����a��3�����%?��67x=������r�Pg2ރ�T{<��`!�{�w���]���Ց�qnAǏ�����=扔�W�-%��f:��k�Q\s�b�7K��|P��qc��!�:���)b��?�����}Y���-�2�	���N��[e-��q�������7�|#�+ixV�i�g�8��~�ج4#�0�j��hǟ6��,-taoh�߾���vU���Ԡ �#l��%�$���n���T�)¤c<�ݾ����=�o�|OVJ���C�IZi/t�%�ȼ����M���>ml��DATA�Z%N j��j;-P˃�56_��Z-C{)���Աn^�l�6�S-Tޞ�W$�0�ɓ/_������������b��6���머�6��X�F�|NN�'�Ȝ��g�X��n" �.�
�D.��=��E�כ��������2ưѬ��@���`��ń��^��+%�W���4ND��C�\��u//؃bkR�.j|aB�:�a���t�Ό�K&��.�6H�/�� \��K��迪��Ĝw��v2#V�<SH�hτӄ��l(5����a�z�VD��X7X��\g������	����^�G��P�vj�J����X�p���zE)/�eέ���Px��%� �b�3ڹs��G�;������m��`v]�ʳ�~�?�fq)�͐�Ǉg�*�����p TKtloPP&s��L�����)�������;�[��h��������j����ⱑ, >�wp��ŝ�-v�-c����O?��z����2�&���� ��f{s�7�7���h�焥2��,IO϶�R���h�8�~��ܾ}+K1�'[���?�\~��,�w���w>x�Dn�k���Z�-*0�I�"����~U��XF9�9��� ��b�{~�z�%��G4vx|:E�f)(�.NN
3v��χS7{��Q��|{�_���1o����G�ɄFmg�X�ȅ���4j6ƫ���I�yk�=3�<�#S������4�$K�y���^Y��b��f���K���΍���"��(ꎢ���q����3�a���E�#�Qߋ笇�s�?R=Y0c��i����;�U�be��,\̓Rq�Fs�N�lc7,�h:J���dzH�V�T�-�E�7�ن�0�[-yWPf`���D�ڏGl��<���V���d1&hh2J۷oaX��ݿ�fb9�>;�u�``����u]�p���{�gG����n.e����{Ζ����ޣ��+�����	���F��[w@�ē9B�2"������ϪU ��۸�۷o�rk���!���$�t/�C�LO�0�be%�Z�m���z�K<p��pП�i�,�#�p���^�9���	[�5���h�y,�/��?�fԌ) �5����uu�{��RȪ�S*�7֛[����,M��!��S6�{��S����,��RP\��t^**��m4����!�,"L����,�vg��d-�p��j��.�,�v;'G�|6�K���m�4Y��Op�p�*/��I �p4U3!~��|l�!L�}����ӧ�j	�$�>�\RY:eCS`i֝�[�T�|��������A�h�b�r�(9%v4F���N�j>af�1�2����ݏ:`��0���w,�ap ��r��qyb��5N�k�b�����{�O�#\����qm�I�i=}px�ՅP���삜�p�I>��J1T�]T,�P�ۥM���w��"/l�_�U�峯���͢q$��l>�
�	�Y^W��cK|!����~v���������x��!����鸋U�.<u��S
�*��Į�Fu%�^h��!���P`{#�'O�0���ր�N0.��O�P�X���G�A�#�[���B�����M��j�C tvr*݉bbܹ[�	�R�5�rk)����)p0IR_Y�G޾}���SA���nO�U�l2'yrrF�-�X��;	�������B)�����A��q>3���!����4�'pE�DCo5<G9�+~��_�[�A��'VG�����*�Ӊ)F�-�y��Z&<*©77}Ӈ'���@��V�O��.�
suuM�#u��m����x��RL�ɍ�u�*6ݽ{��x*�|di�r⑥�8pd8o�L����@Q�.ܨ�H�BG���%B��Rc&J�Y��X·��X��T"�*("x������L���� �5*�r���j0_%�1�4`���Ւ1Ӧ�U�_
?�f�6(W�/��������V��#k���������ZY�L$�I���}�������<g������5v��X�
�b�:�MX�X@,u��f�0�Ͷ�yq}#6��~����s���ڒ*��1u�QE�J���e�a�������ё��,���lc��4��*���x�7:,ʾV�l��"ubr�V����~S-��y:H����{�Lag�kl��{{�7������\�� �}Ùq�0�K��a��������o�>˘5�;�y�R_�}���>BDӍ���O���W�W6�VsK^�I�ڨƣ���VD�E�e��������k��Cͅ���L1�/^>�[��������}�6���[��U��f�����۷w��&u���f���g�/�=.��xO%���a�Ѩ�­�~0���bks��N1PiZj]d�ĝ�[�ĵF�5ۊI����d�Jٙ���~L9Il;���0t�rJv�Y4K㲂Y��5lQX=�
��T���[�"�6F���w\�K�E��g����Y��\[nblc
�U[+��;���[o��;oٷk&d��C�+���oSd��_}}r~����ZZ�O��L�&�"�A�o���l���H
�Dk��|&O*Œg�[���66�,J������0�S�p����="�r����Cr
�Y���] ��'��5�Y�W��R�$Rj���[�Dao��5$b�HYPL����2��2J�FS��#;��8�0#i��v��-���'�ʥ�����e��l�D��`��h���j��+�U�YU�L���p,�}�իW*__��^�I�{]��q��^�]��Y��� g�O~��Ȋ\��J���7R2Z��ׯ_w��NF3.�b� oH�M�i^��7����K��Z�����ݍ���4X���Ag��C�l)�G��D��`�~�g�I��?��S�'�i6��䇊U����18�E2'W�'X*���O2��� ���Q��N���Ǐ��������'���'��tV,���L/�J�{G��o��c0PL4�}t	IB3�)�Rnf]�^�	kO`�x��)$K"��XTx�*؋n�JU)~C.��B�
��[b�B�un��_�0�cq+Vc�\�(���p ��m�q��$I�^�{xh��*KW����Z�%�@����=�߶w�xX�bĐc FtwuWui�U�Be�����"m�f$3f�,;3���'��'��޹!�x���;]�� *�u��$�]�	�!.�S{��V���Ǐɹk� ��5�9�ŰX���&)�%��J�V��.��
z$-�e��RU\r�|:r�.��f�D
B��ÇXiwo]��ݩ7��6b�:��q��Z'�\6�d?�ݻ��~��_~���,T<��GO��<�t:JĉkK%OE�&��X�A鯊�0����eqh�U����a�Q��<][��=v]i��'l$�QDL]
�&��8�ydS�{\Ĕ:���_�?�Y�Q�A�'�sMA๬�+�^R`FL9rVt
b �Ҵ���sf�#����(HP�ME5{#O_�.����R��`���[hZ�����,W�?��O��aL����0Z5[���؏�ƱN)�e��~��tr��LF�����f�B9�+�Da�ʒ�U&�\#l�,Kŝ���.��/�F�������S��o6ۛ�sf�N�Y�t
����vz�^'�I%���H �����0s{ۛm��y!8��McL�Ӊ������% .���9v�T��Ƣm��jn�]�5��|	?��׿�/�_���oa�c�?D%ǽ�׿�L�ا?��9%t�`�c���������A��lo�L��K������Y"��'�х�%i&U��!,���/?�;��\�V�.wN}b�ٞ��Q*ى�.!��alb�K���� X����&c��ŗ�R�Z.�^��ݶ����שi}�Lu�0Z�S"If'��ū�l4���/>���0��ޱ~�������q�/^���p���B�8���&X$�rѲs%^�I�(���/̟��ʋŬ���L�F�瑏IQ�F{�\�����Qo,���8Z.K>��r�SĘ�a��T|馫W/�}�����gn��"�L0�O����\��7ΙЬ������'���������t�X}���{��ϟ?�v	vb�%NWJ��Y�MF��8���dʵo�)Q79a�i(�W۳��Ǵ��ȄI@�rZ-|k죏>R�L�^�(^98>=m֫�3Le��Ƕ�����!��պǣ�X�Af0���ظDI]���C{�(\��I�+��s�7^�¦�;+��(z����-�5©V���g]r�U�B�tx�cC�ˈd��B>u�:���~~gk{��e�Us#�����5�$VMޮ:	�ȇ��*!����b;�qM䣄.X��P���G��������e���S8%�2t��^u���@�\�Wb���������^��Ta2�YP�͍��-�92��������{���Y�|*�������Y�\�e+נ����hq,R18$K(U}�_�cMy��=�ץ�|G�������=������%�mNЃ�#�z���,���WE\2b���Gl{�V��'�.
),��Mf�m�ó`��P�9۱��0��~�m�^�/�DTQ����E2!H%&M��L��d��Z�y��U��šީ4�%��ɚ3Φ W�JL����"����?�S�W;������ 3�9
��N�lǢF�ݮ�P��Y�޽���ʿ��Pd�괧�Z�Զ"��L�B�&�-|�uv�Tƞ��]{���)�;���/��/����?��d�9��{5�s_�o���VΫׇ���w����+0D�9WE�B���ѧQ�45u��۱J)�ڟ~�)l�tBqfa1����*��l���06j%�<x0����b��]�t�(Chi�Ƃ����!�+��Tg<��2�+yij��,�'F)��C���b��_K�����SN^b4')��۷�H��J,��R:7����ٌ�ɝ2eF1�f��I�N�9���h�U~�<a!j�f.��a��5��Lѐp�
yxs�;[�G�s���G��B���M��H�2��r��Q-W��Y�B��`�4����0�!�KjX�req`\�!��s=�s����K�R[�FmQJ#�|��M�������.ie���9�x1�:��t-B�m��|�=Ŷ�6�f�T>;>����ܾy_���=MV(N��C�V{[�tT�A(��a0_�0}7o]ñ�D+��s�;{��!1$��/��?M�����O�
BxB��A������F��I�'4w��h���O�>mԷj�B��߾���&^�����v�6���!�r�F�X�36aN�XB��t5_��mBY���~1��9,BDf�\�)uC��b��
��Z%h����>N �g䁥������Tc�U����K�H�J�È���o,�$����}Q�7��g{��Q��U�U��"^�g7۝���.��nR57ڭ�mP��/�o4���)4��?99��*9�έ�5�f���x���o����B��&��������:{_�U��*����F���g��r�z9}?�����9"���m#�r,DY�a��XC���G����D��?����կVq�駝��7�\��<ɲl���6W��8�J>⸣���b;�[}�l�b8�c��3������LvaQ(�s�Xͦt��4~w��_
�,! ���՛�[[$���(
��
e3$�wg��]��{��Y�Pfl�jPU��
i��<.��х��7��&�4V˅����~�wV�WR'U(�����+z�����CUOa7�-l.֛�q�T!������g&n~{��|Dι��Z�!:���~K��j�����r����ڨdg���1�Ҝ��␊Z�_�����>|�HIK\����.¹�$%��R�_��v!�{U'���p袛��Z#Aap`J`��G�F�<� `}[��l�Ns^�<��"����e]'
oܸ�hup��/_`X>��3,��O�	�/.\�Ǿ���Wzrv�6��7U��{��-՟p�8?:-�o�3�>��Y=�ḆO������l�7�������Y(VU��e�����Fx�$��7��W��m�Z��PN\<c�"ED�!�?�����pV����=7oޔ�6U1v�X��J� ��e)�`��f��*�]�ԩ�"R�!�������	o� ��gz�М
C�X�/*$��:wr�e������QMB�[bSv�9k���0�R����JD9"��LD����]k\on�$B��(X������V���2���W_����g������I���M�Yt8<��9⌇�=6�?��8���pr�(W#
�AX8f��w�1,QKK(�IO���KX�O>�!\���_�����m�	c���B���-�����YI�$K��xN(-\��pM|�e�I�4e�0���˫�6.�OJ�`�XW��Xgb�Z.^6h�+{�����H{Z(05���ŀ'��$c,��±V_�h��ؔ@���5ǻ$��� ����%���1D�b���-͂�*��W!����,�c��_�>�4f�Ӑ/�X,��0~x��5RT8R��^�ayU�ea��t>���r���+1\P���Қ$x�� 	�Pr�J��}�QZV�8��\���ͼ�q�2�����^�YW�Z@d�[z
�Ju|s{۸�Y iWi��	*Mam�ڙ�c��`���;;f�|6;;=���۬է�jF�R�ur���o?��˟��_~Y�	��e�qO	e�c�BtUkw3�˓�3㢇?rҜ�=~������ԛ��O~��t{���<����a�5��sl�M2�8M�g���B���V�,�l�E���X'[.�(�)��s2�V;����FP��q�Y�TKJ�:fk��ha���N1h5���V��I�\�w�.�^�R*Gֱ�h�����"��<7=:>�G�0�
E7�?�:��&	
�8��+�jz�1���%,c��݇��������W�[�+S96æ1BLh�����b�=x��\n�Q�N������II�8�^���0��������z�,͊eޖl��jP$���CF�Fu�
g+W=y��?��_�������V��a@�ۜ���C�^�{�?�Z�߇q����}�ݻ���~�����޹��ss�=;Ô���Њ�8��Tx�t��o�������1��s���3,���SK4�ܽ
��h���P uNM_kp���޽�����8X,;��7d��<�J�����5��ݭML�p޸���y3^��5[f���b�1�h��iBZ�$r(�q{>���3���1���f(�k��$��� \N9��,�s��i��yf��Ul���b$.و}%UՁ,�a��1Ļ<B�&�%���>0~��G\k��_��ɓ'�����vM�c�������B�ː�]�-�w�.�����V+��$�6��r�Q�Ҙ�?1A����?��<��3!����������sDԕX]>|%)(#:J�0L���ݕY��\E'�L<����n�"�2a?��r�*-�x�9v�Ա��&�8z���{W�~�sD?�J9w1�q�\�� S�"�14e=�q����᫿}�_�+�`%(-�\w%��G�5��V�p ꈆ��#c�P����͛$���2z"a�ծ!�)B[�`Fu_p�x"��<2�@ڥp��K����9���TǼ�E�f��*1�A��Ҹ~���CL��޾�z ���67-�ΩxCV�jMۊI�
���B(���>G�Ll�j�\3�QE5}�Ҧ%�� ��Z�T�2ģFO�4�R?���9~�ZmӺ@܌�΀D§n�~���ݿ���΍�|.�h�8���>QD�N��x�����g�^�~CHho�����x�0 �C��]�u�0��ٟӁ�����1�8��Ӝ���G'��
"S��It5M�+U�
ͣb>��D��Xg�Rʼ��Jۙ@y#��,w6���j��@
�Q��E@"<��?W{f���u��G���&�Ӑu���a�ل3�	�<��&�h�\���G�I�|�Jήe`U���~1/'oP�n�����+��a��������M��t��S������t��E+�������6���>K�@�$��W�tA���j����������۷�~��/B«���.k��n��-��`���궧��`(gG\7V�,�0N���a<-�XU*��>�["�F�S���:b1� [��ͼ�zkg������l��т�b��GLg��"�1�$̑���XΎO��8�v}o<�z��bY�k�"�`7g�{��jn�d�s~���O������o��z���ݷ�>���.b�&R)�����*��C����{C{��
�����^Ζ��0^z�{p�:&& ���E��v:&ų��9�\�ڍ&{��vGGV*쎚c�������|3���=�#XR�x+V#�G�QB��1Y�|!L,޾uWԁ4�A����)�oZ_ ���l�;�y_�M����ۍv�ū�®+[�X.C#g�9���f�+`��r� ���ຫ�QT�>IbfY�V(V67Uy���$���QxrMVDF�M�c�$�/
���Uv�K��e��c�u!a��z�2Zla�Љ�"8�-�9�Z�%�JMm�F��@#�:''�p�{wn��G�&ٹ�5�e�4�G���`}0�-ɷ�z�O��7n8=9�{�ܹ�L �R�Z��0��7�ϋe����V��n \�^�R8�H�����'���7�29�2Ds5��`~o:?j��<�^ S�|�L��P,����7�����4b�Ar\��T�y���ᕬ� �W,
�nJK1#�@RW��)g�̲�oW�q=��w�lGI�Jm2�O�,�g�Z�p4NǄ##�G@W-�s��c�2�!�drA�0����"�D��IG�1���|[�m��l��<8�ts�=�0�X�~�[e`�0~8��rpdv1g�(��x�j����<P	�g{.��ѣ�>!G�Kr�+yin��rV/0�A��f&'�gǿ"�ML��W+KT�l�b��u=�+.��޽�  ���ӟ�O�ZR<э�r�z�Bf���p�g��d����rJ6雷��O,��j��b�8��^)Y��bΌy�Ȩ.pVƻEQ�6곧�S���@��(�p��	��g��b�3�U�2Y��]#�6�C4�׮�"����C�(��(s�i�XSK�N3�4.uY+ݏo�a�0��&��z8�������m���)X�yR���zR0h�5�8\�=�O�u܌��yShw)p(��D�ƿ�w��O���S�*W)"5�8���!��Ld��x�5��J�"�2��M�H�!��X�&�4���bŮQߢ�?���F�C�S@cB��"�k�0���S[b�e�\S���I�|�Ǩ�D'ȭA�j�P����%���3���6B�0�5%3�hI�4�zY�s��#|���3�۩Z%LN#Qyns6�X�aD2�?�+x:��eN.�&��
���p�2��2�h������e���~<�T+�M� ϻJG��,��Z�d��@�0w�`At<$2�ŧ�̓5��5y1%m1�Ha؊��S���b�7`*��W�?���JT�צ��	������V�OdMO����]4n�o���3?%����_~)~����/^��Ž{���~�+��i��$JbV+�|I�ʨ����h����#�	��RÊgW��5������	j�T�zٽ{�0�xpö.�E����(����7���+X�;{�L��8\P�Q٭7��	E],	3�L��(����?F���_��.>NpȘdy�v����c��~�����p{{�j�g�[[���?8]�N���_e�k������#������|>L�wG���*���r��E ���	i�)�Q���IҌV�,�{�!��4v���:�]�Þ�#��WKX�R�>]�frc�l�u=���j�/��W�+�P����O�#��,$�e�伋� �<)q`���?n�;GG��f���d2�U���Ƙ�;���1\l�]a�q4�y��m��pY5n	�r�7��=������8���0D���CSd�;Y1M������D70��xw���z�vxz��A�y%��.A�^ ��@]���D&��I�r�X��YZ�L���r8�b�Q��*�Ofx��z�8X%�fK�f		Ƈ��INc��p;hR�DǕtGp��w�`���gϞ�y��9�8�1��*�^,�&�Ǻ����.��f+�/0?Y��q/�X6�$�;;[0���	Yu8�l6�K�~�z�R݋�Dš�bMo��B�I_��`��y�`��N�j7��r�=G9(K��N*.j�Q� ��
1�bp�����&�|ǣ�J'DF	�a����d4�ҭ����F�T���dR+U�uK�:Y�Q�Ug]�V�s�q2_R��c�#Y��%���j��)EH~����"���W�>92ԗ��+��I@�F���YC�7�� 	�7o�tL�O�|L(5��t�k���T-���C��B�"�-�B^��/�,V�������A���LkL�-&~�7c�H���I�O�>E�����
'��]�9�u7o����:::�@)��Tm�z���Ҁ��Di1�D���%�D�����$�̪6#�w��ɽ�19��r�p����\�j�8�T�Qg����T���S6w(��F�>:e���lh:V~�i됇yŷ<���"�P�є�#�zܿ�{U������TP1�H�"2�W��i��WG��r�T&Im�U)�,N��2/>Q�5eZD+17�aa/���F�z��Ɂ�$ۘ���y7#-ջ�%6�Tr��؎��uIz��C��啾C�(ZV܉
��C��Ѱ�Io##��tR�E;[[��h����ؒ�5_,(�lu�Pk��߈G�I����0���*���܆-&��4�,�V-ϫvWm(��::a74e8~Y���z).���BF|���bNR��7wɂ.��I�b�<eu���dds������Q�c�O�1��dB�^�fw�����<Z�A���Pi�q|n���.x84�"W��z��+.d���Ʋ�N��ֽ=�d�Ϙ1��Z�c�X��f�^��@����g�E�;(��گ08<��)'!��?�K\���-��O���R�Oq���cV;�R>I#L����xj��f
��>��S�?�p|��NL���l���P0�W�آ���4�S����Bc�0&���"�A�Xu67�O��ew��T\� p��E�jU{�/>��$6<;�:ׯ޼�ǚ$�RIjR��Q����yy��wt.λ�<\�����M|�r�@D_�XL'�<,Z��+���������O-
�`�I >����r^�* >/[����]���2�:�����ҫt:������Jio{������gcUr^^��d:K�l��H�gb��Z�t�XL����a�Y[M��Br�q��gK.>Q�]'�P �Wy����8~t�RV�|ܨ�a��c悰VKł8�X1�<s~��Ŋ_��Y�K��h`}�1�_X�Z��:Y�T��#JM�2p7p��,�$NP�G�6�5����h�����uX�LR���O�F��r�.NB�%R����]�V�x�7i��q����?����p���&���y��l���0�拓�9�\��	'�js��B>g�山;�)F��b��ݻ�������w�����On��b���j�\9�Ej'��ey��"����sk�cfrc����C6����>qY��d6���Œϒ(Y��xX*ۛ[�.�KC[�W��[�n��y��Ġ�T�k�7M��Eo��*J�����X?�p3�[��\��;!�)��^�Y�\��N���w�9��׿�OI�v�6vv��(\��B�F�����$$����.e����
���F��z|����`�a��f/�n����"�P��@ސ���ů\T��cڨWcd�p���3�L�Z��Q'Le��%:�@_2�����⤲�ΰQ6�U���!���R!(��������4>-2+���B0R.�Ұ|���kI��pb��'?�����o���Ӎ��p�KIbf�����Z�����c����'aQ�o�o�4S�%3�P���=L����5S͈g#��ՍQU���	�ȟãd3��UH�ܠM��ciSΩ�	`�.��b�x��Y��'0�����Mg�Z�*3��xS�֔zof�֜w!�:�2fC��6�m�nT��{�c��޾<�
:*��Wʈ�!s�C��C�{��ivs��Sx�Z���?�
"����@ǔ����/e:o��9�lZ������,�35��2kx>�į��9�ˠ]f�q�ɛ֕%y����7�m�DX#����4I/t6�vR��f!�Xa�ehw�3��I��`
�hBȡ�$�s��������5{2��V"g���g�)�����𒀊G�c"N]���.��������([?03م���A���]p�p�;[�LxE����NY[��������u�+�(���R�+�%��~�3̔$i����$�E�_���*��H�����d�YL-�e %����/���o�~����6�rN"n�s+������s��O����ɖ�Z��h�On�x����{��&N�X�4��fL�&�v�s%Q����G�Ә�.U��n]�E;�lp����I�F��/k��33��[��=�ݯ�*�d9����\��|�ς��ɛ�O�����}�-��r��,u����YW��DH��?�qk{#���x���h�
�d�z��{�z&��չ`�IJ��� I�>c���{@�||����Ƈ��_~�%�3I�'O�ߺu3}��m��g��������p�r��N�0v��M��
?x��Q���
l�͗�(�ͨ�k�~���q���	��J�-8$���2���V��n^n��f�ZH�f�\���d^�r���yȄG�ݨ�ew�X�[�:�O޼}�DY�2r�-WA�QœnooȞ��Y�Xr<��rƧ��
�7Ϻ]�������|_�~A��{����ZRh����LӘ��4ZU����MC;�<������������G�޾o�2��Ra�Z���Rf5k�;$������tF��8�X�+���)��/ss��s_<z���j�0�R��ϼ�͝���e��|��8��l�lLNO��*u^���s��H�m�f.��gi$N� ��6����$Z���j���|,������ā���y���Py«�6D7�͒.bX7?M��K/pM޸y�����Z޼y�9����� s��%C�\��F�7ofE/>:|��w��'#�,a�O�]��V�������S%����M�s�B��'�.O�k��ު^�40�~�D�l�ו�K[+��:�R]�j��%�����4\��ѩ�[V¥`��&Y.s��'+U��5f������ٜ!u�/�?�N�BaY�Z�99�be�����:�r��<X���뻩5*�F�P�r�����ŶO]2�|�΃���W��&�����]��:���
����Iw1[޽{o�dM����Q<(T���h-������8�Q���Ƶ�,�Of�q/��1�%#n6�D�X>$�Y�6��(0$��m����]ڼ��9����~�im�������KV�II˱��EM��v�X~��	^����3Ub`y�WQ�׽R|4�,��Z�Ep�ժ�IE���pP��L-����C���������&o< y-���F����H�c��Àf�b�I޾�
����	�&l>�G�t�8[����܄W+�VvAȨ�'=As*�S4����x4�K�F���_jS��o��E���(�Ve�CI�h�-���rs��rJʼ��4�Yk��$�&D���#}�ht�F+���K��m5����>P�C�b�ZÛ�$c�ަ +6�+|���s���,<���֋��Z�����Z��XJ��@�0R����H0v��l�TtI��3H�T�Sj���?rرHm�8YST�ͪm���g�D?����Ϫ{�.�Ma���r�"�RT��Dʒi
���N����b@��+;oH��U|����y��k��F�RlKԱ��ڵ��u��������)�#e<{��4����i�-��s�j�W	�%6#|/i�rE,]��c`�$�ʐ$d�B>{>t��4h���L���Uyٔ� ��h�����a���q���ٓ��
l��q��E;�X��^ �4<��ƖՊV�}b¹� �S���]�D���_|1��u��r;\����R�خ���Y���&~)��l�n���X���A�"X����+�ſ�����w�O��O:m�B��p���F��n�r�b)ȹR��_�}�Y�:Iԫ͵�"��Ydb��b��/�D��%v������S��d�	B�����3�AT����h3�2Y:�ml))a�{݁��J�B��iT��ͭ��h@v���t���=[��vr{���93�	U�d�
��b>��Y����YiB�Lb`T�f�7�d�,�́�:�%3��(X*z�"���L�oQ�S��)�v���I�d����A99�1�<b�J-_�t[*N�N�N�-��$��e-m�l�>�[��JyFk�0��ң�lH�B�aK|���v!�/�3,���6x�����	�+�m�'�S"��
˶���� +�%�t��.[�S���b��-��3k��,yHL�u(��K�K��u��^�ӱ�Q�'�Z�P22g�Fz�~�\a����:i4P�|� �b����H�,Y�)�j�9���d�I0s�L�i��BO���$�M7���kKh����aj(Y���r}8D�8���0��ᑊ~�Uo���f���Z�޽{���c' �z���6�IJ��B's!a�p�*����'?����,������>��n+��]���\��\&~�7o^�Q _V��%��Ń�#�Ƥw��P��$r���h4�A�+U����`��ޙ�+J��>f\�*�:k�Qg��(�=:|���9����w1J������������*�*E,N<<I���-3V#�y�fˀX-�P�Ĭj��y����b�~,�Y�����k�)�ZU#D�K��g}�����o��6ˑfУ��q�+�움=J�����eU�8�b���!�ݛ�(��$�scM�W�F$aWbr��:C](���{���ÀG��֮d�DU(R���<G1ݎΉl���ŌZ;B�]u�"�ҫօ�2pO'gv����i��$#������������/�����w�f��V�j��[��ݼyS��$ZcەM���I]�¢�?�/*�f|�i"T�H�nSMbeԡ�]A�8N�>�`��-7V)��>�XBܪk	�ĥN�������Z�������:ZT$g�:
�ESKG��5%��-�KL��@�N�3��wV�HM��1���O)#9�c��sYeX�f0�-�~���S+V�^�U8q��H8(҉���
�d��E<J�H�����|�T写e/'�5ŔҾ&�`<Q���s1i�I���`a!yU���KV��#�C��f�4Q���b�}�<H�FBFyT!��UZ�A�Grha�\�{��]��E�HiI
��M�֭�H`�i���pe�rc����]29W�'*��x.�c�+՚�.uJ�1W����\)��Z�����+h���W��O�`W�cu5�^���n
a5�4��?�J�5M�i����RQ&�&}ͯj�j��|V�U�ö5�T�/���G��f�#���3_VU����UKRP$�r2��?�c���駟�b�7�`��O~���~�
6�֔���ALF�~��F���.���l2���lo���Ѓ�
�F.Bf��t�
��\'񯴳&50n&	�ڍc�=a\��t�ۛ,x�c�߹s�G9�����/�-��/��f�X��c���Ex������j��G'`BЬ�,n�D�}���c��u:�������[V-���-Whd�f�+�.��U)���El�2��6�c�"��Z�+����� �ܢ� G����TМ��1 �R�ʶ�8�����.�����[glz9�5fU�L�67/�����N�H	�4��,r�OX��o��������i�W&~�����"K���)�t�&�T5��"��޽{�!�D<%�����cSJ;g�p<"��u��r��HT">��;�{���`�'DQ�<���X(#�<>9#1O���Z-V�
�!��+;�[�nJqb�CD8��b���2�q����a�䘮�$�c�7�*b֗�n��g�c�BQ�	�l����e����l���R��C���L'�?���z�y��-��劕|�P�E���QF��ĝ���j�.�$A�R���"����c|W{s�P.~ A���Q7��l6ٔ��iZ���b�P�#y���hr:��S�)TzS9Cz_-Pbg���cU'�B��l���R�F`�ȯl�^!z�pC�r����v�{�����
���D�yA�dv�łW���d��y�޵}����dt:p����[�F�÷��g8��|�4o���]L�k�'c�f'��3��K�^�@I���<e�G�X(�EIB\�;!1"�/]��l��u����C�*,8��m�(����ȓ�����#Z�����VH�h�[��?ߺ�˨�w�b�CW��cU��(U��RO����u�1�׫��)��D���c�",#�k��ƇAA��S�b��9�'9��5�I\,ت6�Q������ �}��㬑�b��|Mޜ�a�*H����F9J	^���� b�p}��W5Xs�#�X�d��}~>P���8��F��%<hޔ��ج�9�
�:j^�'�>�L@�y=X9�e`��R�`��Φ�a�lIN+���)FX���0����*�p@�(���zM*�rSZ�����$*תL*Z��6����3[��%c��D���jqL%k0SF	$c�j���E���m�p���/^��{a�E�z��NO[)'�� E��K�� �:��������#�-�
��<	�*���Hb�`�_�/X6a��F9=u<PX�f�˙��Hg��sH]�U�O�k��f�hF����w���٩��r�e?J�]!�o<(E�(̏n^����%٠���rrw�\��\���"Є�n]�ʉI�np��xh)/˙F��l��s�w��G�?�����h��8�p9W��]�p��h������X|.�	���F	����t�0��!b���qD�J��)Ya��>V�S<{��N��d@��H��e��UP�}2͙<Y���/��y��R �X3����i�5$�5.I�[�M^����4����j�Z�� �.��ݗ9��_�R)߸q��l!�dY�quU�:�6��Y����2���&�x��A�{�xzz�{ƒ���x��b9O�8�����F��E�Bng{s��Z}i�Bk�&�b�&VE�/}
 o���wߑ�νn��Ø���]Qq4k�4��1u�S/�Q���9��Z��@��V{8���(�e��8Bry�"4�	<����l�[�
���	:���wL�1��ږ��]${�ۢ�{��%�������P3�;MTl���d�\��}O�&>"P&Ѩ��	g$�k�G���2���%ViP���������(��Tc+RF^���X�0�c�A�S�SI���M�(��f/||��S.���k�s<;,�ox�8��)lo51;�MҦ�ٙ�td�cO�Άc1�j9�y�����式�Z晧"<������mߌ��4�Ux1��"���C�H��Y1�L�yk�[�+d��"�A�svr�=�k�~�=S��<l��L:��s�	˃��d>���cw����C\YA ��v��B{ͱ�Q�C�u��bwgkň�l��ݪ7�V�c����i�6]4 �n67����U�/�1�r|��ePI3��Jc8�L/[���;[[7��c�o��݋�Ph�fqq�`� D�xZWK.�X�5u��6_.������'g���˛7�s��NG��lv6f�i�V�����I������Q�v�v��%�VA�RFl���g�����gGT:�⾨��t����I*�$�d��}��8����ӧ0[p��ga{���ņ38}�R�v�#"[�e.�RŬ���;���./�@�?X�wnR=m6eN~k�\�Իo�����t��3Sl>�|�.&S7$�?0H�[E��jS���ӱ�~��>�q����7��tQ��HY�1�G��2񵹉/�J%��ζ��T��*3�/2]��	��A�~��$��>|
a>����� ���;w�E������؜S�`b���R��r[�}2p�����<v���p��s�1y�z��D���MA|��?�����S�DG����g|�zJ�&��ݕ�>g�+Z`��|�Z�Q��c�(..Bb�y�YvA�-	?ǂ0�YjhJ���(fSb�;�|jՆh��k��ǃc�|��|H@��`=�л��J�*(��]ʄ�P��k0�;�Q��PRA��sU�g��H�o������U�R�NVܞ����8���g��R-a-�±���C��f&��p6,'��0<��_,m&�"�0�0S�jY���dzΊAIBq/��Q�^�n>2&iݛ
9��Xщ&K���������Gd���.t��uf[�5$|P�_K��1��id*�zq��?p����B7�i���,����O�<Y�><��ŋ��ŧ�$��x**�T]v0�Უ��������>W��0{ts/ָb���U�T�	���#��hbEb+v�=�/�Y��kg�U�흆r[�tϔ�V˳9�םv�2���<�J΋e[�®�u�Ɗ�rd=eW���g*k�� �<(��ˑ7�6�&.�g.e��k��[m��|8�̧�F�6<�Sq���Sc �ӱ*��ͱ��sM��FY]i�ͭ��wh�:����L�l �E�gg��Rag��#,��u��U�
����XX!��`��{p����)�~goC�h�����6Ѩp`�}��(�t��v��g?��|#s�NTq�a��m�`�����A�76j�6���[gT_X��y��V�� ��zM�gq0���h<ԉ-PVL,�X�V g�<� n�v�+�$�6�(J�!v)�j�QR\�dT��'�0�Ӥ�I�~WQ��c��`<�S.lnu���h��{�>>%���9�����j����{��h�D��
�%��	�],&ggU�˕��ژ7n\��ŬE1-`�f���Y�R���QX�"'�D��;�R���!ݵ���w���Z��Xr�p��4%�I�6U+��t���֬ɋBXH��ɉ 5�o�GiQ��9E?�N����4����7�I�'vz�H���Q�TvM�I�[�ZY�<��/��/x��q�m^.w��L���˷L������h2�=~Y ��8����9��|<y�/n��Ԗ��������;y-������9LF�z�s���޽{���(9����7���ݹAr�d��䭺�3�UU���H�7Zmm@J��R���n��L3��ė~�Z� :Y�A��"/��%�
#̊ZvY��9��)0�!��v����{E��7uelAt���̢�^�T�R����|�b­YS�R"�j^X�8�r�H��a$�.�Q�;;������oܸ��P�C��h��Wl�加F|����T�Q�F C�����~������l��2��
�+֯��mU��:5��b���������˗l�����bs�%�����f{F;���%�$ܘZ�ea���r�\��W��n���=Ý����lE%���tM��gA��R�6Ҽ/$>�Q���%�CM�e�8#£"w��'D�8R�����jv����e�n1"�&�# ����j
m�|��~��,u���J�-�����-8��2m:��/	��D7A�  ��IDATx�^e�$f'�P���BDU�����C����A(,��ڏ�V{���S���f���:��~u�Ȼ����fWf������1S�VCԓ!��2ci9��v����������n�T\��D��Pb+�U�1���R�����ŨUE'A�\T%���<�����1. ��~ �ڪd���,����Ĕ��"$P0���z�kr� {Ss������/#9�����q�SNx�4����u���α��*I)�ɮ�o��l�������!�&�]Ɛm�
��[gV��	;����Uk����S�8I3?��x�/^R��L����&(��ˀ��q����fX,�p{�b�)�R.�<9��O�vj0k�h+Ȍ&�;��U�
���L�v���{����rK�<B���Q�f�*%
;	gq�E'i>�?�E���ngQ�]�| c�ă~��=c0;'���[��^�6��݌���V'v���Z�Fн<,a
�`M(ʦ��N�Z���F�ɼ�`T*Vnߺ���K؝��{�v>9rRM(���=���i�0���V�������YO�Me�	=8����Ag�_Ja���ZS^�ui"�D�����((CӃ���i�	 ���8�$�dl��-~�!5��huK(Y$f���AN's��*ks����;&{El}��,���bV��Z�޿f?Ž�9��!=���>~�83�V���#�5��>|���D���PY�5����5��uQ��;F����^����g��͵4J����GV,`4�vv�8ѹ�,LjK�iač;��� ܀��B�ԛy��r%X�(�M�\���?
qs�O��و77�1����Uĩ/W�p2[�BB�g��N)���~�2M��r��p�Z�ɘO����G'G�[��,�q�vo�^p�L��n��������=NƦk]�s�"FK���\(nv:�T������d���؛��w�l5L��/��b�(>G�0w���b���ٶ�bw�M{Ě��p��Q&
��,P��q���%9?��(�R,'j�P�C��AO΃Ƥk��0Ùq�})!Ly�����
8[݂G�e�M�Y���z$����3�j�_0X�t=ѩu�������Q�T\󢟏���I>�r��X-p��l����E�H<zF�_��NA���s�����mu�sf�����`��ٱp����Z�b����%�L,[m���bMhrb����b�N��3#a/K��A�]�X�N��<���M!�
$S8��بs�?|������^O�^�{���_��Uw�Rƥ27&�{��+F����,���ˏ���e9O�*n��N�^���&O��h�ԑ� 6�e�'Q%�B�(������>y��P+�D�:e2��q'B��eVq@r�լ��X�+���B�Kƀ��jEǰR���à/�6Sw��}X��)�SֽE+.
��z"�ݶ�C�˶P���:��%�{���r}����Zʕ�b�kt���������*X��_�
C�
���Ph%K�eb]�I�>:f�ukg[�S�m���������$te9B�S��ϲG���4�jז��8譏�lD_Ғ��ʂ*_�Q��TD"�O�+�gǙ!$��"E� �&1����O����V#^j~"�ɴ[�W��c
���L�=swO ���D1*D(\���u�@P�r�Y�o\M,��Ʌ���o 3|���1��9w�u��89O�,�:�U��YI�����b�sҦ�E���"��6��zI_��	������]���5Q����ZwK�B蓡�"���Ə���p�?P̆��1�H���_�X״y�S[���j9_b�E�z���;���|9o���fE�B�4_�۪���uL�Z�	u.��ʐ:r?�&��Q"���_~���[���_�Llo��ͧ�|���e�f����t���jEH���nmmt�	����4��lo�Z�A�6�Z4���԰^�z��W_���+"�*i��|:�w���o����QA�p�0��sx��C�bXg7�2��}�`�?�}��g�����Ѣ�N�z*�1�U,z���}�&��i�TX����0J?��`I�#u���O�S�$*D��~�M]k˳�;D�M�g�T�bfo��*��?`�� ?T�5B�_������PE���*r�1" >t�X֎�O�U'��dC��ĩWb�	L"1�D%�Ȱ}:J���h0������~�8<��w҄�+��D�x���v�o�X��(ym�a0�$^���Z���G�A�ωK���'��{���F��%��ǰ�8�%�T����0��5�Z�^��r��,v��9Mc�'5�r�ڍ�Qa�b�x��R0�˰�#Y"D���L�Mf$!�����2��0���,�/f�O��~~�,��e:��~���>�#�g�Y7>�7VA8��㝝=���loo�	�(_��[z����I:�qob.Q���tLSC�G4;�A�P������e�qd�0\!�¹Ł��p �{��j�*��>d�ڰ`CF��~nA����6����S\��H��X �G�H����O��JՊ��;r�_.q�GI�3m��	+v��Gj�ro6����l~�-L�w<��:�M�&���2�*׀{;���.�Pk�aZ=L�c�	4¦��Mn�{��I�v�0�Z2����\��Nj�h���,��ɻR-�Y˘���~P�46ٟ��^瘉/����V�lN�xl��[7Rȳg��͛�l�xr�A2v��"n���߿��St�XZ*ȯW�+on�7��Nn���.N��n��K�&�4,s~NErlX�X���FxU_�5v�b:�|�2a��Q�"�� ���%�GM!j��}�sҏ>�H���p��Zu����si�\�"��\��� �
�^r*7���p>��"�V�@t�L>ZI?q7���έ�C	�i�����)��VT����,��Y���V���ke%�󾏣W�#�D\Ȇ�D\]C���7m���8K��!/�Φh�1p���lׁ�����g�^�W+ˇ!����!k��sZ��+�'#�4��<S���@�
�sYp��2�0�c�gh
��F�9��bNT��hR�w1_���ma�$�� ��cJ�*�a��R�gu��l�񽈹�A�����X�{O]�Z�J��$���]����쨢&���{��U\�k(�G�̊K��� ߸v���������T��������x��>��_%��u�*����` ��_�&,�լ�����f:ݵ_T�P����.�k�M�y�m�0��;'Y��q�֍e�bKF���ML;�!��&��$����Z4��`�]c��X�P�#��&cQ���vq�4ۍgϞ����Ợ0�C~�>�O���7�\po���Ѱ+� �P�/8pS��dN��~YϑBZ���ׯaa�/W�����r>-� {a8�yN��^�G��@ݸq���Jq�`gs;���8R�q�\ќ�VK��2X�}�!z��n�X�V�ƤJr!�����=ܓ��A"1���:M� �^��<K�h���Z�"U���jY�=%��͠�@��5##֜)&,S<O�>~��2���x�o��O~����U\�8T	�y��S���1_kK*��y�D�D��N���%e�ݹ�������3�[���A������������=�}�L�?�Va�1zʙ�9ǌ���~�X��U�OP���y)[��@U7Jb�Y�I4���G@ ^&�A�GǬ���z$3�3_~g��h�\��Z���,� n����o��r>�Y�.����_B:pѰ<f�%�n>��.b8��l&�� X,�3���S����5q���C��h�����?>99�,�W�lbZ�E 0��KdɃ5�����7�	�L��۽ݭm�t��re�\(\&�kF�_�����\"8m)�0�&Z��*�	Bb��s���A��X�T&���vQ\�OB�;a�tmW&��`���]��g_�	�&A����d~�|s�,<�S�¸�^d�2��J��/~�����\1T"��`Eb/�j���|S] A�CA�;����.~�b܊Ն��S�+D��x��@�j��k .��w�>|���S�Z�A�PX.����Aݻs?��U��_���m�s��8�'%Y1�;��淮��i3+=�T�1w..�{f�wus����xB'K2�'�.�	k�Nb�Z�T�i��b��x{��sM�2xa����v��uv�'�'�Zr o��-5�1�0]
0��r�E�$V�
��nK69�VVX�3�65���`�DGc���E+56��>2��������S�nܸ�#��;�s���櫯���M��>��W�N�������K�4��른M^q)����N�8f>-2���@B:U*5U��hϞ=g,e<B�����eCR�o˻�O��p�,0�GG�d�Y.D�º��|���kYD�RK���y��=Ɨ���f<�È��e���[|�0�Ϟ?a���m�\�X�]�iUHdPQQ�á���RI{�9 
�>�?%����	__9I:_��pYc~��ee�`�����=K4\�_qRuK��bS���$�'����t�~"w���0TlL�X!8�� �D�d��t�ay�,"B0���RTC���� u�q�w�w��|<�������ב/9'�^�7��kǢ%�T���Q:a���^�����OH!X���6]λJ�&&@������	v�[׳��ќ���&�6��s1�iH���B��v�"3�4X�kD���������J8��c��q*�-dL����4�&�S�����5���$u��&sh�˚X��Ɋ�C���Υ�8jի��9d�܏㇋0�oL�K���UO`��,	))��tП���"�c���\�%��睫lݠ�"�)�X�&ޛ���FȆG/V����7.5��ۛ��gs<v�����V��7�w7�hUϺ����]�mF�����W�TKX �Ū��"&���f�Q�Wo_�tZ�Z�gg���ځ9�N��ggj��ɿ�aiwj �9�b_�q\^��z�E�x@{�,���ɭ�ݗ�_�Ǥ1_NG�*,�Z���XS�[-���qx>�opLnݺ���wpp���~��{���Vo��t��N�#:/NF�$���f����S����g0:Ϟ=!E��l#�:>=�V�P�P��0s�ɍ'<ͼ��v��Bl��M��Q����U���^��0.?�������W
w~fET�fi\�U��9ej-c�n5��|��D�qۦJ{�_��%^6:=-�+"����d��`�pn��xX(�oݾ��n�mln�%t�ˢ4��na�;��h�e�-k��W��V��?uJs_>::f�~���9v�*��$��N.
���cH�J8e��r:�OgX9���|�Uf�9�5���xT�Q��Q'���v����>EP�t�*y��G��Z.5�B�:�L�2�i�چ_am�I�(,)�Jm������%(/Ct��7��ܧ�V�#�˔�ss�b�,���Ӊ��K� ���Ǆg��n��ͤI��nV����.aߟ���m�����3�ܬmv�Y�+�\�G�~�Uw����lc�K��0[,�eV_f�˒劬].~��^+�8�l��uo�/{��UH���O?������,����{�$���r��ò�0vk�f�����y󈊝f���dN���&�l���Po�K�?��d���@Y���wS߃͈�r��>
B|��1�&���y���ʹ�"r��/�'S��[���ϟ��y�����[(7�&X�ªK�@R��o���3(g.�����x|N�����Z��j^���U�Bh!.��S�����6�;�<v��r����^O�����a���`�����-Z-8�;;[*�R�Ѣu��y�N`|8���JO��`s����V(��h��@x;bQ��#6��յ.=_9��7:[�:�q�#Apxѕ�sz���ӸI�7#�l���sj��Q��������?���gc���JMp)	������A��f�Z���2�����qz�ۼ�_���E�gE"mLgrK����b�������E�(V!D�(���4
�N���I�qC��S����7��혧���W�iW�eI��،_ ��l%���3�`���6D�9�c]��ը�.qvVR9�j&7��R^�MbQ��v�����h"2s�K���a
̴i�N�_�m9���p�$&V-5J�.��<�v�)\g��ӵ��H��:(��D�V�	�XIcџD~��58(L𞞪 ���K*
!�ER�c���aB�cƱ�å�{�{��\.'�	�u�eW���4˯ZXH�L��q��*Za4�v�1;��#>���5�;U�2���߻w�ힾ������
�V�sκU@9U.V�S�Q,Ğ㹍V�|8�ᣒ��B4j�:ֲ/ޘR�$���U�i#��&3rh�����,�3���<@ι ��5��ģ|���Mx�jJ
Ѿܺ��H"�	Q�E�m������i��$� ǎ5زJ��:/�&&q�6����S>��d�4��r15�g�`�(��S��6CNY�`Z��wU�"��zvL�.����H�,��Ō����W�R���BA��y?�)Է�"�%���x��
-J=�L��`�S'�R�bL�[��J�l��:m%�������>���'����د�������x0bj�?cA�P7g�MKq�����i\�x�~��a�򄌜�\���`�c*�)~#KQ.��.�gU�8�X�c�e�A3�ĝ�}����8elp[xE���5�[�/���:�$(��"N7��נ���	���&(�.\�����=���N���a3�u3���9.J���R���*w)%Uo6��#S]^k��e�Q��v<fb��d�t���fn��Ƙ�Ղ��4��?c��`��L�!��5�l:��Q��&��^7_�&�r��f�jS<1}\��z3��41o\o����������m��5n��������0b���o*�-�7��$��Q�s�U�%8�͂�o*�E!�+jFH�x5��-,6�R�X���MS���7��߬�8�/jw��I?���j�2;�:�\-��p:9�u�Ōof����*M�|T�
�G���>���O{�� ���T�7�ґ���ll�q{$�V�z�L4���z)�sJt#����b�-weǆ v*�;d���=6a�-�nȅ'T�fsɎ�F�"'3��4�o��*x��"��Y��1��=������}���E��d[��{{F$f��bw����b�A��a 	�JX��+�X6��gx��9ω�3�sD!q�{_���Gt��0�0�񯤘�R�F��mBƚd1��k��(�P��/�&����]��h$Ouzɶo��k.�Eث%<�@��HQώ1lui̭�C�펒r�<� <���n��ģc6��}IoB;[U��?�̕{�X�}���'���<��P��LM���rw��E0x��C�|(�^�2��G���m�,EX�*��`���[�W�^�?bO��PtM��,�Y�	��c��78CQ)\���Ql����SX�m`�Z��	;�������N�ұHV�\q+��I��99F����"�K��K��'���>�ފ
A�+�_�"��y>����D��N-�	�d�&WR��F�z��T�y<� ���'O���2��6���I�.,y#$�ڹ�H��+2-�4� �Lȉ�Mvƀ���UT�Ƚ�m����Ã�~��Vӝ΍��3�乎
qT<���&=z�)�DE�Lf���B�I�h�5CC�{�x ��o�����c!��E���+	9�J��!�n!�ZQ�H��?�P� �{�O�<���؜H\�;[rl"��r9��`k��//��1���%�����9n�xNV0œU�C�	a���a<+�}��/X�s�/����\���w����hTu�X�]�˕�����r5�7[�8LEZ=��hR�5�N��m�G��/�uT���B�J؎0�U�3s�i���®�}�бu���>u��ڝ;�� |��%�s,DU�f�O86�� �ڥ=�)3�5�t>ۿ���'s����2ͳ����J�S�k�Vo5�0'/�.',�I-��|r|�.�p�ݔ����h+��%������ؤ������_I҇�+�|��ho��X�>\3"�����$��x$��z��^Dj����Le�$Q��}ä�$zp���s�0�cމc���J�;�I��ƯU�w�G2��VJ�޻w_ղ��]���	d�bI��l0Au0��
,QI�V���%�Մ�
��D܇i���W���4���c*$X�2�J��d�r��BmE� ` P���1Q���m��b�
A�Z������ب�*RƄ��i"�?��ZW��4�`1�����2b�hcXa#��ZG6[#Z��Y�Tu2���L�Z�Ї3L�v��+��V;�&y�0����%���iϕ��R!����6�������e��h,���b6�?��?��������O����U=�ꎦ3�A*v�ɥ��h��Ό\DeK��Û�3�?��ĉ`�\�a��9����M!����{���k��L,��8-a�/sԿhou�w�^�ˎ�eHꄈ����g<�B
��gM�������|*����ߧ锥��$�rB#��dj~���`�
��g�䦛���ȯIJ��v+{%1���Q�W���]��1!�M�gY�Xx'5�ql�b�kzI/�z�����T�b�#t��%�
���B%���ۂt���`s���;!�&t�ZR���ނ���!�3bz9�M�d2��A
Br���w��:+��A2��r���$�XU� T����)� 7T�-�)ʑ@=D!� �y��c�:�З��4�d?��O2΂�pY�8i*�g]���zB"��*�7�XZ�_Y���\��J�"d�}��'�I�"X?
��Pl۸���υ�;��>�l@�Fy���:�ixn	K��n�E�q��ǀ[��g�`�N�	��S����HMpe(�H{��n!z���I�������h%,G2�D�C�"�	�����1�WRךq2W�>KA��d�����X�Lc"��M��8����k�q	+��۔�D��f��)
'�c�<(��Z��4�9�)$��<��.kmPǊ_^���������?����R@s�4'� o�o#X7�)��R	`�{�O��c��ֆG��"h�i���5���۷ �1<�QȐ���/�"��!-�O>�dC�&�_�*���t��0,�p2J������J(��~��-��4��.��e����u��d�xUq4f#�U�s��O��{c⸸ם��"��p��X�j�2�I
�{b�jՂ-���>��w�o��H�r�f�TB~�,�D��-�j�c* 2&����6%������z]�F��'�⶘{��8���^��Jw�WN��{p8
i���������%��\e��Շ���l:�Ϛ��NVq�IN9�liCj������q5<��2��2��e�~�-��a$�>��"]�@
��R2�x9����U�U�Kt�b>���$�N�L�d�z�����A����V��1�$�=��B�w~����;�n�+ls�Ǒdg�3O�o��=�Ԃ���h9� �A6A!$ܭb9�L�����d.�
Ax���_��� dЋ/`K��@�
�I�ѣ�|����,��hT�<zd�H|q~���i����]-�t=�5R��W,0"�X�,YUs�Z���sڡ��6����Q-˕� !��F	���h�^ʾS�����t��dN8~�葨t���'�)���p+�Mp0F�f��p����*�|����^ `:R�ͳdeX�U�H02fVǞ��㊳�(fS��r����'��T�S��Vt�\-.��A���%�xG�_,p�Z�W`qk�,Bn�@�<��Ck�$Eh뵪bb�&|���?|t��ݱN�@�x���6M�a�^���i����n(����}�z�������vv�s�
�&�9�W-W�U ����w�={6�^���l}p���;���>�$�<�Wdi�U���Ð�h���Ě}��˷�0��m����8�P6��$�LX�Ƞ�L᷐A
�
X,�����ƺmXn�w*�r�?Q�Ql5YTyf���B��?�D�������-ؘ���F�xxx;S!�j���3���X����6�1ԃa�ր���]���������r-�������ܖ�2���Lh�
;���H�d�ݓnP��g�kA*rq;H=՝(܌�b$�n�*l�ݘ�.,.����
��Nٔ�+�3���J��'�?J�=[O�|�9w�K̓��D{�㩪��
A$��-�&D�ax��i)�1���������k�t���v�u�5��������L2HrW���`��@�H\��1*Xx��e�=��NX�����Z>�GLP��Ė[ZOߖ����v1
C�a�G�/��BM�q��ea������k��| �Ϯ�T� �Mm����[����ӧʟr=���zX.�r"k�(��λ��P�	%̄4�y�AO����D}����N�t�(C7��I��!�x&���".�W��rC����"V$�����&_.to�_'}�9�#P_�a�^f���sz�v��d�|��z���a�
~`�:�������fK��7oް�RT�Cx*�̒�<b
k����32ǻ�ѱX�"�VJM�I�'Ă��V�a� Ha���`Jc�޿?�N=lb��SR�I֬�n�cط{%2�bw�low����ԃ��Eb4�:N���"�0����h<ɖ�a�zcg���h���:�:_%�ob:w)��Q�[����s(��f\ai�Y�����&��(&��D��ޤ�C�'��L��MX
L���l�\Ff��z`	>����dP���$w����R��l�lH��N�­�����8�I�����+�H+���܂f�ݨ��#��P���(,�ӳc�4E�b6�l�S����G`b�h�ET���s�R��Jʗ2�x8Բai��j�T#;/I���k&8����-<x����`hsa��[qEŠ�W+%��3�����I�x�z��_���p���6-�:�ׁ�\%kk�\\^�<�cP ���UӷO����������_H[�2V���#�V=�9��bş��4�g��s����VC���*^�v�Ow8�;� U!�a!������R`h_��ˋal�9%��M�C|,�<��*�"�� xj��ɰ�Aq[V$/;�%�i�el�0?�߽�x�^P��-��")3���Xx�Q�w��.�n3g��,��j����*���׽��^�u��9i����rvCT *��~��X7NF��89;�ӵ3��b����d<e�밀78�<�UN�<z����"�ʽ��Zk��Ks���&�����p���u��3*���U����!�8���>v�x۠a˙��NƄ8�T��&��(��o��F�c�u6�{r��j�k
;֔zE	�k�����]���"��-�I�(c*;�f5`��G�Ʈ�o�ބ0����t%���n����o��RJ2�1v�j��������~��@��i���IZ����J0��P�Re���CQ���+NT�(?�T�n�ҡ�wV�|d��"���<����7*�H �9�p���tC�Z'��˗�Q_i|M���=[�ဘ��۲�� X#�+�쓼�-��v��q�M'k�&�Q��Z�:^m��p,a�}��K:KC��Uz�#��ِg�=���*�&&:I;[9%�LH�p��]�1��+�_C��*I�/N*�W�,[�hEpA�i�x-U�iƦ���Q�C(�t+���B�%�xI��8�L`�v̒h��-
e�.B�;�$���V
Ah%1Ja��+�Y6�~a2qǱ͆:�_\0���D���L��˨G^�)*9K����{���d�t:~�q�F]ڡ���5� ��C���bm���%��ƅ�S�V<T���A�.�R#@+^)J�?	X��24�$& Ck;�Ysy��a��1rho6�*zd�z|���<c'S�+ղ�t�C��������1[!!�^������u���\�R`5M��?~̑[=6v8+r�L��2��+aʔpp�ɓ'�-b�1��~oO�A���_�%�-"���:E, >0]-!��3�?��C2,��/����g��L���qR�Sʬ��*E(lY���I������v�vvU�2��VF�@S�J6r	�(�A�����i�,�U�ݫ5�i��S�����F��r6���Y��n��`�˦���U
'Y%^	��n'֮
����y�f���g���b6Ʀ,GaΌ���h�I�5����wp������q?��!��e��['��w�P&K�Ԇ�w�'�������pg�*\����|>_�szr>O)d�����-�=�%�̈�J��J�V�-qK�C�8VX��&O�b
���������a?�[�_�$��s��}�� ���9��$�TBD��b8p�7:	�u�L$E�eK�7G$��ΗVȒ)e�.��2�����[4LI`ňħ$��b:��Zb�ybq	��P���YT���ad��ʌ������T��D�0�d�`��
?O1>��|P�Vj���1����|(��ZNǨ�0�7o^��_�j.�A�Xpx
�PH_��A�|Bp�3���$��VdF.�0ܳ�d��iZM	~���yx��2U�a�Cc�ǹJB90&�3�\��� �yl�9��x�f]W��ݬK�H���BT�u�i9=���;�skee1�12��(�LY���j.\��a��6�i�Lf�1J9�c���MP�Ϛ�x��"WN{��n�6�/�J�[��U���-�T����w[[,$��G^�e�����m�{7�O�U��d)�L�ňuK%3Yf3���vHD�*U!i�9�T+�^�\&�Z��x��m�V���aۑix<��AD}����&��j5�ۃ���M� B�i;���~FQu���}��By\���{;[�+�j�
�cC����]I�B7z`�P<W�&̯)�����������D�؄��	㛲��I�,�A?�9���!3��L�YJR�Y[�6��N�`-Y����1'P$ز�D� |�8�l��������1Zև@��fy�D��f��}�K�l/j�T��Z�nt�~!����dd��!��c�Eo�=���g��i��aI����Y`9��5;�'�S��TP☡�r0F�֎�+b���k�t�,nFl�����Q��mPF%�8��?�u��c{س�1�2zk�01;e�d�T�Z0B\��xd��S�D�܈�Ņ%l���(̍�H!�T�@�X����T�LK�o:GR��5�U�Efna+�����k�U`Su�Z,O$ɭ�}�A���)ł��t��Z �mx�b��W�DR@bB�D���P+v���4��j�\��(wRL��}'܎�s
Q2�U-��O�-G,����>PA������Xqr
�(Дꡄ?�T�ݰ"����Tzch���_
��;�=R�2��@V	ܵ����.���2�1A��>Ƈ��aj��<��M�/�,0UȪzIn��&)����_�V���7)�%fX�L�������j�KC˥��ي�k<��%A�*U���ĺ��;t*W�*��Ę�ۣ���1Ff��V�	��a��:�S�YX�>�$�T(�'���AQ.�=��%o��Z�2?���	��l�ل5t2ͧn����(��Q��q"�ݪ7��jf����p�UL���b�V����{�2��O߾�mw����f	* b_q�F�اsj���P(>~�1�$�����Ζ��M��jM����F��������o������?��?����;�m�z�N&�R�,����g����{����3�F4	�T���s>7,�o��C��<I�8�K�]�0�AE��l���ϵ��Є�&��(�*�K\,w�܁�vusd́i̺�r&�� ���ʻ�ͻ�����.��_���,ɝ���U}�������M'<B��P�:ɂ�Q�ѨbrօN�r�o/K�Fb�Q*�4-&���������:���+���+��is��T'`n~�f����kFD6�:Rx㪞�ie��f�8��η.IShq���0�C�`Ŵ�b���nެW�ZeS�ǠMN�M�g�%RK+��p�1	�����}��)]�z}a؁�V��=�s�cu�N��L�{��	��R�N'3Hp�2���o�����j�v��}�"�^���"<�e�H]o�Z�;9.Y9���4
��Bk��lT�y���F�{>[���E�s����&�^���u�	�].�
�5��v�"����61��������lJ2b�6���̓%�I�Y��:p���X(;9��Z�q��K�:-�h��O~
���B���6VG2�t̙wR:��j]�
1���l>���܆�Es'PH���"#�2RD5*kԱ�ieYe�b��9�'�8�l4V�oo3�/�����b�ׯ��x��"B�u�ݍ��7�II�1���|��\[3��0�U�-O�Ӫ�oKnU�� �|*
$b����>/^�u��FW����g]�nVA���2��A���Zd��,[Q[b;)V��&	���_^�����1Nu�*S&���b��q��Ђx��=���ڂ�`2Ð]
RM�J����:�U�5���TMO�Q.�L���{�|G>�(��g��w���q�sݔ%�R����/{ [Y~j��T]��]1����yP[<Q��Ml@Yc�	䦬�M�D�lmU5)���;;�޾a��N є�W�����'a�,����
�+��*�^�戬�(y9X�R��
�r�3n�vvz�cE�j�O�Ր�/��*B`oBO��td���0Fo�=�/�
3Dfé#�t�Mz�S5E���YA�U�m1�dˑf1�ˎ����C���U_R�����>@��*�I(Si�[�kd #�$Cj�(�6Ѻ	 )FJ�Z���Â�lC�um
��d�M�7��UNAH�V�g�+�ư��XݢkQ����$97��i��߮FW���[ #m��m+]V-G
Kl��?����ێ��xf�Z��cj��Y��L��tf_L�]��l|�@�]n��'�V�"���C��VB����?*����O���$�N'�k.hYm�s�ޥc�-�������t�<::
�z@q'��<}k�N"��JJ7�<��^sR)CK���5���$;=>�/�t� ����]BRt������N����Hl�����[�E��~x^x�x�����?�C��u�#X�j�����a�;pl�\���H?�{GD�����ju��eV��Q�<e��R�
;h��a"KEr��*�U���k}jя8	<�������BH"cċu���*NT���綉eQ�=_7m��Ba�^�����]1I>����
���N�~S�R	[�����Pq����X����|&nֺR���;;�������X�-8&���`(ЧhO�((�,���<�c���8Vq�Ț�bOr�7Dkn�E�-������'��, ,D��%>�4k��� �X�f���tv���-`�G�{v���a��ܓ��%����ׯ�����q����A~��>���� .sp ��"1t��z�k��Z�Sx��=`�`7\^��v��]	�R ������1��^�����ѭ�~���X%���N�	JS#sr���ң�!h�.{�R)���l6�	�]ī<���3���׻8��!��Q�=�SN�>�jrC�6[-�w1g��z�u�[�mC�@�AG�0���ۇ|� 糐%�|��~�9��P���P����RD���e�p��SHWs���d͉�/��"n�S5��xt��M��֓���D�?�hg3�U��6ܲ?`9��֨���w�Q��;F(C(�z<BKy9�Tu��j�a������s���2PU'���ҭ�o��"�T^�3Ͼ��Rak��;�*��7��l�U{9♑}��X��khȊb��f�1��e�����*�5B�X�"'�qŲq���o�����-�B�)�7o�@��˛ HīP�!�`H�c!gִ��S(	���;`'ꀇ
�d|q!�>N�W_}%	 .yl��f��l�RpYs��͝-q��I�n4�2�5u�H�HYa�[(�e��2�$50��p�:���+�:I#V:D�%�+�^9���Of�k0��q%�e�(��qU�j�L����3�~��:7��j�
��I`��7ݲ�I�1e���Fl��rnRcB��~��_~���Ź��.�
��n���?��H�7��R�~������}؜j>�#�J��l<U�]@�$m]��?��?.3�k��KZ`&aѿ�>�g�4ԅ��f�F�s- �����ͱĘ�q�8��a9�D�K�4���r�,8�M.(D�2+B�%�]��`�o���䚶�1f���s"cK�������@;b���[� #Y�)�T�n贴�v�;`4 -c��.P�[�P,a82�g�=Q�X�h��6}�l���)��bq�q�b����qS	SZ���QRc��2��$�ɿt�۾���9Y�\H���\������*�"�	=��͕ﱫ��{���?;~�C�\������%&��Z N	$	 $Yz�u��Ǔ� �%��{�_-O�>�C�^X�,��F�J���p�������:�-�ñ�c�Ve+��<��95��s[�w����z�^mVG�^F�R�H�b��/g�p��H`��Skv��G��g�ܹ�7�q�>�s�����x���bbA�/.�E�Ņ���
Kmq,�A�L&aT��%��d��ŋ����X��j�r��Ad�(�K���:/'�G0�:{[�+�������	�'�m�9��G�i�wޟCA���2.��-YƂ\^\$YPot�w�=
�q����LW��n��?�:����+R�
ͧ�	��**۝�O>�Tds+Yj�nuv������(k	�^���wq���=�p���@�¶t�$��;˻"���~/*208
����h���)U�S��=�`�p��Z�m�Y�O&�_(AB�ԛ�/�1I}k�6Z�r?%�i��|q1�e{��ܩ~J�A����yN�Q��;�j�a1��:���fql`3�!�4ػ�C/p�����U[@��*L����)�e�h�n�\�.ptq�../��g�E����"�_��ѧ�Jr��i��e���ϱQ0��h�;A��>�O��;7�^�;^�i�����.O|s��w˵�����t���KSck��s+�9Ղ�1�:���i���'�)PKИ����1]F��U�\)Wki��M�@��+.m��J\]��R��n�Z*C?Ȱ-��R*U�--W���Z�6Z���W� ̧�e�t���<�Y.���i�[)L����9�<�X�Aag�To@���06�|�K�&��7 0�V!.�������_��_�;\�菰�Ƴ)>|��	S�y�(U&I��G�x�H���G��C�G�'��<���ݝ���D�¥��d^�?zV��r{ ~*&&Q�ـQ�)�%�
����ł�v�*�8����Z��m��{CްA1�	s�+Og�$M�*`��5>zw�B?���D�H1��kdME���f�NI���or 8������+ڀ�I�	%I�����5��$d���y)��ӕ1<K\�Bs�*�_��׏?���hm��@�N��:��z��I,���\7��3�Ռ���'�
#BPLm�U��`(������f{��S��P�3��rc�]����BFVe脓�eH����vS	.����˗P�4U꿸nň[+�����j��7��ϖ�.E'T@ \��o�u3V��D(�[����
AԐš=�+� ��w��'���k���8��.��If8��'L�j̮�|�}`��qyգ>�qף+��V>�))"�V緿���%�^l|m�)�P.�Q�2,\hzQ �s\��&�lZV(D�$s�,9��O̈�*�3�Hj�D�Yg�4�9�ge�6��@����'� a���n�/��/ޟ�Zxm�W�W�)�P0�ֈ���?R��/>�j��˅i��ϔې��a��ri j�5������H�9%G�����^����4����><�soC�:�UF���-����Ϟ�''*�R�F�I�7&c�sa��E��˪�
K��~��.������j��(�1�tacb�=E �ݣ���`۱���EE�朞���6�n<�X�$"61	8�Z���x�W�������L�@� l򃝖W�@9�E���0�*>��-�K,��S���^`m��F�E����_b4m2��b�A��{;�sk+�M!P�!�(�@���r8].6ʺ�
,�b���e�:�N��w����t4��;��^�	�{p����ۡ�
����{���	�,V�+��b-����T*��$|���s�s���k,�YلD���woc~��O?���o�a-^{k{kgW��,��	�_,3a�*b(>�r��M�:y�T#�eD��3�������n����|����K�i��)Վ�Z���i�h�S�O�A'�%�z�g�;���~Z|`.l�"3댭Kf�X�z	?���g�U��`;�E��%�@і��b��:�\�c9dX�UL~�O����~�&>������WJq�Mf��#��X*C��窶c�;w��v��^8�w��V�:OD3>5��~���}^+�u	15����h�ۮ��a�W�D�����F�&����mñ��_~�b������IvK���G�������0��}�ݳ7���U�dQ/���dAC2p�rψ'����A?
����|�����;����/��.��_����������Rt�e�u'u�Aya1O��������<�$��<� %R�i'5*v�(�_uf
�dF�X$�P�{*vtvP���z��JXh�I(+����:��F�<CaQ��lG�2���l���)���)�R���Њ���<41���6C��O��tL4|]� (�{��͒�ۇر�߾���8>q���͠u�$��28U���L�h6eK����n� ws�a�Q�-�ؖ=d���%������0��������j��ݿbZ(��,&�%tׄO�\@G歕w�2F�\���E�-Ed�o%�>��4Ƃ��v�Р�������2�o�~����ٹ����Ψ1�{c�5*ݼ���7��jLN���j/ ��m���I�3�A�C�`Q?x��7����.!����R�61�����{I�������j�����o�5�a.I���K�����2R[Ғ��5Á���]^��ɧJ��dȾ��NS�[vZ[��6\�*P�31~o�^�_ȃQ�Z���4^�x�D�l&.&I�di�͖c�32Jݘ����,�&�?�H���� _9��z��E�!�M������@歲xlB��E:�x.���!�r�x�~�&���X�*��V�W�o��*K��{��,Is����U����#�1����r*��ު&1.2B$}k��Zی�U��|�1�A���~�y.��#+�g�Ջ��lRJ̺C�\�����.����d'�1ށ��k}�@L��˳K%�D(@*�9���*�Wsr�[��8���H2������0v�f�{]ƺ;�-�{?�š��j����Ö��\\���P��R���(����{�WW\�1D��&7I����R�0��	/��'�a��Y���ȹ��5ǝ#�bf(�+����8��+�{$)�Ig{�e��w���D]��	G���Qe����hP|�%�^*�����U�=��_�"��ta�>Ka%t3��������)��?bV�Qw,+�� 1��7�VDϗV�E�nF츹(��F!/K��"��A���ɷ����i���bn��#p�ؙ�Z�р�����(��q�'��Ïf��������^����d�r��bN-�:a�٣|:�֠����c�8�t\����ܪ�WK�2�u�UKKҸ�l��ga�٘��g�=�:����������"tg��|�G����,m���~�poWR´?��7�����g�u��?>��[�nag������;���d��/Gcu?U���ߖ��Z�1��d�Ҋ_hwo����9 þj�čZ�sf:�������(�k��(Y�C��M����e�������tg� V��f�� ��s�<P� �h(��V���x����O�p3^��}���F���dg�2%X�I��	�I�نԇϑ�乲̰���kt�5ڸ;��Ւ�UvvR�I����?���p��u��7S�fs��l昛+��������Q߾;���A�\3}3��8{���\#!�X��ҍ�:�W.Tn�H|cH�{�\dqհK5Y�Tatc-������>�-��n��3�$f������!5����/.���D��*���y�����c�˷��rw{}8�x���7�B�&˝;�¤��9�m��Y�����=`N����9�&�Yƞ�F�6(�d�28�V2�Kj�\Cߓ;�G&�w�Y�RW�;�f�DJ���r��1S<g���é$�0)i�G�i�,���;@���`3���ω�j�[{��q�X.���0�l?6��d��*��
rD��Ud��@F����:���z$q;>eRˏ�@`�b %�<i�^��&�zt��x�el�k�tK3Z��($p��˖G[۴�Vˑ���)r�;���$�U��&r���^�	CeR�������Vѻj�Uk�g�ֱP���㊣����V�����w`>��_�;����.������0��Z�kJĮ�XK����쌳�����<}��,�"�69�8�j�!�JycΐV)4�mɪՁcxx��?����(
�m�|d̊C�7���*ЎD�r�N����+����bs����:>U�?i�[�z1<���Zx"RJL�n�:#�:B9��<��ڴ-����%���La\UDcz!=U�l��`�
��*��y+�V\�K��`��ًv����Ȫ�PVf>-�c���.*�\��QGϚ��V�0�f�^I��M+W��/�z����߉_�3.�؊(�������G��:NbV1�_d`�t���uO/�E��8%B�c�x���+�}Y��v�k��O{�/�h�s�j1]
q�����0���ײ/]�m.�����xM���� c��O=&��&�'"�[��ѝ�)��$T�f�u��.�ʞ�pL�P��z�Yj�Ѥ� ���k�w���g���)O�Y���ɓ'Jxjqɰm�H��`��J2(CN*��ѣ���WI�8�T�Z&/��ĤI��r����Y>�l<��[�uo�1��� ��B�1��*�朢� ���h��݅��4 �"�����x�bE���������Ll�<�)͓F��>A��&��-V���A�Y��Q)�b�Dnp���x�x�|�48�����\)%H�����4�J�/��ג�0f��|f��F�Ν{��wLQ��� �˺�36�hÊ���ywr���D�V��=	�3�
����*I��j��q�-o1�,h��ǟf��r�$q�����fey��ɶ�
�ɻ�.&�-ܬhQ�AEp�ϰ���[�P�&k^z�YhK�����Z�sYU�u3��k(��b����7X�4�F�R�r���(�!��wwTC
Y&a��
v(Y��H/�O��<�u���45�,ntx�.e�벚�Ǟ1�������wO�2�kE��U�2�U��j���'TAT�i��ù3� ��JੰG�t��$Fu��}8�o^�#擩?�w03��Q��	�Zmh�EJuK��V�XI3/�ha����')�����s��8�|�=�������*Y
?+)h<M�rٻ��H(-�;a�2V�i��z��}EB��q�P��xH:�Xy.7}����J�ܣ��ڨ���;#g4��?9�T��=�Xi}X􋌪�g�0��vv���U���3&Ϭ)�F�ZF,L@���c��YI &A��={*eϼ�j���!g'��DANz��4nY����U�S��J����ZN�x�����X�PY��pDY�>��H��/����|(�:?�^s�;�K�́����e:�6ܣ���=�>�2m��i �dm%i&;��D	L)"U3�&'������[���w�?�x���Oҋx��-�������{�"��J=��d�P�^���>#o�<��֚��3.��I2'1�������2t����&C:���H$K"��_!(1������`#���/�r�N��[�q}!��4VQ(>�:��=|�P)%��$z"��û�*�0,?�/�ˮj�����IpA�X]E�P4�E�yM��X7�-��6΍�X�� Q2�(Pշ��6�|���-��bqx�>�Z?GmA��K�������~���A���M��U
�;e�K��w%��?��˯�R��C��0ZA�l6�zz���=��!�>��oḴ�Q�ݻwtt�1�՞����ÓR�[q�T#;d��j,��a���nm������8��*���i�@��D%Q�F���!�j��٣p�h�r6N�(s�֔�{���X����E���&��,�Eh@y0��c)�-�����rI�B��ڶW�h�VBm�O0&pw�?^]i�r�l���:��ǩ��|���c��Z-xo�9��B�T}�c�Bah���J݈�M�v��u��_��,6b����U�B��*�i�&c+�V�ތ搷��Rn���~�V`�I��w���1�T�7ֻb�i��W����'?�i��b�R�����ܜ����(�5�r?��*b�Ȟqʅ&���t��,�G�&���a�-�*��ġ�p6%t���cJ6�ZCa
�e޼.$���]��?��������cG��n��VU�����N��+�(�]�i��H�?��,g��i6��`��0b�s{���$	`oX)G�e�/v<8��~��ʽ�������'�5@E=�?Զ��?���ꫯw����!���ke��O�0���U�S��r���[�-����~��j(;]*<�Q���HL�h�q�EkD�hυ��nS�~"\xh��b�3J�ɩ"�s��?ؕ:��WåBĬf��]^*@!;�3��b�� �u�&��@x)e��<�gm�k���C���h����'�띾?6&��dBt���FT�]�&�I�H+`5�.
�m�������o#ᤅ!�&��KT7\�%�~��U�W]ǟ�Y{�\������*��@��jU(M���|�P�İ?����rZ3��O���U.a�wX��Fk����d�ԋQq���^�\f�w�T�fMC0kQ@V�����8Q�^�ƈI�`��Vj:YX�p�T��ֲ���'?����w�`_U*{Q��ԑ�Tj�qbK�r�6�������|���]|�鏆�ѻw��d�*B�C�`+��<��+���0�0?�D�F�0�.�y���Sx[�<|�
`�[[��u�'み\-x"<ok��f�h4�0�*C�������ʬ8H�]�o�b<�1)�ս5O]�-[;�#����ަ�8��`Z:Y^)���4��旪����,�W4J<q|Xǰ�25k�b�"�"K�?�Tpkx�H��Mk�2?Sp�Ν;�F����)σ�*8���>l^�W�4�,�'�R$��7�y��l�M��/��7G�D������z7�r�*�N�g��%�4%�d�(���I-�F��ŅuͤAc֢�=�Ct�����d`�·��,6���_~��	�	.1�����/q�eh����س��fR�ב�.
uI��`>,� �x��Z��M|)�!���1��S�I����O�t�������"�ͬ�} ����LP�V�[s�PC�\Ƭ
�ȞN�������L�յ}�vG�[1O]��Q(l1��<S�*6t����ð���!ه�1�ƚ_D�i�����{���PJFl���,cJ�	�����#9�JEb�娩^��cb�(]w��x�t{}��ao�ƗJо���qb6��mň�m�߿ϋ�U�CH��d`9v��l ��+��^��ÖS�?�pfM\0H���e��qE�*�c��	��F>�=|��\��>�R������wϾ'�jn*_,dF(34�f&��I��K��9��Z2d�8��ہO�XgC9C�ru�R	��y���ց*���-���{ⵦV���Y�ݹ���T��%p��T9�ҙ�GZnf>e��l��R̭x6�c���0*���Yk/<�^��0X�(L*��v�hI���2t\�f�\-�X��tDq��`r�T�S��1E�m�	�|��&���g�'��!���݂���臞���%l�0��������w�K�Jpce5z�M>��l��ɵ8��pxa)��6�l=��nv�+��*�V��%�pu��-�f��6O�~ϰ�G��~�3�L�����{���Sa�"����Yh���;�T��0;M[�փ�d�+�Y�NP�	A�l�4���x���q�z�Em-C�x�iNs2���|#Xdp�AO4�DT/�471�=�k�ԛ8reX��W�{%�Ӏ��l��],��R'k�T���e�v�}d�1��� jG#��=�Y��t2����x4p�w���kؿ��gk�4�S�R&3�V"�ҏB��?Ǖ�55�ѐ��X�A��������B�
0��J=7�$�rF#�P�Ar)�s�R��������M�.���[�c��x^
mj���b��}�Mr.���HQ��jTk�)���������S	q_2�a:�w���LY����jR��	Ɗ���b�3����*M�Y�M��Z�lGGEy�1��o�H�,����y�61iO�?c�0�7�o%q�aDH�'+?T�#�{�V(V�EJ"q:_�h�L�����$`�{���.�oV�����n����Tl�Ԃ��Ji���f+N `Yᣋ[���S�zVSR)����?��B����Xn�1���;|���k\�:r}�|��f���l� wQ)����Zvy��F�<mb��������Y��h�1���;X}�KQ���@�� �Ƣo����L!�,2H�8K6,~�ط�5��i��~j̚yF;���� ��H0���������<n�_�uq��x)Pc�m,�2��Ѓ�{N�L��n����Dj-�@�J
o�>��C��>z���U�g.0��O�	d�3��j��$�ay�c����?ǽ^��^�ջR��,�S>cv�W@4�u�(ׁ�_�J�f��J;��8�feЉiu�T�"����)�g�cdU�lѩ�XI7Ԗ���"��ӧO�em��к4�ԣV%����Zvh��h��U���Ҟ��
���Kho��C�t�-{���1�f_��Q���/��b�l�Yb�q�X��ٳg�rwdI2jJ�d��a�/^�fDj*R�\�v�*DOӪP*��Bމ�C��L4�*�8���9i��s91�����K�\.T�+��Ks׽(�������m����X_�5������׺
n e�w���Ʒ�ܑ|by��B<V��V�,H��t̕f(E���v��29�2��~tt�(�^��Y��0�jǕ�B?P6^�P��c�ᅔu���i��d��I��2%���G:���[���SQ(�}]�2x�j�X��M!<�3��<G� �����t����핌@^���|Vy�1�(����j����4M��ψg��ew�p�
�:sXw�B�]wG�p7)\���ۄ�[�D9O�6�(՘� ��LXx�������ju-�P��(I�I�pAyk�$��u�$��6�u7o4G䝎�b��^k�u��}++���k�a|3-��j��Y�V�r*QCVh���������g��{{4$��{9�W[���"u����"0������0�� �X*����{��aqS=�r�'>��3a^A�z}'�c���.���_�Ű	�>;�b�� �?��O���	v��V'���]R5&S8��l��}�\���O��ݦ6�K8n���{���I�E��g���e�Í��@I<�=���$�b��9UI�)0hA�I�eS��$���W˒S8�p������$�Eww�!Ξ?^�L��0�EO�3��6j�tۨߟ��Ex�;dۙ\��[����L��2q���q��ae�����{���V�f�����Y�٩]��3�'�z+idщ,k��~������
�R�i�aǜ�������?���Wo��׿�{G�n�G�� jT�}n����>�l��|0�"���ˋ�7N`��g�nk�i5��M��f5��Q�i��x�����j���c�`)*1.�Y�In�ļ��H�`�iI�9&ĨڋL�����û��q���>���t4���do�`a��LT�8oQ���$.������c�dc�ǚ���%>�ϔ����^o`8������p�����,��!�K�yΪ�ǏCQ�_]£/0ɓ��\U�묩�릹��Q��&�V�R�ۿ���H��U�k��3U9aԨV�[�b�A	@��ٛUFG�ȵ�`+E��̀)t'1:��xW�����"�d��/y�Vd����o��A�.�V׺�R��+�<==���ci4Z�P�(��Rꁕ�$���A�c{�)0��txs:#��*q9�K��Ā���?��~��߲��aL��hȵH�9ξ�)�b�A~	Nf.!	WfS���2E�@M����f&�_��_� �Y��Op�Mos��:;o޼�T�(�?���$�o�1ӟNF&H� 19�d�2,��>�L�A	�Ǽ�c�nI�}*ꔫ��ӻw�e�_k��Ǩ\���Q$Z3빽��rL�F^��[�MQ�R5��!n
j�`$ٹ潑����Yp��Lf̤�;�H:��U�&�¨����"��u�j�r] i��n�hJm0�a�Fr����h	�[X��\Q	���z����90R<����"�)Z�=��n
�)#M�I�D�s�\���dĚ��K7w���S]汊��jd�B)ڠ"�\R�6*fS��_��R[{LZ�by�F�MD\��i���l=�zE�Lԩr�O*��P�c����0��|�wy��uʦ��R�jh&c"͊���� �\�hD��Ie+�������a�r��Th�l�
��=�s�.�$��׹��F.�4J%)�5�6S���՚��=�:�ii�1�<���-����l���N)�p���˹��S��RO�5V�l�5��h"�9_�F��ó��A��ȶkF"Rg��b��":>�	��El<Y�}�HcgGW��F�������kV}�w��ν<�ͺ�s���g�d������ng�EA��wز���F���L0X�Q6zk��/!�����e��{�7��,u��A��bp�v�
�`⛟��L�7X� E����K�0���4#�Yo�E��<�j]���U�R�ٕvowK���gg'S����˗��ի7�A��/D%�/��G&�wv�;K����/{0p�P�D�Ӥ����=�Bh�ք�v���R�u)�d��u����#$�	٬U�T��f��C�e��{D�C��I�l�9��v���3h&��H���rK�ioo��%��u�����z%E�D7���`�Wq��_gOC�v�Y-E5��5��e/�K�K�O��V��K]CA"��T������P&,]a��حa�-�/��3�.T)V+��ߞ�|�~�֭���[���z��r����7ϟ=�Nn=|�����j¨\��īd1���~��A���p��U&�։�(4��b1Q��{�6�����1VIgJz�c{f�q�`)�a�L�`Ϝ�H��ʥ�b�GiSm�gg-�-H�(�%+���R=m?S菆=�<�)�C�Y�r���[��r�4��al9��︣	7���r���.I�o�}[�N%����`�D�J)����d�f1	V�|3�#˭Z�ږ�NS��s��x��₹Cߏ���e׬��a�Gh��)d隇?Sᑌ$RjٞwMgVcoP����azh���Od>��&@j-�;��^�'��0n�$*k�Z�6����Z���р�U\�l2'���*��x�ss/��܂��ٺ܌�A3�������v�t2&UT�Md7-�'fC�y�(�K}!���!��H+t.79�nC�P�p5�f�����:�~�)[~�tطㄶ�ں������J���p|��i�:�w��c$�1̐�?����0�N��Ж�ݔZ��֩V�S���Ta7���V�����;~���"��Ěu��K&	"f3\Oa��pþ�+�C#n*R�`7D�Ĳ_�����?�hX]�j|x��eq���5�?T| P�J����:�rIK������S��IF%(��BpJG� �������&n1����M1�clx蛂u)���SC$������EVJ��lT됡�7�6�ߕ�^=Srev��4����]�6�\B�`3�	�þҡc���,W;?@����0fI\arAps|"�ɓ'�_�C��|��?��_��u�uT�f!���ı�!�]7y��t�!��^j��41�ˤ�4L�|�7+�#R������� ��ܵ�r�$�%&�msϺRvx�� �Ϯ���Z:�Ƣ ������au���T"�F��z��e�����0,��3R��{W��\�:��T9�T�2��n5G��ҚS�^�*S��ɴ^	"��i�vv.U��@S3�x;�����az�2:<��\�O�<�w����?��Yo�������)�V�����G58����j<��Nq����~�˟������"]�����Y�V��Z/L�&�����,9yw�iV�قx-D;��C��W���i���9��-w|W˥��{�ݫz�m�[��-��$�޼{�h�t~ry�����f�������}���۩��ʪ�3'=z"^�?|���w������.������7-��A��=,��[�#���0D��^b9K���{
^�o�;��iWk�Ѹ���/q��d't��ЅpC^��x���C0Zx�O�yo��׬�T�6e0x��"��;���ƪ�2�	",/��q+n��tz�V�r���7�u|��l�ƌ��!+�0u, � �����t��Y���d2�0ڝ�x2��Z�V��B|9���JVK���5��<����7[M���N;
ݝ���gO+e�B�N��C�ZAT�����x>���j9X�R��bZ��vw:�߼(���$N)Tu��l�/-�Y�*rVT���n:�W/��-���x�����H�Bi0�����zH�Z����z.7g)l�����TX�]����eb���2)��#��P�MH�R��Xΰ�̮3�����l�S�n6�vpZ�''��4o���b5�n��U|��޽{���
�S�>���6�b6zqJ�Z�,�E�J��Hn?
qL��R�.�TK��@�^�£3ȤS�2;;��<�S��Q���=���'�8Y�a9W�^�{�|{ow6��8�p���5JWK(�U�U�B���I��/\&q�V]&�����},+$p��|Q.�׭�G:�~���3��b���_С�
^�����V���+�*�V�
�B��p�^HL��Pb�i<�m��~�
�{��cw#n�񽻷����y�FBe'Kk�:iH��"�e�[WŷI�~���o��̤Rc��Y�.T���2�n�j��Yx�]U�L|>��h6���~�2�5��N�]��X�h��#,�j(V�U��{1\h5�bx��F���nw�P�"l��c�t�oc�v狡��جW=blF�J��ެ�z��R9�c�+�1�%�~�-�;�@X+��F�9T�@���'�c+?����!�W���� m��نEJ�x���K6�XAFW�y��e��,c� JɎ�lW,兰���CA���$�k�]�3"�f
�,;�H�Q_�2��u�)������������u!EX�T��YM[�ھ*�4_͕S�dcT�p����Ǐ1f1�I��LW��3v7�a�(�ӧOE��e�;��k@��(�9��o�Zt`�l �?��Ϻ=�a�BӴ�-$"[�îc�۞?���,!��t��tP�-|�����8Jo޼�\vpi�
��9� {�7������On��8���:㨀�M��[�ml��H�|
���V�ݰ�FGE����kF"*��k>\��j�"���BQ�$����-h)��`����"��e��_��SI9�B{�'�=�%��"^T�2Q���-i����1����l�Ԇط�aҢ��ss/6K�H�IT6TK��h���F� �i<�0{J��W�~I�030_�O�)*ź��'=�i�`��!fX���
D'�ySt��D��BTV�?�ڂ������w8�E����pV�*;y�������w��/�͙��qhw�Ƿ� pe`B.����&�x|�L��������2H��+ֱ����)�V9A�\,|7�lΘA-,�s(YKSgʖc�>���18o��'32%��:|p����k4��+e
���_~�����{!ug����enLY֦���;:�/	���7����h����t�����  |F����*dx�����.+��Z{5��IrN_���������[�5���I�hۭ�{o�0�c*���|�	F����~-��#�:	�QU��h��`�@�;&데v(o�$��+��S��q����!�	�ǝ;w~������Zy+?\���1R"�M������{wt���,����(]���剨���% �U�b��r�RB��R�祲�4Ƒ���z�ťr
#��a�3�:a��o+���Q�wZm<�)H8n���u;�|�&�!,��c��,I��Zlͷ��"p̫K��f�c,��1KFH���:2�<?p�dϳiL��:ɝ�{>���7���
���3ݐ$�Gf��l���\������x����҆�a.�����'�1a�$H�ʕ������.��и���g�&� ���	̃4�҂����'����I����Q����CE``p��퓠�3�fM�P�'f GRTE�xؓ����$j���x����;��x ��H���2����L,)�VU�(AMT�7��y�dm�%��X;�Zҿ�!J��r
�l:K��fQ1n�!@:��Ť�B�sM.�C�����S]��0�~2��=�	R�*D�Vk�����@7��s|g�Z�ቱ��SKO�>hb�v��4�Y:_�ݔf�*�"�hH1��t�I�`C�C��QxjӪ��A]��'����j؋#y�Nm�R�w��:$����+J��b��Xb�zY'j�L;�:X��S��Oe(��-�����j��W}���hm����c�k�a�G!���lc�0j06acĨ��!�B�&i�+U�g	_�K��܆p,�*�B�
�����@�����b�[%f�z�-�7<x�@��m�6����cb}�}c?͌�?�716&������`r�̮� ����{��ԡ�ۉֆ4�����ٙm3�&��|�ϗ/�K ��=�ĕ&v&b%>Dd~��k�=��vkW���E��Z��L���ŋ�E�W`u�Бj4�'����P��o�s_�ׅ�z޾@@�����x$�*L�۷o�ɽ{w�������U�� ��JO*�O�-����N|��M�F���:\�uU�/͌J@$/�Lv,T�
p�
k-e�<
�r��b�]Y/H�G�?S����P�	fF.�����O�s|S$�z�1q�+v�??���o<x�����쒭��,����zj���R�/��L�Q��iH���V���k3��V�-��LH�25��t.�F���|#T��s�W��%��*���(�߼y�e�jKC��4��075�C�0�I2��ɣّ]ڄ�u�rA�2���8ἱ��ي�i��k#�b�ȥ`�&��斵K6%�-{iY"�\)�!U��m;{)�Y�!�������p]8�J�-m:�)`#K�/>}���ӳ|��Xu�<,il�z��8��X��h��)5j�@�2XA�&�l�Z.�'����ݽ{������V��U���g Kh�����h�M��RL!����d�U�C�ϡ�Xs��^���f�M
{	ǟ���xVb���z�����[��n��`G��OO�������Vk���/�%ӳ�G�l]��h��s��0����bJ{��<���)��#��2L���w��	�1vֶ1f���)+�ӌ �''��;���b���Y��4QK�˳���tξ�Kv�s��c���y`1�\�\X���Q��n��%�"�h�{�$�QǓ|.kD�L,�-���*f�$ ��6|��c��%K��t'���Kq�� P�O=�*|���=��\�f��o��Unauvy�X��Զ�gW	��z.�?)3���T�ۘB&bv�z[,"��� �A=H�Z��g���,jͪE��v�,O~���+�����u���ʣv�:�Ʒ"�>��q�2V�<��`xy~�#�T����Z�����}��@y��"	�\5��G�Q���&�F�������w3��P��N!�5�4������������
���ňm��@	�ͮk0P���b1Ţf㹒����N��i�र5�h���f�E$@��V�6Z;<k��?�/��Ҧ�4_Ht���].�bH^������C�U�λ�֬��C��;GDF���Q��$#q/�	c�I7�01U���xAw���1��j�/;Eza���0
�ApȦ[şK�#�y�/�TMH,�!�'Atn�<xS�]K��.kJe6��.Fd]#s�wQ��q�+��l�b6���BTQ|yja�<��Z%qd���qa-Skx �~j��ӹ��Uq���! �IVg�����a��jX{�m�I��"�5�Svf���[!��i�@���c`lh�G{Saq#�%�H
�1�Np"��.�X��H�Ԫ�d?eCPp�x$kJ+yH,1iOͣ�uɛ��`DOj]Ԇc����ܑ�/^�P�ScM��fW!�w���������l
%�jPlz���
&�/8O���O?��%��Tه��}9�|�ږ���`�^��2~W�l��v�6���L^Ӌ���n���\�͘���A�t�a��uV[�Bk'�i��U�3��yu*CakK�Si�R#���9(��-�K!n�Eжї!ߙ�/�ϴ��`J���S}K�⫂�1�2밳C��d�j��S�a�nL�R�l�Ev�rjuY�}���Ԛ29��}���}��� %�d)�HC��'������x�Fm��u���$������3�����x�g���R���X-��/Ѐ�G�u�,��g��K�=Z�#�#��t�(�3�V1:,��0���yH2���� ɓ1�����'���ܸy���$�%U͠��g���3�:���ǵ.]�z��ⴒ�2�n���fk[%H��d�Ɇ��;�Ġ�μ�un�an�C�>ho�K�5�|�9���p:�X��[֬M�V����2Ӥ������3�d�Q$�"%������zz2��	O��Ӟ�j����/��]'�aK� �G�	VZ��V�,�,����������(ɀ���ĸW�PiƀMj[�}a��d(j�Љm<��M���pD��E��� �l�TT�C�O)~����~�l��pɊ�H
s�8���)��ub�3���U��\Q���(j�B�\�G�E"
�����)���A�^���8(C���H8�2�I���A���*�N#3B�&i�5���@����ǌvP����{����_���j�@�^������w�'�����0o��I�ûw�	�}�M�'�(�:����t�����F ��Ƹ{�����>a���K~ik�����f�P=���5�e�"c�(99u�x�D<B�4X�x�S"���,V�#�IӾPE�l	\=�l3���n�Va���N�*N,����ԉ�9vI�RyŦ���ޛ���ʛ��֒W5�;i�aD�\	N�d2�P[<9"�+�(8��s����i4;�8���f�.��&\��#(y1�U�E�e��uS��×kT�V�rp߃�
k�q<_<����?y��٨/b���>(���O����;���6��g�9X��H��I3O����v���k"�$g���p͌<e�������K��Z��޲��g��W"5�	WZ�
x)��nNUs�-!�V
�6�����;w��1n��=(�{����L�w�@P��$Y����T�M�=�/���p���Foԭ����ə2:x�o�������~��)]�n��ݻw�~ �9�<� �c��D(�_��yMM��J��9� �⊹B(J"��Ɔ�b]�̰[��D�B�3
C"�
2�S�����|�+�o`�`T".elz��_�=��@�l��Qc3j`��W�:DH�J ����0��!����X
r��%�E��KI�#кh�B�WRb36���u �^�x����?~���a���(nTI��i%*r���˩ǀ�e�L0��a�<�%���Vթ��0i�a�6a[�cw��q�5iZAE��kU)#]/D^6`N~���a��[���T�u/��z��ƣ��d�*�YIgx�(���CEΓ_ɏr1��y.���j#ka(�f��Z1+9${S����vGڈe192ˎ�|�}+ a|�RP��S@BP��p�����a�<�*��@H��_�t�֛?#2>Y.��	�3X0�q�6{ZC�bxs{^9a��6}n� �}}�m榦i�:#�1���{�)qs��LVTܘ����T�m����^�����CȖ^���_<{�J�F�~��9��C)X:h y�<�b��pH��r��r��"PTA���e�ߍ��l.h�8Ҭ0�t,���ۜ���@ա�/���0"ۻ���*ö��'�]C�޾}���ʍ�{J�
�8W�q�w���m@g@s(& �i��uvr��gأ�r��&C�[K���g��F����,zM�?���p�&d=����|�I%���n����$��X��D섊c�9?��N���d�2���t�4�U�(Xq��]l��?��-���HU�������7���{E��B��&Λ�7��pv�ޞ�X!��R�,��C�r	 ��*w��K��@LH�H-�l�J����x�Q`
W'.m�K�G�8x꬟Q��m�4�g'��ȇ���O���_���@�6Q�@XX�u(�El~w1�/�ꯞ13J�~,�K*1���}~*����EbX2H�U��ҝ��
f� �J�]i-0$�r�=Ve�����s���w���*(ʼ�琮���e����ݱ��Pp���6�T���N�Z^.=;��S��#G�^��RҘ�u0th�/3o���x��h´N�3�5�J�WJ5����sl�T�^6��GGG����t1�п\��0���{�����d�=�ׯ_K��;�*��{���Fdb���%6��p.�Q๩/hh��b7��o6���Ʉ�2�2֚�,��� �p���<��3�I�a_f��x4��T/Kӊ��J�NA&#�����h<����|�����0�\.v:�7�_�)>�÷�6Ӭe$Av�؊!]�n��~�t�]�
)��}UR�2�u]�X<��_�l�`~��p˦�#�e:���`$����;��*���q:\�G����������������0u�x���^�2eYg�C||��Wx�d������Q��w���Л0�Xvۛӎ�8Č��U��4�Ƽ��u+�g��j_JoH"��8K[�EL��7��V�zѲB%H�)�ZY\�{��������зoIN�C�Zf��m�}ӽ{��_�����	�S�[Qo��D�����½�#�+!}OU܎�VMr,KF��X�(��i�V���{XtQ�k�܄'�HGd7��{�+Uzػ�KErd�;�	p�9��-�T�����2�~���WFG��n���H8J�Tk,E��s�}����#I\�u�����J�{mr$\�1� E�3}�}��o��FA<5�k.U���4o���k�n���'�iKÕ
�*��ԘxZuͭ��gg�ک�nt:�/�m7
j�a�݋�b�<�&[Oq#"�rI�[d�t`������g/n�nW�2V�[&�Whrs�a|��"�G�X|BD��^�z��$ͼ�x?5��r������+��[tt4&�1�T���cآf���{���j)g�4V�<���0+n]Ί��e�x��R�˺w5dB��D�KGL,�J���1��5L k���n#��X���^-v��y`��������ZA�S�/�B��1!p��?`h�"��2�be�gc?����kM�	L�\>�)�`N��}c��ؐi����E�pĆK�1����>bS0��V9�Z�Ȯ/�jśLF�p� ;�Lc�ȼ�x��b�]�4#IJ�l��vM����Lh�;�c�Tr�E�٭w4�B�� B�M�0�Ԫ��-����}����i�7pL8ʊ�]��7n���Ck9��S���l��{�/6��<�����Ub"���!�Ni1�30�T|���S�`��1ZPr�:�RI�š�2��q$)�0�O�����z�۔�Ĩ/7�{��e�H�1Քײ��h�Q![䭲�"O�*I����ao8P�E�
�S4�D�	c}6�X����b4S�bq�n����]W*Ub�R���\6H�K#���5�W5��~�����0��8�^�qLUj�̿���`��y8�˫����gs��aICÚ�]͝8sYz�+S���u���#担��ͨ ��	�3�����U!��V�'O�Z޼9RZK�.#��9�7[�qr���7F�(�l����K��@���+�ì|;5'֤Y��-��6���0�!p����',�/�:�>�k�zR3��ќ��[����`��ž�5���x>�A�e3�h
Ǌ����dy�p4 ͆�����7w�?����j��$��w0�F�e�g�YQj�Ve$g�f|��������1F�>��9����&l�f\�MU�������YE�i��ʏ�&=�?8?=[��a> �j�=5�3�e�ڠ57��|���8�Z���~cM-F�[`�0���R�$��h���H��D�v��z��^�9᷃PV	.���K���Û,�^��F�h,��~��l(�����D!`Ҥ
k�T��XYzp�&�C}1�a{��h��*6
c�0��]���	���j���®V���$xR�n�Bq�XK�����}�~��T$Q\xe����`>sݼ�cI��LZ;�أ�O����\\"Gf,����6����L��sE�[�	%��֦��Ç�X��@ �$F �\uIR��f��H�z��T�g`T�Dn�.
����:x|n�%�6��W�C0P�"���,����ķ�#�A��Ȕ+B�ŻR���Ml�hg��0�K�l)���z��4�XX�;rp1��
H����ũvoe�N*�Wq*�)�\qLm`~^�z�rbi fݭ�ROOD����l�&�
M�:Ҡ��t몣�qe��Hm������6Ro0dS�=x��|Mit\��bE����k�#��Z�
{Z1oN�!� 촘/ύ16L����D�����n&�^S� ��N�T�����p�"5ǐ���-Vr�t�����(��B�����wr�}���+j���˥�.�:�
h��w�����;�h�R�a,�������p�,�k;9��;f/��X�b��͋��;��o��V�V�;�����`2,�.��+	t-�U.Uء�O��*�������쪜�<k�̠b>P�Z�m3Ϻŭ�O�[���x��i�RJ�R,�&_	�۷o�x��i._P� k�^�+2C��׿��/y����~��˕i7Kgy8���=2��e�������{G� �&׬ak�+���di�4��	�Q��X�	�{�[�;;NZZD3'��t������L'T�p����_~�U�W���\��g�h�B�9�fx|!�J�zF���ߨh��f2��/��O�����/,�P1�M+���u��pTY�f�[�2�1���p�O�[)7<w���UZ��r��;�F0䧓�l���g������2I3ևG%cB���5�&��X��5��C�a�{��H�#ff4dV�ϰv��bo>L�"`إX(2�'�� ��D���H�+�D���+嚻cy�R��%{&q'icc� ���H�Nb>44��J	F�qܷT(�Ü�m�*���q)����zD8
0��o�� *w0R�̺���Ƨ��,S�^Ґ,��DCa6*a��8�-��c�X�%����]�4%6L�NU��#�6�8;+���C�zp���!g��0���\��-�J�v��e���\9J��/�̆>�	Kz/��ި��q �����!���w���[O� �ca�*�;u�x�K�z�f�Bz��4����a���?4��q<����fp�q,�l`F��=�-����Y�[,�L�����u���ƨV8��$�~ͅyL�ˤ��2DB7�+�b6�O�_��7(D�Ce!�;��^���4�wj�7Y�y���c󙭚�ap{ُL��V����a�`�n_agr�Z0u����ٸǲ�(�x8M�|61	=�l�8|�篙��]�F�Q��I���h2��V����yE�Ĩ��Jx`����I�թ�-��UzC�
�F�Y�YR�x���&�<:�:KE{)x�n_���
ԁ7j�ި3v���!���}�,UjR��S�E3�0�1������-�*�J�>����kC��B�lE�%�PX��@h�񫯾�2A˂�HKl/��kT�&�f�(�È-��{���ﾓÇ��`ð4,��C�C�`w�P����$�\���x4��UW�JH	����_èr��{B���n�:=�0��\!c��5��]eʻ�A��U$�����D5��b���[��&�F^S�
��)A��'���p½^e��`�b��o�e�d8��a.�u!�W	�|n����!�c���`���'o��g�jz;�X\]��ĬuM�@J;,kL 7��&f��%�r������e��?{��Q�0�_U��y��}����C��(���|�ο����|���Mx��?��c��7�|�bx�p͓���������NӺ@����W�;1Fʾ/��+k�qb_��^�mM��.L����g�S�eՠ(�fl�-	߇8��bb\3�6�������9�K���-eK�q�bb@(s#�J.�Ơ|W/�s�:ؽ��ҊL�,������R�j��EL��&��Ǟ̆�Œ+U�ݻ'9����۷D魈�E =Ii��ٍ����&��M�>��D��I̛V=�'����B!���l���_���R��֥����2ǆ��\�y�y"2
�斎+iˆ�]��B����w�6���$Ip}��NT���p:g�c���ǟ��:CӪ�.�GWWm'-+�"�ӲW.��X��R�XE��S���MZh�"i:�����d��L�V�d�'���4����9��n_�L@�@Llo��zM6���Q,_���t���)a�А��|���!�(�z��B���A4�������<n4�L��}��wN�����J!����U�4��2-A���O���W������P���!}	Y�9h���@ƍmKO�%�µ��,'
�jQ�������8S�K�
�S���1	�1]��h�g]</�)C��H��N����LF�v���e���RI��U.W<	3�S�s!�`��TcQ���)�:����ǩf��\��p��)f='�l6n�
�Ln6ܳ���?L5�$��x��+��͛�ќ`���\��0�nO�GF1b�Lb��d����G��j�}�9�Q��N��{X~�q]Rboy����������O��AV*�ɔUĭm��Y��e���Y; %��~F3#R5�����xbzT,[��! ��b�,��6j��p0������ܽ��6�w<|���h4��G���w�LQ l��.dI�n����'pk�-�:
��{��tW@U�DF,���F4_�B�_����d�0��"���f�#��'fϥ־)����i}��}��'�����gԧը�Z�9H�;�/���LQ)�Ė*�@H��F��
,&tyVcʯRP�!_Xk� ,	9�V��_|��F��z³sB���j������O���\4�]���q<!,ߏ-��Ȁc®Vn���Q��uF����͉�dw�
�5�/ϱ~�x�d���[�ݝ��+����AH1����V�I<7u��į`_�m�T���l�C�ջ
��h���x���#�.|�A7�Q�p�b�m�r�9
��#�]��u�9�1b����3Z�Z���q�+.�-��п쯒ո	��z��B��vDpm����g�}���-�2F��Dv�DX��fk�C)ǩI
m����TX8�J�岡����f�ޛU,!����G����5 �ECEA�)��KE$��*�c�G�H޼y�+��$�BR��xp�n��ܱ�,�vt�Ꚍon�lɭ�ө78T�q2�Q�H��Z-�h���@�8�
\D�4/�E*I����K{��?�\��aj�*��҄"ØՍ��w�	a��E���x�ǆj�J&,��Ǐ>|ȖY�β"�B BN�m��X�"%*vw�m<S��,���%"�[	�J3�-��F︩U�ܒ�ݒ@V�;���/��~����f�q����}P���q6�5�_I��T?�}@"��ϟc��Q8���ȁ��B��44cd=�(�y�KKb�d`	�frO��
�0��ɸ�U	r�r��K�۽䬛Z { w��mQ�JDo��,�L�t8x��'�Jd`�Z[�������Nk�=MaT�$Ä�V��.�^�0��ܼyS�ܭֶ���R�\̕�����P��ag�����"f��s�����t�K��t�'Z��z�ہ�`��r6̦��7867��`��~�������)fr�^~1_%������hP��t��df�|�d��w��P��d|��&��F�o{gg<�{��ݺ�l��ܳ�Q;4qF�Ƈ�;{7�'���]:�F�:��n�n�<|{��߅~��׌�Yl1X��|���߾9��
���Z�&^-�[�~�Ѭϣ1[�,��r�I�{ˈ�����L9�d��.�WZ�,����g�p4&Ԓa��2�Yh2���Y�~�N��8�su�&�Y��bݼy{�����bg$Hv��z~�,��1f0�l����t���=��U�^����l�t�f&�JV;��?x����ǃ���c!��_,�~7,7� bH�Ydf^	��dT�53�D��.[^�v=�������e�M�����֊mYGTN�y>k����~�lͪ�c�:3�N��ⷰ�vwn�Y�OO|FG�L�5�����|�l��^J�b��0��g�Zj�p2�U���w@��*)��N��o��Ψ�;7s���|Ի��\^v���{IJ\��\?��՛�l>�&�V�q���0B�����*r������~���hU���f�^?q�ýC�^�'�!6�[*�:ا��<�I_�y��W�˅b�}?L�����|b9jBf�y�7����2�Z(�FJV�vU�8���$��=~��i��L�����8Y}��0X�����V�ћ��b��|�IV^�/W+�A�	�Ĥ��z��{��~�0��E������4�D���J~�������0j�p2p��/ޔ�A�~��bD ��R�wan���չ��+�Gq�J5gVM�\��ًDT_�UZ̧��M���v��r��������
��-�Ҩ��^���rE�֌1G����h��v�T��̪`�0a�}���"�����b��h1��*�e��[7oݺ'��`�X#�����nl��ǎw�+~b�B��v��5R �ܻw��[�j�Sʕ2��0	��J-f�l�&K��?�ʬu_Ƭ�JP,B�w0�wZM�q/�?_9᧼ݠR�b�\c0*0Wq�Ω��8��e���G�>��<��o]]�'�#��8K������f��()Y�b��Ɉ�X�*u�{��}�rO���S�� [W&P��%H�2;R�w���"&�,�a�<�o|Gk�W�5|0���њ�J�?Ū9{>���ʼI�߻G��Td���N�.��ĺ�������L>�\C�����F\��� �&���_��-���y��tV�l��{�ln3/d���[�mwaU8�mWWې��yD/���P~��Wp�J��1r���w.��n,U���㡦Q���\�F��%�i4e���VS��M1������yƽ�}ҿ�`���9F���y��	�@��̙p��#�o�qxGfet�r�}뿢 �0��d<�Ր�XϨur0�Ѐ;����WS�}b�m�ҟUV>A�9o)ԕ]K��Pt�D�<�5�❾0'�1D@v��%�'*,��quzF�w�.3��h��K�(�� �>�&�P���pX���Z��DH��Ct��3V�7#����1I؉�%�J`8�s�k߬7/���(�W�<��$x��Ȥ��TO% �	8����f[,��t�l��3��bA��[��d�R�3� hև�y����>��]ڜ���V6�5�=?u=?.S���"�OM&S�/��
�ϧ���l�hmOg�`8�ɈY�&�&ӱ4W�`x=Fpa��W�����	n�0vj�`k��Sf��3I q�����Η����Q�8~��q������fMFÈt$S�x��Y�i7��2j�D�<f1�35�`��ƍl��x����H������<�J����֐�|�lg�w���,۾L��^�{�
q��T6T �SAܺp
�ELS�(K��D�����;�O�X�̩��0�ng���r��]�|#{m��~�֨�B%G��e|PsW��D@[�8T��r�s��֫dgg��o���xT-�� ��	�c<�&��w.�[���n��Y;;9���Q�`�p�9�\�R���|�Z�4ju5I͘�'ā��K!&� �iZp�n.��S��)[3���=F+`ˆ�Q�1E���k�p�0Tٱ|�T^�����	B��H}����2��(�T/=�x�-Ah�@^�C��]�5��4j�#A����_��Ҩ���lN��p��hԝ0�c��S9Q�N�mf<=��:��5��`T�$N�^�"��ϛ�]k���\; S|x)	�2���z�8d6_�Y�Z�q��w�u	�E瞷����*�ˎٻxuMeR�:Б+���,8�;U��a��z���y�v��k<�%�U���=��nK$6�uذ
��\�`���*פ4�r۳s�In��.���z#����|��yg��KsSK:)[�n�<����>Vu7��L@C~�7�o��c�1�q�[d�cKS���sv�Ú%��$�t�����Xi�c:��y����3]
��B���L��c�lh�K�}�IU�J�R�{#���5�F귬Ra�땚�,S%�v�T'�lǳ3R�)�W�^�$�����h��8�"�1��Ћ�e[u�THC[�W�.>)4@�e��|�c:Dݴ�]!�6��dV���>�Ί��^��� ��sK׋:�
�	7�OC6þ貧Ū��,E��D#�]�EC�+�;q5��x��F�$B-��-��3[�J��na=�|c����+~ ͮ|���.N��m1��w�Q)� ����ݵ��֜����L�in��!���h�.V]�8�\�r�����a~n�w ~����5W�!k����[a��B�E�����@��K]Q�nU�͝�>�s�ɭ9.�U��_�o~��;� �&:�Z��*��	���\�]����a��U������M�̖���� �O�R�@H?a�����^) �|6��E_w����`ku�����O?U�۷,�r9:�N��(i����+�J���'��Z���f3Y��,ՖF��N�X�O�T���p�>|�q�蘌��g�]�T"�j�T�q<���%|s���|�y����ǥJy2��"������ӫ�Ʀ��fg�Q���X�E��}�2�!�P�0���/�aR'^��a�S�9^�X� W$(YG�R��3�̄u�L��d�7H���Hr�g�L�+�S�;h�i�Z נTȝ[�(1��qϘ0��]ƸBv'De���Lf�n�a�\8��A��(�*E�?1)�5��R������|���f��p<j�u@NMS�\̏�}8*�@3Y.��ٙ���a��=O����ѱj���6C#��|�����,���!�q���0���>��ڽѸ�r�j�2��v����~y�2���m�fV`�n��P�׍����KE�Q�^)�Rf��KXV��oi-2��9��3`{�(��~��a�}!� <;�ײ�w,,dgL��$�|�Eo_\�!����i2�����߹�
Mu9%���{0ؾ���p�d-�=���OInb�zU\��J���`7[4�T���$�U��!aӎ52��cS�.Q��\1^%��m>�5S~�F�*��ܲ���.��a��b�*\�yl�xF�����c����>�s�h�5��u�.��x��|G�  �U �ȶpÆ $�^�J��جXscC��+x^�Vk��V�����U�QD8���qtr��j<�P�g���I���ʪ51���2B(����^���_W����U׬ �O�Y��U8�"l<���TeL����q�p8Ʈ�.:6�_|�'�D`qfD����=g�����Rżw�>Ȩ�� �bH=V����j`�u�]`��L�[h���W�)����ݻw�RS�3FBױ8oɀiD��p ��·�$��0����+��{Z��M5@m�=���ͭ��U\M9�e%2)D����`*����a�yy���������1;�֫U5k�- 8
����ou���Vk"�Q����%M��9��8v��A�Ra-	;7c��8;S	���>�f���@bE���f���N'
l���<��!��h0��#,�U���4^�Kxf��E��wa�>��29Z;���E㛪#���3[�u7Y��f��S*�m���|�]O���&B��GC�L��'a>���,9��������Ӏ`'�\\���6Uy9�r�EQ@/Y�2fq5+�g�b���WmMUe������AS�74v��X��Y���o���,v$�/<����sLU� �#�<H����Bۖ&���*�e��,����ҼҪ*�W�ɱ^�1g�hB<I@V$N*�0UA
Eʟ����$��}5�Q ���`N�/,Qeu
��c{SC���9�L��Cȥ�Ր�leV�bT�QY$:��s���?��?ŕ�c]'+?l#ޭ��X=
v���*�a��cjs/T�fm�8]�~W���@!e�(̬�������VI�����m��Gl����P^�P�,�>��/��f?��aD�R���U[j�$J���/y�ժ�ؠT4 �f�n1�^�xN��Z���%�(���\��/��Ƥa(Uk�E<�[u\M�7ҟ�����-��>]ݼ���_�z�﹫���37x|��n�g��L��x�zlW@\�p$z"X��Bq֋a&3C�Sk ��jB�a�2g0�¸�{#��W�b'���0�U���p��*fT�%��e�_�ҹ;�bH��`����sv�H�N}�#3�Q6�+,���ĺ~0�F'gg�Ng~��1�#O�����b�
�W|�����$�c�
8��GG�[t�.�K��8�g�*x�DY86*�2{t�E2���NWo8��HB����ŋ�t�T+��Ϛh/��mҟN<?�0�o�=����4^-H����e=�!�ᐭR�Z��b:sD�����P�an+W�[ޒy �D�,B�̣9�ݝ�{w�O��G�z��5�F��ڪOF� %fW��K�n�?]����Jg�IEv��������ޅ|��O�_(���op��7�����ju{�d6B�TkF.Tj��f��u�,��4��Q�BI�֐�2eT�0�G���&�u�X!˝k.n�g2d��T�}qRpa"�}/89>SO6���p����2L84�-+%��l`���5s��O���"��<S��D��3ZB�`0���vD+�8��&����B������~���;Q�_�y�)K��?'���d����63$Q����¦7k���r,�H�JW������1��.S�1���K�n]*C�OBa(D$X
S��9\M���B���*=��Y��ٖ�O��8���נ����_�+������9F�Ѳ���DU Fl@��܂2��I(�\!��f	�t���?`4ޢ�%h�{��'�6��栕g1h<5��7i���V&JV��\+�
Xo>�q�kZ�_�j(���+U��0����$s1K���U��3��¾Q��?�<Y���x�G����7�+���4Z��
��G$W��ݧӕ���(�@��-T�7�PV�P���"���ؕ�'����*91����%��	Y�D�����l\O|Z����L-�������Ff%5,�\A�*U��/m'ʻ``�u�g�5_���0�nT��(X��5�(���`�``PWϞ=S�h�m��,V�G�X���з�t���@A�h�~���t�1��Z�	�EPl��H*���fa;�h/��ࢺr�&HV?n!��TJ���I�ÑϑZiy!�S��&�H�+�zJ_`�N6/jf��N˂�K%ò�#���^��2�S�n�[�U�(�D�$N��TӚ��2�*����w$�u�!]�>4v�Se�`}�3�A4�I�B"}���T�`��E��N�O=m�V�����Q�3ɘ\g8jTd���w����$ t$6�'�~�4�lL#��{Ė���Y�[kT,P�\U���O��� ��y4�L�-�;+"�6��|c\v׉@��^'�e�1��Z`SC��:�"O�O�Vk�Z�O����a�X�{v>W���<y�p:f�"p��ⳳ�/��l<b�n�����y�=?��p��<p�Ã����J�4�GK�������l�TٽV�?R�����ש0�MZ.�&��X�?�������~>\��P͍zs�M��`İ�x:\����Ȫ�+V4�;9=_�hV�B�^�7ǣ^�Z��ݘ�%���O��Y�sL=|����i5I�,�)+Cl.�.Ix�M��.��׆��W�j����pS�XU�A���g�˖X�u��-��/.t�T�@UWgU��G�4j�ԘN�2�]nk����[�w�z	MU]H�j���c*��}�.�dpss�j����� O����bQ���z�K��G2��"�Έ����h���q��=�br�]�`�Bиq�0�F�PE�nBB�L�$2K񍻂I~�75����a���hB�[�S2a�7�+��8�j%.�J�\:=>��n�0�B�]Z�Վ��׭���9��.�����F]����	ø��27+���;\D��Ik��׻��+�WWݡ��ʚR. Fi��łZaiO Kϟ-�\Ν�-�_[N���҂�r�{&�L`�/��V0��8޺wl>G(�h?V�o�v�߻���� ���3g]r�Hac���M	��b�G�/7hx?�JE�K�E��*ƥޠ�4FXj��o����������˗q�j4�`�*�G�a	/�W��F�I���ݐ8����f�"�$f��R�=��f|u���x��_|�۪2�<�@�`�O�|2Yh.\.I��#lTT�b�#{B�I��\�|srr�����/NO�F*j�I�G�Λ��jy2���u�NIŌ��rC�r�è�*�� �R��ۛ��(���"~$K���W>y�'gC,=���3�z� ��&GDyј2+���T��w���E2��B�M�߻��Fl]���|��?�y����z�ӧO'(,����s�'do���xi���e��[>j>�E�XT|�H���ӂM��!��'�|"FM��.2Kk�d&[���%��D��ժoH�։SZs��V��h�F�ݼy�����\D3�C2Ŀ��R��ɼY��g�LM�d/>�\`\shئ�J/+'`��3 �SPo�$�ͅ�T��Ex%��)^�"�pA�pe<���+D3�,gW����Qt$��� V�;91��+�C#.a5~�\�A2J�X{��w�j̚@m��XK�����b�?�x.x�b�q,[��
}7Ӎ���2N�>)�*B�:p��A�p�
�6?	|���t�b�L�h�J�v��ZYE6�����K�u����L#�4���Qa���8��Ja��� ��}��,\���1�Uk�l*�`� �{��W�]R�P�	���o:8̭���a���t�c�"�|J�(�cJh�#�5��ڂ����\#����#�U�yU0����Ɋ�߅�����)U6��M�İC\�PDd佬V9#C���BE���R}ڨL�"e7-��Ȍ��i�.�Z�_�,<G�F�V������Ȑ�e	yGH*{�`]�v�_�|~��36f���t��vXY��7�8©6^�0���}{���c�����N���U����G�	� �ɕװ���bT����/���|'�Y�݃Ø|H�����~a��;-�b��4?�����>{A��9y�U&���K��NE�Xagck��� �x#`�p27� �E��T5���<qN@rAL���J~$����ɠ���^X���Z�j&�G�گY%�s?�,d��y6�5���x2��
���R�����㽝�*j��(H��Mb�<L�4�q�fb��x(���t���,��N���s�:y�\��j���o��!�����ˁ�tz'o����2Mbs�ƙ*�&+&l�|.�ƥ$��rY7������Q6����%��Q�z���������b?�T��^��.��7U�"u,D��Znq�O9Xʇ��Yn��M�)���`��#c����x���Z.B�H6rW������h-�CA���(�*��`؉�7Go	��-��m�nl��\���Z;p�
a>ʺ���Z̗�I�a������,��O��l�I���@n������v^�z�fN��������쒁��E6�zM#hD�tKh2�{=�6�È��'Jyjې}��t���\wփ�"��O��'�@�V�I�;�g��U�R���0�!��Z�l�9�^�Rf�{ۉ��f�F���N���=2�E��u������ƙ�T��Ȅ��ބ�\������_��S�b�<%͍�Y�,�}�3�3fpx��E�ɵ,�T��eFR~a��(1�b�#��Y�G�%A6`u �𝳫�����H�1':m���.;V��jt�H�"�����
;�HQ�� L���8���%~����R���ku�Ŧ��ޛ����.��8#y��^6φ���wr���n��zF�I6���i��Ծ�Y�e�o*����{\��X��;����?�#ht�2��J&�"�*NƦ������RLg:�,����Ik�_CٸV,+oC�����ǜ5vL����sV�8�S{���_�п��o�$;������W�|K��jI���~�+T�_Y�z�V�1�RY@>���d^Y���,����u8�F&�&�BQ*б���cʯ�~#)W
�K��
�P�%��(��U,�`�[��e���!�u�:��5���~��	���^�%<�w����O0�T�II�C���'� �_�b&L|���E�������v��g-�p2�5�R*1�.ckAy��n@��s*��p�xh�r]-���yl�$U-�������M�t�砳M}no����L��T�?kp��&Y75�)ڐ
/��Y�� g�FU�x�J�l�V�$�*s�[C�Vh1�fX%vJ�~�X�p_�6� .fZ_�
���������O�ڨ�+He@p�C<F��_�j@�RD����1�
=)�3���D�M�Z.�ʼ��1�k���G�,_���z���AOk��'�������Y���~��)��j8*��M�0��N-U���ks��/6}4^B)x � ����9l^t��̖�2���d��}�K����L������u������ �M|��|�b�b�XX�ѽn�MW�0�dB �Ɵ����W-"4S��7���|J��JU|6�8��䰁+���9�\��O�hu��+Qt`i<�:LZ1O`{��T�(0{���7�S���e<YXa���g����R�4W��F�K6���u��V����6�o_�����X%�
�Jh�~IH��`�ݦ�7����v+	噱o6����[��t<����ك�F�k6�-^<�$N�����3�g��dZ���V�G�k���g���98�q����o���J���Q��T	����Uʅ�]�� ��g�^wͼk�z�
~�#��x�'�b/"#�x�E�!@	��W%�粤9%�yކ�4����=�1�X>�����~�ņ8G��M�?<�����I�����G>^-�����3ьr��ŭ��[v�������I/I��A�:2NRQ�����쪎A14a.�'�?x����}z��vg��b��X���?��C�>|����ۻ;F����H��a)"��)�H�%��X����;[ȁ�QB�4]�̀w�*��"e�ʣ��%�EmQ�@�C��`Y������Ux���t�"����dv�8��<|�y��9nԨ�j�j��dokwk�¢��s�on��5Y�O�6�����?���߁������EO��X��"����<�(4�"��6NM����0/{��<�÷��
���$SI���"�*|'þ �Z�!dplF��w��R�Y�g�-
�-U��&h��������`͘H7+	/5�T�eȝ�\�0�TȎ3ͧ8�`a�q9�����785�?���� �ݡ��ۗ-�%������VuL8�2�g�X���`9�I��F�-1�5.�����Z,b_���ӈ��n:;f�94V�d~�n��w�}�֖��a�������d3LT�jLQfkT�����/�d��<�����G���w�全�<\lbY�[��e��l��LiXQ���+Vc�<{�,����$��q�C�W��s����:3�~�杭��z������p��	t��|�τ�pc���9���پ�T�=�Ea\lr�e��d�)4�`H�!��S�jYH���9��e��5�3̳�-��U��X�Ȧ<۰�[ϟ?�������!޼z��l��f�KG���~�;�䓜��RL-Vi�Ҋ�y�VV����Lu�;%:��hH#f�u������'���JM�r�*��M�=�ש6eC+ JǍ�� ~��HCK h-���kg�V�<2È2k<�૴K㷓��7� ����
[X2����J����"�����8i̻T�}��y�=���&�`e#-\X0� �����EM���ѷ?��9�8����r�XeO��c^�h�r�Z�*�L ��(f S4���Qdȱ<�P��Uw��uĂ9��b �@�j
G9�@!���+p��X8��l��7�F��<IW�;����+\�q<}�4�������O���f�����q�peVZM��*ZQ��+B̉�b�ʶfɚ�:?8��Wb�a��?��Ν�0��ǥr��cow?O��7�2G:cu�Z�$|���%���k�ܹ��<����0� ?Y�ِ����93��{d��p, ��E�i�C�'p�Z���=6�]ĳ�(Y���Z�+T����xzv�rt�"}�X%&#���~�_�����[,�ݻw�SĀ_�x��_��T}���>S�~�5]���!(��9�=pY�Vm�Dr��x<_, gͣ�֢}��_��
�	;[��T�UAh`�}:_��ًfX<QB�/�l(y���|)?��� W,X=]�����)Ӄ�g|1�0B#R�z.v}�º��06����O�y��8�d���۳m�1�H�RA��x�	�J�F�)�7���g(�!2h�R	�����˳s�q1��=&	�����N&�r�G��՚���G����W��9�|�~P6���8&CF������!���g�*����gL�����B�V8�Ϫ�QS��O&,H�������ܝb��Q4*��x�QU����ܖ��Х9"�F�o*�4x�lo�l�4����fP�lL�J�N��b�h��z`L�X�ׯ_[���8�xe1�Vk�&�lh� b���tZ>u��M�Hڂ�~*@��*Qm`������xXߚb)�0����^���_}��֋���Q�ܐ����8Ն-)�^���XQ6	|_i�V�!v��WlO"�+YBr>~��1�R&�Ń�(�U���s��S� ������B!ȏ?��C�,�{��j�16̗��o���Vk��� ���;]Z"��HR�p� ���*�"���yg����.ײ��$CJb����9f��L���[<]l�0|��ͷk���*2��j��y���/���ǆ���R9-6E���e��("��禷o��~�l(���S[��gF�F�}XD��*/����'��S�ݻw#9?����������>�L֫@�9k���y�2���p��]�z���pC���d�(�FO������S��`X�־[#T�O�B������q��E=��g��{ Q����:�a�� ������pf/eP5lf5V�Pd����MgL�����CΪ���R/&M��"����}P4q�]�#���[q�}�駘+���>�3�\��5T�	'����"��p�He^*aױ�ǒ�x�֣�DUS�I�(Ϯ7x�����vRD�aHVQ���{d$%�bCd�k�;�R��UȨ��cK�����)������d��&b�TCu�r���D��$��Wuc��c�T��N,
,�U�T��Պ�j_���mQ�n�X͉rl֎��o�"�>�'z��_>y�T�����v���K����O�>0�k�X����y���YG.��V��l%}�|V�B���)_D�A�FH,�[�AL��WKo��TxO��VK!A���Q%�v�f��2t�30���īT�N����u؂����e4��`G�Š��Y
^s��࣏��G~�嗅=�b����y�B)��O}�ds�hvy~fR��Λ�[�[��ޠ��W�����-|&Oo��<�a�����CYC�������ώ=�-�Y8I@��;ؿ���l֓�`尳��G��݁����e[��X�$�8�G���b��U����V�,D#w+
��8��2�C��w��Gt�=�E�8Yu���C��7��]D�� �-����8��a�-��>���R),f�I�2��e�ǝ�	�Ѽ�ݺ��M;����[k֬B����ƺ�՗�"?�x:����^��d�دV���y��ɓG��cr�f���t<;z{rtL�m\��#t��*����֖��V��̸A���\6F�:�Ī��l���'gm���^z=V6е-d�=L�3%�^����u��7t_<}Zb>c����*��b�����@�g��[}�;0� �X�}|�����޿��3������'�#�H�I����Rs8V}H|׃��Tj{�{o߾=<<�/OdvC�,�i�u��p:Hɨ5����Θق�\sg4�M�S���6�,D���~;q��Н/�	|��_k4݌/�r�Q�gY]�8�q�߃ׁ�0_�2�%v#���.���C4葷i4,�a-v;]QϮ���l����[P�6���{Ϧ�d� ^2�1'�����譈 ��ȉ�L�tV�̓�'��C�,�-����u�R�T��Ԟg�P�����F3�O�2�jَ1���`�}�#���8,�t6_^^����2�o�}��^L�e�P_&Kl�Rѿ���oC��7�L��/�����4ƛ�\w�������mxk	c��4�H���z���=���xrx��ȉUt��Y���E�,���u`a=����Ns���>[)Wk$<�?h�y��}��ф^E9��7�,QNXšU+����1aM��M���t�hz����ٌ�c��ޔ9�Z;L!��9vI�~��ٍY�~��E�y��]H(��5M�=�<��!@`w�T���7V�0�T8V��G���s�w���?4Z�t�:t<9P�w�)���қ�͗m���*Zu�J�����8]���8x�jcW��u�Aj@�Q��K���ή��13����v�
�x��mir|R4�����0+�w�>P7�v�l�u��x�������e�1�S�ی��p�C�Z�2.�����t�!~��D����u	)�����~�~��U�a3��� � �����}�nu�m�Ѳ���?a�ø����F�ͪW��O@f�JE���iSR���j���� ����[��r��XMV���4��p;Z���#�iC.��8�/���$V�VVU�䠕20h���j(cE�9�yZ͘<|)�Ê��y�����M�к�b�'a]ԑ[��e�)謤��:�ѿYK�8���{r�h�[$j�d��:�c��_�p/ћ�.x���<��z��u͖���P��5׬7�"N����M���Yi�b1�� NH�ᰯL��@X3�)����_~�Wx������;�gՔ{re�k �~��e�EE�}��Gـ�[�ȉ��G�vUٿ�d�l�"60>��Z�7u.�˿�K�U<�t<���*?}wd�	�ܚ�x�lA2���ٟ�}��'x^߶�h�ҺB>���C�0nK�!7+��.cqQU���bJ=�EA�C�hX,A	y����)�/m�p
�PYԎ�u�CN�d6�q����K�7�b9Ǝyut,��p�*rW�ƾu"L�(�Et	!��Z�ᯉCN�};�{pq��|���ˏ��g�4�Z������ӓ��{!�g��޻*�c{/�	3�ӈY�l�����?<�.�qW�j�����-��Iy�r��9�{��$�f[���@�������ѱ*%���Qe�znx���W$����<���C�XX���x~F�:|��{����S{wo�\����������ά����zk��C�
+�#6&2}p��l>?k�R�fk�$'��A��Ak���'�A�wkg2/W���xM�[l'o��-#�4v}�����7��=xp�՛#K���]y{�j�$�zR��o�E9�j�^A�tm=�}���ۭ�8f�j/�,Uӄ�_�bGXc6�ZB5Gp�q(��l�:^��㷣��r�V�ѣGx�v��L1(HU<K�?�-E֗�JJ�o��op�����3:�X�ֆv	����\P)�تs���pvB�ő+^��U�,�K8�o�O	��d��*�/��Zjlh�<��������L&�O�<4D�ħ���cmu�P�5�27��"}�K�|c��+���$QD�W�F�4��� ���5��Ƣ\�*��7���΅�^���\�^2�<�p4H�b�Go�
G�N��DP�Ea��3������;�����7��[���c7��!���捃G�nݾq���i$/�9j?��X�F=����1i���8wV԰���ۣ$IsYB��U�:�|���s|r��[�R-�X�$�g:
�a:���*��d>���}���c��I�SZ��Xئo޼Z��;`��?YW?��`~�Z
gdYHmt��ެI����p���%���DU���M�5m��L#�����U�g�e6Oz�ʹ�2�i�%6�h�^��2�r_#3�͗9�;��" ��u� �����{��-�;��!fwxRX,�pl �kw����Uz#'��2BM��PD*��B��
5j�YG�i�g)rp���Q�0��-X]\�U�u)�8�p)Z��W���'OZ��{�����ϙbJ������:�)�Cqg}���}�H�x|�>j��,���y3C��yr$Opkk�P�j����5���ʁB�n�#�!����p,b8O�|\?��jT0��cpw�~Gt���;���ңI�踪������ő��t�85,8�aa���`�cn�Ƒm�4������/vpIp_�|�B���=0Oq��
��CO5���,:CU��ҌU��Q���%}��p��q���i�1�A���G�yX*3���(�Ɓ��!
a��%ܚ��1���5�d���\���z�侘J��?�]fD(��r�c4&vb*������!���\��ym�������I��w�}����н"���Y��r%��W�TUn�J����ǁ�"���Ԫ��H�RH���#y|z"n1Ŭ�O���0�^�+�g�޽�k�裏ԯ.��5�(���hZ1�S5,Y�~ \���r���j�� ֯*(8ZɔBr���_��/ QxH�t�%������Y�7�j�"�T����!�Ν[�X�(&�V��"�ر�Qʤ��u��T����8�g�<�W��f]�,Fa�&�/¤��Q��
�����E��郟�6=���n�`�����M!�����u2���r<
�k`'���᯸�尭�_��5�������8f�:<���w4��.���w�#��gE�UF|��_=x� ���)7~z��v�IvZ�^4���)���:�>L�^w���iEG�w4��1��[�2����?>x��:���ّۥ�7nZ��8[,����ȵ�M2G�q?u��Q�)������3J#`I�	m����[5�����	K�n�u|r7��LY��a��`&Iq���d��}����+�J6�����q�o�y��zcqi��
[�x�f�鶱W�j��=/�V��a]#rE��D����+�j|�V��&����p_^^����d�f���_*U����O�)!���h�A���Ф`��k[F����Z}!�TR��OQ�#��$�L^>MsS.  ��>�N5%�ϤNOV�S���/��hN�� YeVox��A���6�trv�����NO���$m=fh�T���7�!�ECT>�vv_$�ha�������%53�nb���ժSp(Ib��TQ��I����%�lG��wɦ��0�ˆe9�Ϛ;�]\C�T��| �c%|4Hb&���6N�S�j#��n�ab%_F�$��i���+�D���K��	�V�W,���d�M�� μ�D]��1Md҈��6O���8����^�R��+r�K����p�I���J>[���C,����C�u��؈�Y?z������g3��;��秧�|�����_�������]ȓ��8��dگe��B>�M�5�s���t�]G��n���:�8�b�����'�|�v�aŧ^�׀�J4��BB�r=#�$�B���\6τf�#JWe�sD���C��bf�?С���[]��B���j�ϳ-�?������տ:o���4[$��9�_K���* Xl���V��ˋk���{'�O�q��!�h5BK6�W�Sˠ+���?SJI3{�F�7��d��xb���ذB{D�Pc��s�
b�����F�8�=9>óP����W�W���۷q]�	�g��̀㼰�pX���M�خ����+��Ic��f#��9�dF*�<8\
�k]��kF�L}O�%��1�S=;e3��/ ���"a4=��h��FW+�v�^Wρ*
Iu��śIDtV�ӱ���1��l�	����n���3�o�;x�����(D�`�CSq���8��4�c0p䃋�Wb:%��\���|�KR�M:4:�G�"�ɣ׻� �I�O#�{�56F����aZ\������c5�\ڋ�����K�B��̈�3vLq��:{DU�S�JY�����H�f��8&�NI��Om���2�N<�����r�X0$����eӰ�L�S�+�G�W_�gA(�Q$-�"|�(f�dan�Ν;q4%��������>�쩯-ژR����n���L��[-̇�7oZ���� H��dT&P;>i�.9��pO_G�&��(õ�?�ުKD^��"�g��B�[��%��!��N�p���r4.���L�]��}��n�MH_m�����Y�+f���b8\EUnK����FғFm.�շyK��C�Tľ�%�$d�/�p�{Ëf����^^ Mt�Xa?���W,_�]_|��a%.^�*��]���t����?����0��K[�����z�88��t��0_��wvr,`���7��[��RE��8�5���Y�ۄ�����O��b����������3�
<�������[bT/������y`��t��*uv���V]���X#U�D"��#�݀�ְ�??%��}������|>�F?�J������	6�k�S��bggkkf��.�@����w�~�1��3j�&��A���Í���+�?���ꫯS\X_X�:Ǆ�ۇ� ����a�c����nG\#;
��d���ŋ�J���x���5<za粅�e��-�R	����r�"_��^��xhy`�UɤOB6v��q�থؼ��=6�F��&��ۉ�5�gd����U�T�N�����Mf 75�����hԾjY�9via�߸��=CL?�I�+GL��{��	Ѩ��Ǉ� �1����ˈ�I%��z]�
�v��갋w��F{�yD���v=8��oހ=������L�m7���E����V��*�M�n�شX��UjI�#qY��b�|tH*��J�kU�aP��&QCq`�5�ñvw1c(�wa)_J���+���������H����U��������'}g膣��K+�����|:U��ƣq.��V*���k�H7�$����Q��O�����6o�O0�����Fc^�/��X]YM�0�s�'`�rVpa�MdS�)m9s�M�zc�+��;o!hE�[�T��������b� ��kׯkk�m��U��Q���mC!�G)Y<9=��E�,�+dJ�kލ��¡��$hJ��M�^ά�A�^qY*=/�����Åaȓ���w?��:&�g����^/�=�6,�<�G)8p�ث?�z��	&7bƭ{&G��r��A%(��#�S�P�>~��wW�����
$��l�oM��Ɠ^(��	�:��Iɿ�ݎ�7��U��t�௅3.R�Q����1����ܺ�|�f��|�p�E�siM�f�������p�bL�ƞ5{��T�U�W�@�Z�{x�r#�T>�O	~HoUM�*]���0k���*=�xْT�~T��->Fn>ׅ�U!��U�Ԯ�G.�JF�5Sh"Ҧ�� O�vt2���~]|^���G�[3t2.`�����`E���2h���8@��l-nݺ��\Bl8�g�}��HӍ�""0XUv;�L<��K�Y(D[\f�pzB�]/
M����*d9�T�@�>���u3=%�,��X�:�h+���RT'BF�"�S�:�Q#�<n�I�=�R(�V�Kn(��o5�eU�f��x�
8(�@�t_sIP�b.����]RC[��\�
w�d�����N�y.N͜k��US�����(��׃��^�`>ti���d]J#��TMt<$�N�:�����h���=�g�Dv�Qr�ǩ�X�^#���o�w���7a�H!��?7W�UM�*I�LH�^���[u~v�݉�V6�Mgd�S��Ή���Ѣ9�i��I�)���z��܇F�8E��V�{ B>f�_^2�#�I��)���_��A<���˥s{��9�<���?���P��k�\}s6l����j��A�A�����ُSI�G�J�
��sG�\6[��^��`�Φ��R��,���䜁�5���(��YÄ�0`���%{_[𒾴<s# wlK#�����3���TʵZ��K��1�=T��Q�͇�{rrt}c�'���/>�)���¦�bV[��Bĭ��7�g7o�#�~��'�畳�D0���.���ֹ^�DϨߡL�Z̦_��`�����0!^.5K�;۴�n
�5sy��6��|���L�^���Q��L���o�#��
���Ո��b�=.�0�(��Ж8��,��{�����M��r~[oy�c�ej��}�Y���<����3�܄�������C��L:utȬ�A^B���{�����Qg$Y_���m�� ���N�H��b0��d�zL;���W�W-O��0I�W�A>���vy�g	!&�(�maNT��Bh��onހo�������Z{<�n�qp|zV�֊��L�n��ݔU�6������&���,�3<����]kbw�+*\�v�t�㸴y�-7�?x��Kes�j�>O�y��D���ӥ�L�]˗o�����e����V0����V13ZW���H|燩9v�����0M������Y{��lG��*0��k$V��i���M&��t1�Hr<�p�Ҝ�G{̨?��Q+UG���93.A̕�b��!�T�0D%w)s��ߋ6���ݼh�(��%����]�I8ek�K�Z�Fqz�+(��Y^�,���t!�$`>zm}	�E�*�+�0�8�.�N��� ���*�zU�ymĸ�K�3�AP#�ݻw���=��m�91��(�&�hʰtx��\Q#�h����G��M1�?��_�s�L X�aw_2%x���^����$�"�:\��_S=ᠼ3�����q~��)� ���߯�X �.��u����V���G�bvb�r='�M2lx~�ES�l@1_�yq������.� ��d�"�(C���h1�H9Y&�cn'�dFv��Cؿ����O��@�����ž�_�Dxp�ao$u�;2^��?N���ϜL<\^^O�A�8�� 0�6�d"1�amG�T7t�XvSD*9�,�"wIؿ�	#�`N�;�����$'L�B����bu��ޘ�5��a���%�-��?�1�D$ uyV��"�_`5�$`.�0Z��Q�E-a��b��b��f��ݣ#��>/>]�"+�%Y�|��O*w��0�%��{��tXE$B%X �!�}��?�G�hp�'A��j�C�A�&A�����[��*����V!&��u2��n2�+ӫuJckȮ��Ԣ/�]A>��4�h ƭ�>��Si1�t�X���`µ7�)��oC\(\EYj���9�^������r���a�Q0�MEN9k�e9F��\ �v
�0�CD4'���xF1"�3&�I����"�s�t���ta~�H�D�X���9�{�S-�c���E������?[U�����	�(`n��J�Ӛ[�����z=�L��f�!W�������:n�x��>�d�|E���a��c�T���|��GF�0�.,ygι8o²�UT�Wi�ì��TH�Z.��QԃAĩo߾����X9(ui��:Ϸ�>{����X���)5�+��j�1g�A��W!��'OhD���:Vx�BU�t���v�wme�W����t�8?�`�ƭťeqB�^��c`y?x��(�gMoJ)|��p�(5*����L҃�c�I��Q�����u��Y8�ڄ��۷߀ݼh],,qۀ��|�4�_~� A;n���sc�h��<,�Q8�)����jk�����r��;���am[��a���ƌ-���l��hO���(�:�T�Q��<�V*�B>���q�LT���$/����	�
�7M2������"�0aJ�R�\���狪[ؖ�� ��85�`����0��į�so����F�gV0�ƈ:݉+88��O���I0��dz�?Py)�!���ecr`�^"q�鞞��b���|(d�=�7�〥ύ��w6�k�L+�a)���)?�ᒶ�WW�k|�Sm!�����p%�y,�ݽ=���g����Yr�x�d�a�̉���9�tPLH"����{�E�n�/,CHB(�n��d��&�|vme%r�.۽��r�^ ��l��ȱ3#"綡=C?[C�%I,���'n��W�C����
�kí���h��[���.�ȗ_~�E¢Ő��q��ܻ\���v�:�C�b߃+GھNި)�<��Q�@J�+<e�L�^���K|�ׯ_ǘ�Rq#��ṙ�Z�n 괭�-���rI�^,0�Z(���z������V �iU�	_�lS���'�r�EeNl40����BK��]��z� YC����s "��)�D��Ncc�S�~����?��TVMQ����sٴ��J��sj�,��98<!6N���� �,L*�T ����J��&;�䣦e�d3F#�Å��x6��&S��LjRA�X��F&@�_���=k�a���Mm�3&(kvc���'�T*=UUQs2ep�e��菧��J�Y�*,,A/T>�
�V�b"�-��Ly�7��J2���0�0n�Mr�ڂ����!\2��
�ɴRj�A%1�"k5Wٲ\*����S��]�2Nj�����ž%ܠ�*�(�B�e�S�^J�K}G����c|�*�y�Dg҄��. ��vf�.�"o��vPb��o+��s8,�!�����)$-%�u������^��d5�<#�t8A���J�cl��	n����9Z�^ʾbJ�~g��&�	|(�������f1ˊQ"��4�h�P;�V��5˙����rc�洎	���B�l�l����(&bԝѯk^��zD��c`��1T�EEF���$��0�6沙t����17�0�#�"�(��=�X�aIv��R1��xx|�~�F!�4^�hJ.�:w�22��v{�2p�^l�켘�V~�����.<x�n�RX��G`�t��L���`� ���9�m�a�w/�-�>�y����E`-���{0��l��0N�t��ãr��4��q��ݨak?=eMHmY�ɒ�y�������+�ȭ����%{V5��66�V�8��a�¬c��L �~	�9���///⯘��K�<'us�=���|cn�]<��+k~2���an�-�l�<LtYa��o!PH����T������U�5�?�a�� ����5�:<��*��H�,/W0D�N?A�w��R-S�å<�3�E!�q��Ѱ4?�����g�p�XfxS�s�l͌�+:n��G�V�RvMX[1�po浶��ӣ�&6 �+����C0�nq�s!�<��V�]2�f��T;��'�ۭe��%��y�Hҙj/✸*���s��ذS�t6_�v��E���� �p�Uۆ�fIlW�`���v�;�u1�ցc�"-*�]Ä�=�h��J�.�~ڌ�&D`��K6��m��X�*���f�Z9<9�qdhe�D?#��l�V$g�|0�i������qH�E7��L�\b�b��u�ޤ6W�W�u��0.-��JĪ$�J��u�*_������&~�׭v��Ͽ:;m�2��>|�����?�|��'��k��CF�i aоh��US�qF'\�����a0�[ZLz���)�#�L�k0��XJ�b7֮��D��� ���/�8����	���nī��W����;IX��HO.l"�$���H� �Cx��B?΁i��@�Ī�y�,$�D���K�8�����S�&d/!�>y�󅵕�Ua#��Zk��:^ă��R{���1¤7W���Ks�U0� R(p��{��"�*�0�(�ޣ��O�j@
3J���	�0d��?>+qˇR��r�LĮ:��bX5��KV�,4c*����W��1F����)	H���˦I�f��մ:Ύ��;;;u��UG1�g���k�f%^$��	��*U	�0pm�o^�ME������E~�"���F"+ f�ݝ}���R���ۀ�S��A�Kn	����(L{Dm� �D6���Q{`:�W�����y�h"l����T��[�D���A߸�J�*�*�!��W�YDK+g�%dKJ��:`5;Ξ�u���≄�$u
��QV��T)��V`����?�*�N$�� �6�4���z*kB�����j�<�a�V$��d��[o�a�1����>�]�w{����y���NU��[�c7�+݊3��J��d2����vѴj=���� 9#�W?�B�$���q(�eI!�&�Z����X��/��G}��T���_�WM���ob-���O,\c��^K��T����Z�����~�3����B�G���~�n�>#z��!9�Q�K ��?���s�Bz�"0�6���q����f�H��94�&\z�EC7F�x�����`��l6_no#t��?��������Һ7
�'z�6��[�/}0D4�`�1G����T����S��a��_�V)�0�beo������<�l�b�8��S}�4�E��D�+^~����X�݋N�<�����]�Kc�;�r1����������ɝ�ǣ��$��`4���9��Y���gϞX˕�k6�{����V�f��D�F�7�JW����@� ���Ӧ *�A��S
�+;_0����N�Y���o\S�JW�}�  �IDATc�aU�g��YiS���)�;0CU�lu&A�_?~�{pD��T�1��f��9DN�?l��!��O*�Z�T.#�aNfb�G�([�>��:���*LyTZ��ԮUȕ�}n����Ū��Y(f�,��3١G>r���`�����9���w�y����X�kGWo�tƭƃm��K�:݋�K��3�.Lfll�M����eM�L,�$�{��q�q��s�B�5���HbȈ�I�B�B���j��©��9��q� 
M�o8N ��c�d;�W,���m��p#M�h��=��,�&S)�`)�,��Xz��^��Y���مt�m�	d%bqh�v�L�}+�ْM�-���v��aK_Y[#Ƞ�2;F̔iB�����VĊC���(�a��e��d�ϧ���\�psc�|������5ޣ�j�f�Ot��Q쵪���R��	�����c�S���ض+����QM��WX&�%"�d��r,�G���dJ�qe����<��£��I�U�#���q�@�Z�h�*{gؓ^�D'�K�y���y�����̚��q�b����@,O�^��)���p��m
ѷ[�0abݻw���)�\�l%k�iV 	ǀ��\��Z�r�<�urLķ��@���
���`���B���cp��j��-p���9h'D(�Ig�0$buc߾w�~���#�Si�0����J�S�-W�\,�0i[�*Uh���.�I�� a�2����i�ȑq��H�|ᦔ���0�W�F��p�G������;h�8��>�GXYYÉ0/�t��#0��Ԣz�WW6Dj�[�#HV���V�����(4v��@P��
v�h.~����BuX����n��w1��-�)�
;����Td�Lo0�DkA�o%y		u�;�Bx��i��ny�nwt�z���ˮ$@�Du#̶p|
����M(].L�P�4�k����0%�� �d�io�&�+��cz��D�8C�x¡a�:mMBq$s��5q��p��\[���^��P���l�eV8�a؞w��]�+ۭ�&jHy�,Q.	+a����Z*�8��Uc���pGu�{Fv�a��.y(�C����0�����6&�W�8��(Ih�
#k�gTzs��~��+��\�@�u���Ve1_�e���S���v�}煉G��Zv?����-Ƈ���Sl$z����7���\��5����#�,U��<���a���Lp�u���\�5�&��"gW�� ʾ*z�f���O_W�G~"�ygGx?�����L8�߼y����_��n���|��t�;UKΆ��;AJ��o��x�r��?�O�q��ة�-Nb����T��3&d�����>� >����\qF�RL1�;���Rm4�g�Ϸo\�A
̭
��������c4 ތ��ul�:�-�iy-��W7&#.���.�?���"���ew��D?��[x�s0�{=֐3����ԑ9�������'FF�^(�66n��R��3�����N�;J�٭�;�^�?UV�P��F?�,'���Y�R+��V���Q����6Lĉ(�zTfU ������4O��R�t.���������O�n�HQ���T����Kwu-�L�(hv��ml��QZ3�'��$E#���a�_�d�֥���t�qx�)���߶���k��Qtٹ����a�R�4_{�^2�Sǳ0��X6~�?�C��|
����V�g ��:��Ɣ8=8�ħWe
�|�t��i�'e��GG����kp��ȧK�y����$3|*�&�7{rz<���9x�l���NX�f/5�,RYYYj4j�rqqq�ݾd�t�_kp��;�_8=:'���B4h�3�h�v;��7ߨ.��)�r�C'<�3�<;��t1WL{Y7��D:���`���ÂE0��#�r��T�+MR���![7�'�S�)���-���� W(Z�F�^�d�o��Gz�
���8*�s�`��b�+r�������qk�2L�e�J���L&N$B�����\
��P�p�sK�����ޅ�F�a�3�z�66���:v����+��!/f�{�]_�-.4���\5`0�77�`~%Nx��x�۫���?D��uM����FߐHƣ/��i^�o��Yk�}u�����S��+T���Tjay���8;y����Oz�`4�;�'�e�쏇���;!�A���e)WJ�v{m��t���%a�RܹY`�v[�V3�_��vcN<bYl�r�J�Tˋ٬f�+��8�۠?���d����9��!��}6B�q���dU�����?ē{��wa���+ ���0R'3������P�ŤF̲O����}�%¨�h�Ա�V
Eca��ﺯ>��w!>\��q�������T��J5��\��+uc�JKC���p3$-��i�E�|Lx���JwA�*�GME�N3�O��LABm[2
���tZj��#��}��� ���K�C�Ʊ��v�ked�Wk�c P�(G����=�E'nD�魋%	�ER�pڛ��>yL�#�c��)�"�gow�����~�@�n|�\���d/���+?�̪ 'W<T8���ik����6q�0�pf����h��� �զŪ� ��r��>Q	TE5
[g�"�7�0�^�g/�,�Y��Pj�!��=r~����Z*�d:��O&����X);��v�K
���7B�kx3B��84�����"�ĉ
I՚'�$�K)�N'g+���><b��Ri13�90v�fa���5�3�+q_|��ֶ��L{qX��_��$]���DgA1�%�m��ǁ{�q��Èaa��E|ri���䳮�#����9��h���z"�=��Hv�NF֖u�;��0�D��\4��yq̐����y��u<V��)�!}H�؂�S�������dLDumy����G����Zȉ��X���*<��[79���nFb6ku�|�q�}��q�ϛ$��5����IH~�I���ƾiDԘ�ē`�9���0����߼���Ӽ��yqt��}7�LӞJ�G��������}
<t*������)��o�..Ξ>}��{��0!��X�����\��9�zC���/.z���|'�BN��O�������Y��f�($����0��E�c���&�� 7�o�}�d��9v�h4����3�(ݓ��~���8�����5>!e�$]��jW(����%�	��eC'8�8�{FSq�Z�0����l����@�n�;�R��%M��Ã#n��Զ�w������������g�R��;���(E5����e�J�h(�6��5D�g���P.-,��1�F�J����z�Z)T�a%U7�3>::ff<��ɴ0!F ���X,��F
��CL��^�*�|6���M���Z��H�3�����@�34�'��G��D��	q�V��[�9 p�ʱ����h�vB���Z�Vc���V�.����}¦��xpj�Ɲ���7�ܸv�7�����%���.Gq���Ma-`�e)Fc���3�M=�l0�G!��X���C&���$�F�r�*���dĀ9~�ZbK]��r��#���Gx��f�g��,p�J����ɡ(���\�OX'���R�V��9j����[�6@��+�-�0��l����Ǉ��\�^^h�`��=e:��H뢍��V�O/E_0�v��yk	v}�(�05���:��7��)��p�2��{ۈ_s~*"Ӯi��	JY�]������p~i>���7�{;O�z�sqz��X��:���Sk�`�?��vhe��%ZH�=P:�^�Z������E�fwڔ�e�4�Cy�08pp�W��$Y���\m�L��E��9�m��7.>�B��/��j�����e�E}�T{;N,�:�Z��b�����&�C��l�;L��ᾪ�8~�#\����w��=?��K����>\YZ^Z\b�ữS`���bD�ZuW��\�K��|yh��,�W}V}Zm6�M�[��������\��/D���C�}���Kpuu�r��C�+��.�T�(+(��m��;�Ȩ�]=4z�����@�j��9NZ��ɿt����v��#�:-��A?995�'�Gss�_�j���S�0`�G�A��(����7.�9!����"w7o��	!9����J�bq�t��5�ʪ���/.��p���j���gg�����-<bp����x��^��
��,�s쥆��"T�-S_��d���6��l2�t3i�q.��Y����ZH�?��?�?<�J1�!
��s�krYv0��g���'�F,Q�ݤ�r�����8�Q�I�ǊU�4�>.�)f�Y"=W��,93
MkXI	���BE�L�q����;@��p��W�Ha��Z�}7a���)�є�C|��won^w�{ضK�Z�lЪ�O�4�76��oȳ�@AC���a�ٯO?������)���C�kT�r|�m�d_^^��OF���	�����W��M��C0w�l>����c�a5��8C�G�11�6V(\f�>�-y_�Φ<�����w������כ�`�b�+<u�6����;�`T�T��~T�7R�7����*a?�����6�xcuM�1D�dË�(��TA�����p��J����׋x�ۈd��~��G��������/0�=�Ǆ�f��hf&�[<x���a�[Y4�����$�f�2O�I�by<�~���Wn"ݨ�}/=���/.�⻷߼�������:=eձ��`<1t�}`Zvk����Q4Y__1�=I�\���w��N��$�;ϧ��MU���M	R����E���B�"�\�R���,|��\d�
V�h�K�	<&�ܭ���9���']Z^����|.�h�Q:��rũ�wdA����]�u1��q)�0���۷��}�ٳg��
-�Ȼ�WH��.�6���7�.&+T��8���XP��z�Ҩ�0��i�ǾՅo�₠g�"$4��eN� ��Ȏ�F�C�W��\̽n�T,�-��;�a�	_����[UF�RP��T�S(T�症�����O�d�X���>�m
|�|�M�"f��
N�	�t�=�Ztr�@���e��X\ZO&Mc��l��Ι���C�ϱD�i<k���_���sD�����ݎ�k3�L.�I�1`[���ҙj}no�x��6w�Ȅ��H��iW�9�8��Ξ����G���p��yv^.�1��w�y�U�Z��3����oݽ�i����Q����2v��&����j�:-	����+�6�w	'�o<u;�;}�['��֛`捇O�<J%����^�����l�VOg�gs��i�0�Ol)|ӌ�pan����B����tnmlb����~��s���y��M��R�p�:y?	�X�5C�Wh��WY��o���O����& �����G����X�7���U$�-L�\����h��~iw���Je@�485,��E\�O~��G���/�����_��9���%�yc36���C�}�J$��dB��S6*:�z/^Rm͚!�����h���FEե�L����Q���Z�W�4����¸���8ð�C�6܄�e��8r�>+����~�rnR��[Їб�)gF>tu�b�#�*2qܔ��q��b[OR��<�5�+5�<*�;;����0���8��x$'��Z�;�׌�o���G�#L���5%�TP�g\�W�v���r�8�J)�3��"k%����gg��%��W˰��i��9�0����u��R5yط��l��b��8�ݻw7nl����	C)*b6�9�:�%��#��qqQ��Ī�kظ~�������,|`e��&�#�'{S��`�s�[��q ���mŲ+�F5D����DX�E�)N�Je�p��2���IS���yq.t�0Q��8�)�F8�#�ؖ4�����U�+�8����Ʊ-���F��{�R#��P��s���WH��U���Lv&���X2�F\(iG�W��ÌY�%�+Nğ}���[o��6��a��DJ�l�I�7�U���~���=~���T���k�غP}T�(</u�(u� ��Q���Ė��\�vM}�2��}��ʶ�cJ�:�~�Pd�?fvtʫ����+���E�b�8޼sn �!1���#�b��0�fJ��ĉ�?|�z���
s�&X�"+Tc-[I�[D�������#&[��ݿ���޻W��OO�7o��ĝ�϶p�x�ʷ�����Β� �E�w�分nwz^m�/�)���죿-�熽�z)��P�_`�ؾ�Ȥ�p2�e��C$H(���Lꞙ,�#B�9������p�✑J0GN"�'�J�?/�a�Y ���������A��7��dHl���e�L�%�����}i�K�,b��.y4�%Vvan�s|��$|f8�a=E/_���A�0����
>CQ�t����ǣ���A��S:.��oo�<{�m�m�r�����(Y��x~�Bzͽ~���0���l�a:I�sP?������|>�붢(%LѰ�H���KP��X�&�T��G,��I\.�:w>c��e��~��o��|#\j��>�Ss<BxM�����kkk�tj�V��RC${�;0�_~���A� �T�p/g>���d�Ĉ4���UoԪ�y����B)�ݮOCnL�<��K��{�r���r��0���6iN(.�T�}�G��Z����S�|1��=~�9��a2�d8&.�\���>�',ml��kժ�lj�R&�$	#Z��t|׻� '����^.��i(����ʤmG\�����dB���k���ݔ���묬X+1��Z���F:q4��'M�7?�<6�0�j@�9m�w���Zjq���p��b�ק�/��%c��������lv���q�N0?���QH-�~��}���e����H{�ׯ9���%��N��d�<y�p4h��D� b�o���;{fT_��4��F��N2�N��Q\4�)p\x[�-���g{{�m8�$!X]]e�o�i��˖���>����xx�F��ժu�Pź7��������2�����[Ϩ:@ɰ}�Dwnߢ&B�� �ӗ2��x~a����NV�V��3�ޝ;w���)V��P~����s���'�@�|{<�~��adD���J�BTA�T�c����Q�B�}�ir�%��pL��y��B���K�Ŏy��-���1G�0���#�)i9t���6f�����p_r$���/~S�5�ἤ#��B�G�?�g���?��h���X]�&�-g��������5�����m�6U,,�cQ��]����W�]�F㰈�T����
�|g̨����a:����+j��p�h4� �1�ͺ7TH(���T.XSbUPG�PF�:�ByuɈ�qO�b�#�8�������O��~��X��Г���aٸ	��+g�ɵ��Ċ:l `�HK�Iue+Ž�(�(�
!٦jm%r~����z��t���g�����7�`�b(�K�P�+�x.Kf�҂É�������m�@JS�����J���#B�0��3��,f���H��b�E�?�Qm���=�f`e�T�hK�Z#'G��-��L�f�,ϓG��Ƴ3ٷ���\��sO!��c�[����?�P��jyb�o�Z�XPM�Xf^���^l�5��c%#�ܶ�Ӭ,��u�@�C��4y�Z���'SJ�.�W/K����y���T������xN�`�9	�ⲽ0߀{��b{qy����N�:cd�_�.��N��i_B�z���B�R:9C�NZ���B��*"����.�0 7��`��-ܻ=:�ч�V8�r�|��d���,�c�Z%�����Q8�dاE0����\&}�	��f�Mgf&jv��0�=��'Q2��\���|���iդ�C��nwD(B6/�яe�G��$˟ͦ�o�y�Z�8q/���Ƃ��+�j*I5l��u������&C�΄��Bs�ƍ�~�k��)|�."�L�j^�$
Î����׾g�u�ƱK�3�Y�ǰr)��"���b��ZC��)���A`�1<��qw'�<$��|&�a����t>�H`q8	�_{~|�:c#D�R_$K&�����t�8��FqX-W^�*�y�RZX$9������<�^��NϦ��!��C��kה��&/f��HZ�Tʣ�M�浛�L~����{�,��`�JBl�n�d��w{s�F�2����\xR�7&��J�N���Z��y�&~�y! � Vf'ǭ�ܕ"�Ȓ)�@���雷o�׊�/M/�I��U���(�t{-����|�`�9����ŕ
�g12�$��I�c���S��;�J��Ck�O��Q�Tc����"!���1I��������0\_Z������7�!w��%��h�o����
����`%DH������}�-<�O�����8/ѝ\&Uk�a��c�v���G�+�'{8�Թ	'�l:�G''G������0wt|�3"B�b�U�͂�V�{�?Li)H{`A��>��s,��1*c(m-�Cj�����ͱ���G�UjB�1�>�ݑ��R~7�| ����D�R{N�������|ssS�`�0Y�śAx�o�p|/R����X�+Ч(?�/ӘK�L^�M��<�AH`���]�gd>��N�̸4�:�Z!&�j�l�Y)�i���=<k,����I��]�9J0Q?��BF�*'^1�D���B��*s��S[[���cSJW"�Bͩ΋}��ajq����V��n^��؁YLD��,-�?���#��ι�R�2�Q�@2H��jc1�_��_`b��_�߂ƳʠM�vK�8q��Z$G79E�Z��:�l�bn<!�B�r����)D�!	��~�e������S5<L݄K�frU����u`�T
�U�a_�uu(� ���^Z��'�P4`]�l�裏<�)K"&Q��5�q1+8S��L�.����6B�b��ݩF=�jP�ǎѫ©�q4�&��U�i��6�ix0����ر	t��˷�~��Ln�D^��8�>Smn�l��������zyW"��<f�;�\.1
�_��תԪK����pW�)��5R��Ǐc̱v��,X#{���ꉛTF1�'�'�^�(��믿vl�c:1�3XJ�خ0�?��OH.�l*i�T��;�4-|}g�1�e��~?�˔�����L����[��0{[T���NO����\J�y��L����*f��}koY[[Q�6�O�1�q}�:n�Q1�;8�����/������Z���>���|)�8���Q�m��㵽�y����Ֆ�r���nV��m�MJ9�K�N�����`2���\��`�����ӧ[�T�9?윓�d�n�A�����k�&�������5ͳ�h��gK��B�a/v���M�a�Ġ�o�ƍV�y�|�-{��i�#�d������}/���E����Z�
���ˋd�F����Dt|t�g����þ����l.#���L��K0y��6r�d��ɍ��A�z8��q8�u��^���������L�]Y�[7�ԃ���!�tcuA	�`��������F]�Rgg'eӅ�����FcV`
���OO���Z��l^��mԖɲ޾��ݪ���~㎸=&�̄�.��Ѹ�#|�Y��~���{Q8�f؉�I���xd\��2#$*!�7O����g��J�^�5�(�9�I���;�ͣ����Fy2�a������Me�zc�Rio!�l����ꢍZy<�e��,U�<9�3ڋl��z��&=D�5N	��J�!�6=�ZuccId��M�燈|?ZZ�)�F�j�P��9�[o\�M���q#Z����Jeӥ�^r��5lXﰏxF7��ԪTK$ܗ��Π��c��-��Sb���7<G/�=��u'��9��v�sg���/������ٜ��>_�.o?�|2:��6�0�����|��:i^��*�|���Q�%߸y�yq~t��>_̉H�`⻭��N�c���ob��x�#&P��6��bdt>;�����{ￋi��4�z+i#����'v<i�xT��:�h˄Y��g�~�J�@�BQ=},�v��V�03p�r����X��7��� sF��16\�c�hc��'��J0y؟)`�&gy�o�Ŝ�K[FGv�Y���R�8a����s��M���j�et.��2斤n���>!
E!Pɖ����(fܩ#|y�c�:��ȴa�&��(��Px���i�0Ec�Ebʼ�VAׄ9'�NӬ�b����W���(G�������nuu&#_(}���6�x��oݺ�i]X~�b<dG����f.6x��-*���x|� �Ѩ^+���˃u�8�n޼�X���P������B��d`9���L6�4TB��7
0�������I��q.)�v�^��k��N���a���&β�����笆�<he��8r}QO�Y�MP���x���l��ɵRU�������#�kyy�!"�׆�`%q|/���,���J\j����1�ڬ����a,c����2�> C���_\P]�����@���T@�V*�T��"쑸p�O,-	-�%'a�G	F�DS��j�W�DB	:WԼ,ږ*^L�󩎪�����Gj+_V�m盾�=>=���W��{�=��߽|�R^2�Z�S"H��z���:T�V�&�=G�1�Ҡ��,+!��1O�$�TpR�e��w�y[���VՕ�'��-��:��7�m�u:�,���� ���~�B�}�j)Y�k���yS��̓��|*�EN�K��h"8_?�����d
϶%���V��/��섄hN�c�2;�c%����o���X$׮�$X�K�+��Ã���n�Rx!��`�*�\�)�p�4�y�Q�8�T�6��`�I��F^�O�"��j�B)�`�{y��76�C�8����%������j9=)`r�+8�8�h�m'�$�N1���`<wvqq���$Xa�h�_�{�25a��� ��0�����Z�Iױv�<�6o\�L��qm����_[_X^i��3�=[(��d�ɺ�����`��}fcZ�"��T�1Wn�/Z����Pƴk�Bz<��O7ڜ�����X����vݬu�$�g��D?��m��7������"[v)����2�d��~�dƟ_����u��D��J�꺷�pC�$�`~eO�R&��ff�޽{�1Mgc��e���8�d�^�R���
i�B/�O-�̧2i�Ε�Uє�r�xi�8i'���Re8A���Fhm�ڏqXG�=.������8Q�y��u�<���@��ˋs�r������E�Ѩ�3�b�0�tr9��7���\�b�vZ��B�T�������
~�F4�-�LO)�/ͯ�1�r�B[�A��B���9at��*�*�u���N;�98W*�_�{ݍչF�M��y��D��)�t�k�T2�&�|���ؔ���h]���a`��+D�c����u#�-R| �$�����_=|�y��ng���΃/�G���`i�� _(O�(�S�����+ ���
��i]��Q$�$����c-W��<�Ѳ��ӳGO��K���`�F �.�j7���N1�,͜���B�?m�n�\Ev�n�XLlY�!�����m��ڈN��Z�~
�O��j8�J� �j`���O���J)26����ׯ�c�9;Ņ���[��_?| �*G7���,�k�WDJ�xx��ml�Ʋ�����`����)+�XG'��BK;�H0&���G��({ή�ȑ�	�Áj$/������pD�s�X��	�4����:F���S)j(+j���)�z���	�g��*�^G8��3�������$[*VT$���"��g�\�r	rT�%��cL0 �BC��[�U�I�zU=\}�"�:��h����'����?�P�(8�hHXZ�'��@r��
q���c�uV�b������ť��#�zT�V�@���3Q���xCR�Z�J/i�(�b�*	v�xab`]����a���������0�Up�g�/KB�ܨ+ 5�ƅ�L	dP��B�`��	/g���n\���r���h�����욕PC��R$-���U���G����nNєh�
�(.f��zG�JĴ�\��L_'�����8?���iVWn ��w'�e�l0h�q��\^O?2�*�Oh�N���$�El-�6�.b�[���!~������G�E�lk��X��i�����Xh��%i���P}���C��4ۃO$��t&��I�P��uy�iϿ}v��c
G]f�0o>������^?��cEa:6���j�믿�t�������&�1�h���:x�ͻ�3\�T�w��_�77YP)�$���O?}���ݦ+���:^������֌7���P2|��[��8���\[_k�/D�g��=8.�:C�z)e��\����8�RV���h��X���6�s�Sf!��Z�K��2���9(O�]����ޥ(�H#��.)�LF"������L�)擥r�M\��fv�Q*��p�S����X�c^|�]\���/�Ǒ�u�9��L�؈47_	��C��X�_����
�<f�p��R�]\�j�s�������B/�d����<9��H��յ�Ȓ$�	K��	��2��jnm��~*O��ݣ��+k3X�K�@���Mz5�07'�%��'��NF�Ra>;'eYѺXgV*�(���0MN��;��
�G�[o���J���A�L�@���kK
��k�C�u&�\Y�K%=��)�%����K�TjQm�b���ǵ��ň�C��=�A��A9�Xvh��e���`�Af3�r%cb_�w]S�X'i!�g���jK��K��|������
���]2�%:�1 "Ĉ�,�3����i����w��v�dL�v�j}�?���^�0d���%��������������WK�����r>{{��{�J�y,�֨�#�o{$	�B�"�~�M{M�����=��I0ə�G+�D��g���dҕA����#@����~�De�c���R}�R��Q��'j�Wr����o����C?�L�,"I]�!�����)��R�����e�V�#vUuO���I�tW�!�9�	��,����0��T�@XE;l��M��>�
h����M����Ė4`�#1�G�s�6��a�&�����j�vs4����o{Ɓ�J*�L�j&a@*��?!�<��OO?�C_P.���Lh0������r��t��N���ʊ��D��9�����%J�� �i�ɦ-��q����W�����Xv�a�N�N�֏��*KA+w���[��3��L2c��əe��lp�%�>S�����2;�]�`�N��J���ᬘ���L|l�9v䕳��O*Y����R��s���x�e8J�ҍ��݈g�,��O��|'�a���h�ڻ����n<��d�f�#D(��<�uL��_�Y���*�_dn�.I�T�;bY
�xΜL!qhI�E�M�������+4��&Ǣ�ePȲh(8i&�0�����,�/�B����TU�na��X�;q��NK�9?�׬�15Š���/?���7o��޽���'�Xה5t�Q�����y��#&i�tI�EPC���jx��|�ʜq�2#Z�Ӗ3L��Q��&�$���Z��0�i-|LQ���X�J�u��6��w�1�r�Ԁ ���µ֩.��9h��KKsx�/��9GqJ+ē5%��K�R)��I�KÓ�e����Q�O���ť��-��\v��~�������P��{D꬙	�z�I�7Z\YFX�sx:� 7��׿�۹�A���)��ؼ�u�!��ޱf����������S��
9x"t�*������B4)��c����$��d�L^UY��e��'��Y�?�lǷ�0��:q�9��k�H�>m����g�7���$3]��2[ֱ��t�|����թ��gn����$~�֥��s���*��� Сd�d��ߨ�Gߝ�B��������E%t�s՝�`K���'��3��[��Z��٘8�d���u~�Rg�����.�ս��7ߺ�o����?��W�����+/��8��g����7@)���%�� :���9ځ�O|���(p(�AA�(��/Z�����2�����p/�?}����8�޽��H��V+�n��b�����}rt<��%L�^S?`�Z��Lh8����5�:#/pSɕk���gG�<V�����p/.c.�I�k�����\��퇑W,����ţߟQ��'���B2���������?n{��Dt���5����`4�P�eo�(���C����G��[��<�|��ڵk�uɍ��J��x�֛8����f3��G�Pz�9��b������������_�������w�9��WJ2����ROS���9L�����Y�M��C��[�r�ff�f�ѕ�"�W�H��;GH� �\ɫ�r���z�b��Q����)ܫ��ů~��:���g���=�B������옳��̶R� �q����p�{�ｯ�Z�����{~Q����Ւ���_��bccYy{{��Ç�b#Kl'"P ��N���1���E�����HTC���C�����;o�,�F/[��<�����m1R�5��	����߻w�׿����UX��0uj�r^�E�D��_4V@Bޚ6<�ű���M��ia�6H)��9���y���N�ޭ�occ�Hm={Nf�( ����6����4��3Dәlj�&��b7������CzI?��wx��������O�ݿ���?��"�z�!]�o��[��[�o���G��7�d�5��[p�[x�W��W�i�;�����g��ww�ٶ�_r�W��?��o�~�y���/��
21+:a����)Z>
��Թ��o����/��{�<���h��vͶ�͌!)/�R�0�I?E� �d�vU<�A������A_;����ӟ�7����> :m֛o�����O�]ם��s��ڻ����$%Q�,y<V���;F�P�?�����ɣ�h�pxL�F"e��"	Q"�@�Vݵ��Y�g�}���S](��F$ȼ�hde�w�}w9��Y7��x"ƑJ�p�����bߣ���Ew�rY��h`'8
��0B	$���>e��D�?S����D��@B���v�[�u�⣸��$�1��1����WÔ�QI�I�D���E�m���F�¥��wMOOcf�Hߟ_���af|1h�#��a�盓*��|��t�H�m�ad=zr5�~Rݵ>lT����p�{~:R���h��~�G%菂��}t��t��x�2�������$��ƫ{��8]�s�#~��{~}��>����ʇ�,	U��?��G7����Y��$p���5v�R���c$�i�ԡ(ɮq����;�D���l�T�c)e�e�
��H~��^y啟��'�ѨV�q6�E�$(�P�k׮�={�ҥK�o� ��@|�<��!	!�����R�Tj@e�)�{�|��s����h�M��q�����xǽs�"�\�EDzP��A��h��Z�a:ƣ!b:ȡR�qA6��)?!�}�ƍ[���,-_��n�߯�ϻ������\�}�tAT>l'w�d�>l�Nڠ(9�c�P����HK8�ev�|���-O���?���=�����:���O|������L:��=+)�a�'%��C�|>� ��=�C� M!#&����v�k��������g�阦E��S�����dCϗ��1��?��	r7j��(:�o�:]0�d2���\��@�ۇ\R��g|�k_��o\���h�x��Z.noo"e���5���g��mK�0$�G>�oC:�̌u��D��o�����.��q8?���e�V�г��e2[6�c�Z�3S��ps�V���8�d:E�7��J�H�L&j�2�\�,�qWlg�����[o��o�u����߽��o}�[�����3���'�&�R��c7�=���i�~�S�@��t�_�����zݣ��TM����j���;V���я� �����'J럞L?���{�),]#�#�=������|�; z��������-A�f�.j�D-s�B�Z�(��c�q�kDr��;l5��9l�u�gE��믿�H�}��˃⡓"i��ω��E6IJ�A*�s*=��Jz|mC
�t�~R�m�G�ȦS���j}*�IJ���\ّ
��]��r��������o��v��t�m�vq�e*Q�Y$�"�ƈ��ʮ�:(R<2E�G���f>_Ȕӎln�a����\������\���ɀ��+�ꙴG��\�����+?ͽ�'I�OG����#�r���a�O�=��z���0r�Y�5	~R(��u�����/b$
kVa}�W�I�0H��ko]�k����[�;�%������2�l1�JP�,;��c�5�J����e%�dS_!��������ؐEim�.� D�k׮��o��<�*��р��ufi��؅؝H�ؗ^z)_,�ܾ���6���c[��D3?�m���OP����݅�ũ���w�@`�S*�U��-,bR�*gff���WWW!˝={�w�D�D=;�Dq���tHe5���$
��� ����I�ٳ����S�1�E���^<�j����P�_�|���������G��_H_����t�/�I���ا���͇�N�)����R<ν�����)��Ss�'j�H�OGv���ώ��ƽ���X�?{��_��_Bx�3\@^��u������K$q��	8T-̍�5\]��ˣ0\�N%�<8��L/=�N�b���<�T����*_6���=��s�ۑ���ɞ�9v�=zu�Hu��D�es{�1=U��8�i�?��7��+������zA,V����\6��i�������8P�RM��p�'�w ϠDgYu=sl��g�apc���A�ӧJ��n:T* Z�ҵDT�Y*W�g/����?�������J	�"U��ڣw�G>����>?�"p��~��y�9�>���8GM+�~x��?����V��?�	����0����H���IJ �H�<tצ�wiu��_���h�����7҅�?{��v�ٜ������q�;�� 2V��P�7#�y���d��!�N,F���Ġa�L*E��_�O�qB�����	ᓆ����8�D,�3�|E�fk����7p1�{ESs�b�n�U�Q���s��D2	�ygu���/�:u��ۘ�������[�nQ%[�H�b�`mm����*�@4���Eug3���χR$����M.��!��\��2���.0�D�m��aK����Aw�����)��K�F "u˶�x"&MڤMڤ=�����0�T2��^��o��@�@!A�^�
2(#�ZP-D�'�|�����@UU��Ê��r�z�NJ�����УXVϧ�8$��& ��{��5r�����_�j`���TƐ>n�/"<1���{�H��񘾵��*R�\��P�_��Jx�g1�X<�>�1B�p,;�4�( o���Te����蠝0���±�~�����x1p�N1T��/��S�x��Ҡč������_���{��/�M��ޫ��	4�ߗ�_,�Ͼ��	��j�;i?��I	��M��%����������Z�ՙ���,!�u��c}B�1"�M��2�
�fәV��nS!z�:�(jv<g��l*-����"����V*��~�-�6�lԄ-�z�ѐ�Wm-
�lF�(9�=��@Me���xJ1���g�...Bu�hX����.��YT�ka�,۲������=I(�Y�$�G���f477g�A����si�HT
#�T�uL���\�u6�����_�r�R��B@��<F�ۿ��o�q����Go�į;i�6i��	MҨ3"������z�����!L��!wA	�6ۄ����Z������EQ��kQ�3&e(�8q;����^�����H,�7� �yQr{�r���W�򕙙.��~B;������ם��aЬ%a�S���J	:�9�@�f)J
sDV�>�n��7��0Y�Ze8�K,ϣ2с����L�c�D�@,��_0�?���P�Su0s�o�K-\�~�7��O�Z���ULw�R|��}���?�W����?>��rt�HJ�6i�6iϤ�dɐ"���V<��������^}���
I��~���܀,[{�<(��ٚ�x�Ģ���>�;6ێ�$�"���P�n��' �s��P&ȸR}mR8�F��%�� Ƹ�Ҏk
9M	����(U*X���������K��$�`Kj&���3"��i�WO&~��C�c�`;��CQUjiii��IS��2d\������%��]�1�?秠�b�v���7�=88`�+|�h��n\�I���(�荫pG��@�X��si��?�����/S��(B'�*Ȼ������'r���Ľ7i�6i϶	��bY��~���~���/_���E���_��l6���t/#,QlMa���Z�)v�R=c����x6�y�?R#�9���G�.��*'D�J�6�*?.2�������{��E�g8��B�<==I����4��Ol�Qu�V��s;�M�d��٩���s�~�v�Z�VÛ���^8����^'�K�j���`*���PG2T���"}�2����T�s���rV���&�����P��D*i�N�/vz�Ƶ��N�����7��0}�t�K_~�'?��������riq�W
�`�&mҞI{���=�����?���|���sge���kkm������mܾ��U�*%H^H�����)��z�q,�w�d2E%�i��q2�C-�4��]G|E;6���c�b<����nP鼹��3g�l�w�� �d�	��#�@R�p��}��z�!j��n߾].A�1tp��iollL�-�r9����\x\���9YT����AQ�v�^@��UQ��`��J�>�:EA������틪��Fh!�l�Qd��BāD�K/��jP�)�\��o|����?�я��r�V�&m�&mҞICH��ݷ����l�L��ԩS{{{��[__���\�[%���6�(�L�<�v:�|6�HK���)R���0��Ř�����n��S���t!I�.//�Õ��U�J��Ί"o}� ����k�JC���S�`b��j�,�<F�Z��nlb�.\�r�J�TV%ymks�f��K_�=����Q��5m��d�t:Ej��@����>�rgg�:5k���o5Z�,�q�Ō��D��>Q]�B�D��U�w�[{A��l54C+��ĭ�[�Wv
�UН2=|髯\}��o�?���W�u�Z�%9vI����S��{���?NڤM�Ͻ�%�3~�i�����y�G�T<2^�$}�;�����_Ah�g_��B*�~uThkc����3 k7�^,���VEi«��P�"�Pv2F%� �C)�C
���並��h��g�v��7b���m��͝?�����Pֈj��e���3���@u�|��l6��_�%�B�D�R���
gq>�>1��RH��p.�j�Μ9�я��r������@~�v��l���1e`��꿵�Ź��q����T�(����mS�V����}0 ��V,��R�Lr�P�|"q��9Le��cm�9c�4�̓���>�0�Q��͛7��o�����+U�
>�KǍI2ǤMڤ}B��>��$���H�����o���?��׾��Z�v���Q��QB� �䂤aQC�*i��(���bc;~ZZZ���ކ�II���N�rl�Qtd�n��:�����ebR�g�Ĺ�YP���ut�������llo��qH�'�=u����H��Z���x��055�ꫯ��)�MOO�k�������2Q�#�b��h�j�n��ܒ��-�2[���c��x��0���������gP��߭xL�a�xf�S��S�l2��SӌSg�c]J��a,-����������y!��4U�t�ubF�c�U��O��_��T���I��n�>�s��af��P���Ë$Qp3�"?F����я~��{|�7;��	��|<��w�vg�����A���N~�L��"����C��ƹ{d�W�|��9���z� ��2��4Eu%	�8F���v,gl���\6�j��۽nK��8Cmz�7$X�'h0TR>
?�+�ɍTT�Y r��H�à776�����{�^�>�)`͋�z�&�ǋ`"�o#�D�YL�L���T�#f2,0f�v��lT=��Ν_FW��SL(��@�t<�k�GC��5LV�`��������z�W^)������1i�6io⯪W�PQ�8��������"����h׺��N��Q�:u��^\\�"����ӣT�l&�܂A�@�p1��S��E��d
�q����5��N�q�bJ	DdܘM��+����.;��=:Y^^f���i�F��)��	�	��_��(eU�q�f�xC�e�qo޼iZ�o+�����ĝ�g�Nq�n�Vn�;����^&���;�mw��~��Jצ��R����p��e+�x&fX~�c�ܹ����G��k�c�Ǔ	�j�+���������s���.������w�&��x:���3�~��/�OQT0�)d�-�By�*�c�&���Y>q~�&�#��"�R`���;�bh�7\7Z�w��7��z�D�w���F>����޻FIyn���A�{�$>����S���x�u�f�.:�&�.V5���i���a�4T5��-;�J�26G�kk:Q)��l���H:�x��ƳcC���K��x 
<=S��2gΞ
C��B����p�k�F���Sd�ӓ��Ve*C��8�occcj:�Ao��B���
˫�벨��Q,�$�z�E�+L.~=h6����!��vvvV8<0I��0 /�V�Uv�l׿x�z�t��Pt/�"����n�[\|�F�n�C!�"��2Uy�m��_����)�sB�'m�&�v�֋b���]����k��.]�촾��/��d��t�5�8~	B3(�`0��Q���2�.a���ĊkߡS�K���q*~D�.S%=�U�@�@<A��
:���:�.�⩩��H<w����8�D�����]�l���ǳ�`z!��<�9�p*R���:��}'_$�z.��4�v��o���vT�5�+����/�������k������S�L��{\\\�5�N��)�'����g8��Cw�d�4&���Y:�s�@A����*ƫ�~yggg�`݃Z�/,.��������;��xbL��P�d��cח��PMڤ�µG��dEWx=����G=������x��^˔+KKK�djuu��-�n��Y�#�Z�@յ�"�x
Tr3e��PUeM3��B���E"(67
�j�����4A�2�L���paa4��j_�M��F����S�ljog+�/-�٭�-�t:E��X2��Q��gU��i|��"x ������{�P�._�I��w��D{hx��{,�yآL�x��O� S�� 7����a����/���>� ��T�*�*����	6�+�(��K,����nY__g7	�
�����W��Up����z��3��v�|�Mϝ]�&m�&m�D��*(x����߼s�D�|�
�~�냆\y�P��Z�"H;�\.�J2W�&��5�����Ѣh�@$�\W5����mC�.V���=<�׫PbI�$	K����ONz�È�lP�[�,.���P�\�dk�4�D�Z��R��0�S���lO����h`.v54��$Rɸ�M׫��S��y�����SՊ��~׵�k#N�Ms��r�T*�>M�� �`�Xp콽��o;z<n�
E��P,�����qQ:�;�0|��20�J��ʶ�UA/It���h/��9w�9�s�w�j�24�Q��ӷ�8�w�������C>
2��"��DO��
DOڤM�ϧ���<pC�ṑ�ˡB(vcY:<�������4�P��V]�Ѹ�{�m�\������aY�N�����n��TN�H���*�Ry��'�c�v@���a렁Ϛ�����	��Q�0�xli���,��ݾ}�����}0�B.%G�z�F��@l_|�R�V� ����Ѵ#Z}2���Վg	�XR�z�uw/�e�$���+����M0Ʊmݺuj�~K�OMIIF�<(\��H�P���7o�D�1#���mYY��@p`Lh,a�Ρ�ز��]�&tpxC�����m,�� `*i��;� c{���1���ͦӘӟ��g��^xA�tG�cV2�g��5�x-i�&mҾ�-�|��,���x�$�`%�s�����=#v��9� �oDs:�6dY�p��{�g( �P��L1��(���<����>���ܻ��JV�Õ0������3���xb�H���r⸞�W؊q4���<�����׿N���(ꃋ�}���i4	��eZ���j-��������@�2)�o�5����m!)�e�a�����^����/}x���h`k��tqg4�n�X����R�Yh`'�0a"��7����Pa�  �#&� 4�l:��<w����Q AX��Y<jԝ�������i\in}O��#{��>X��B�*��I�Un8��F�� �>
�2�H�<i$G�&�u�������Bf��L�#;�F���TFɱ!���Ɋ5"�s1����6�ah2(O$�C��.����fCK��a�Nk�2�ЩS��DD(g����p����H����a?��O�J�4{�l�����luq~1�XK�r2���P���_|������{"�nffb>���j��	��Kh`m@��Mp��\��v�&s�]�~}���9�����b�����ٴ-�`?Xh!� 0y(4�L_����x6o6�?���D �h%\[[����]�H����Ξ=˖(�D]'.c�&Bi�&mҾ�-�+��`��$9��R�� ���?����֛��xf~~qqqx8 i�G��/. ���U$D�a�[�*�S�3~m4PD@�@p+ϥ�U��o�ͱ ��C3y��5m��"Dt��5�] �S5�t������7&��z���ʜs}�Z��I'�E?��l�$��G�r��FK��f�ƍT�Jrgg*��0Y������.aӦ2 �����s�[q�w	�+���s�_��G��I7�0t���CJ:�)��T�(���{<���s,�_���Z6���+2��2�����]Sr������էk��{�7=7����<��)�r��֕+�"f��q�8<ϧE��F�� �I��M�/h{0����"��P��PTI�iN(ml���;?�����e��Ν�W�=�3�#=T]?t���A�ǎA3C2����݃��+�)�}P���Y�� �T�O�*Dkja�x.$b%�������h�9n�VFg�{۔�(�~��3A� �C������V)g��rY#����g[N�Z�ק�HV"*#(�	�"�''�SXG����U��3h+^�R�@�O�~
J ����G!�˪��]��5�d�2"����pE�+h�3���R�&x~6���z6GթzTQa����Th|l��E�`���8q� ��ի�\
*a�p�]X�H����6ͩj%�ΰ���̥I��I��7��>h�dyT�{g�?��~�7??���@%���|,�i��'t�H#����SX�q�{=��K�EÍL��=����)c�v���0
bHE�,H���s��I��}�BeR���\�|��ӵ�cbs��bP5@����9�p����)���p$18��)2	�����M�c�zew�=����7	����s�v��wށ��G���n�s�V�q]����;5MAo�\�A�1e�r}vv���J�{�;��E�8r,��E���D�`~�l��Ǔ�t6�N�4C�tzo��Sl��
w;h��2오�u���]5�x
�k:��@DX��t(Q��}S2�_Mڤ�´��/8W�(C��f8�-����W���w7D���y"��@T�nx�ݍSM=5nXR䄾�ǻn��mM#�s�Nl~��BT��7��O$R�BѵvW��eڎ���0b�nd13�PТ��TPH�"6:���i�7�.|��tUUj��~�R�:$R��I�����MN���!�ߏў���*�H��*�H\�x���Ô�J�v��y����p��J"� Ӂo$1A��p�ere����+� ��x&[�nnQ%�b��	�r��1f�9 �ٳ�B	���S���i� ;�.TsX���rm�_|�EH
x���.�t�k�_��*��|.�/�i�&mҾ����p��@����7�xcskt`~�������:\y� �4�6@"��a�I	p�1{¹�S�d2	���@�9n
?���O�o]��!�U�&]�N�袜8�=T��SN�K�r�
��h�������ӧ�T��-<��7$M#",���x��)�ƃGqLF�?�����T�~�jAw��Uݎee�]��m���;<�����B�P@�C�K�uj�ƌ$�՘���:Xk*�M�JS3�kkk�[`M���u\����v����ۊ�+�N�Y����>%R�+ECӱ�sKs�li{SS5p�N��k$H��n�֋/�p��yǱ��lKy���4���k�����/<W�V!�\3��*�"-H�0z�G���8*���y{�n�0�D���_�JO��?GG�pw+��:H2]-�d^��DT'#�2;x*$�f���������{�޹��R;{-����g�$���v�Ou�Sq*�Z+!������GQ����EUQ�v)X_��c��xTz/a�\�M$UCS��k��|�\M�O#�ȇk�)����m:������mޡj����[�=�ʂ"���E��g�y����ų��������b�>�i���y8�����<�������>!���,--mmmA�����[��'2!�8�&��=a:f�\c�B�w�V����jnllpaAǅ&�Ω҆�a��w	2���b�p1�$8�����GF�D@e���u\L�:M<,�\06s4>{����T&�1>��ȿF:�&.�I��ϳ�� �ѓ��,1/�q�P��݃�իWw�f^� 
777�!��������^(��dtJ���r�v/$�. �n���K�q��y�,�T)�2ߌG���)��4Zw���L�A��,,,��F��Tr{4��ѩ�*#_�
e�I�
���D¯|�+gΜ�TM���Te���Ϝm��6;;K�F#��g�_����ڵiI��b�K$c�1�83�t*��V�P��iH�\P���`�?����p�6�7_��8��x8�rb=��� �taP�P�ٵk�̱��9�O���{{��CN�Z����c�q�t"Y)�=׾z������Rȧ�Il)_�P"�d5�H���O�U�0������b�~Z�2�Î����6|!�� &�P$Ų]-n(���<���o�	�V��t钞H���޼��H$f+5�4[���I��b��ȿe�<""l�|6W)�ww6]ϊō��
�TOM&��|=8�I���fB	��g@�5e��C�������������C��ǌ�p@��ZY��~�m��T>]*@�.\���������\S�֍XB�\�g�6|ϫ��30) ���_��sr�z�J�ƭ�z�V��`�k\'��n�0*=l��g�!C�P��q�U bX"�f�=�>C�`�f㐊DI��ӧ �`��F�q��T%'�M�E��|[���ߞ���:u
�nW���I�-��{F0�6i���vl�P�#�溾ah������ n߾���?�zn����r:���Ơ +��ܺu��h1���yь8�j�,���C�<�Q��h�e��9�h���T���g��+%��q�ƍAo@֔$���#00�u�_b������ ��PQ�N@?S��/�?���ŋ��d�O2���~��e�9��D&G^d�C�_^>�ɤ���,-.��놺���X���L�ד�c?�^<�JXY�8L��`ooODB��c٦f3U#��_�夐~<}�,f��񼩙�I��po�`vf~�܅A�ml�x<9�����@����1-��Z[�ٙ������������V5���zg0������|6��C5H"��P����o���v��>:	d��Lگt����ȡ�Q-����BPYU��"�J54:��b9����ʝ;�����,�Z���|{w_�sr���'{2[�A|@
 _syP���򙴢�T�¶�
�,�Ԟ?��-r,�y2I5�М�S�p�\�3��(c\����٦H��TA������0r��8�R���`<3�@LK�50�Aw�kf�d���D2>�+ַ8|�ԩL6DT���D����� �����s�"W<�d,x5��1�A��x��M�Ƽ
��FL���]EC�Ds&c���O�V���SR��)�	�6�a��B���	�0p�����	e���BpN�k��6;;{��/_�l����^LWIϨT�ە+W�ܹszq�``��H7�
�� y}�&mҞ��ӛ����o
�(�������F>�P�x�w���b �[����hl���LU��dg<�D.|`�@"����K(���
�׿����)��J�
eb0$@nQ9#��T ;�ґN�@�:��ObY D�@O�#�2�_"�q�*��H���!�7�ѨU
�6�l��7�Z~A�1H�ϴ}�F*BD�r���>55��!�s3���k��r<�ʥӭ�a��o��F���;�R���c�.
,����]?<�AU�Օ��q��]J�H'S�A��"f��V+��xn80�H��[`��Q���i�c�>��Q<��sy*+;c���C��w?H�j��Lf\��o�7�w���J�
v��۫�[;��X��.��U!݅���y|e�f��>i_�����a�qE��ģ���h��ˠ�hI;6�BȠ�C̮NM���ng�ڈ%���F&��$Y��J�t2�<��u=��ǡ1h�nY�+[XX ݷFC�E"�)N�{{�sӋ��M��k$�L�B�$�?h�ds���ܠ�������zn�{[�v�V? ���ݡ�G�t6G���^��r)%*��*����O�W*�Z�
�(����q��g�^�7Rihw,�����,�ob ��,�K��U�y��{��/_�
��!��H]G౤�Ƈ%o���&9'O�����}������:�>\��or鎒h�*�Z�����s��\�WqӔz����_�d\��y��v,�kw ��Ncl�M�f�ÿ�+ ;�"u��1i���5��.��L��յ��W�B.(�k��@N #AXZ:Cu2��@��q���!�r&����P0Jy�T>88���Tbss3p*�P� �n�����ƒ�Q����*�T�����o߾�N�@a@
���>T�N���\&�Im�B{")Atg��r�֭[�}��s"H(AiH
t����a�3d�V6}�h�_�a����GT�����!�(��2x���� ��ۛ`�X'��q�X>_��&�L�K�/a	1�����������QZ͵����^�8]��~x���_�uv�c�`�ɎwN�F���v�����hau�#����������`��oul���cظfe}5q�g�*�2�M��!�Hr�B�j�v+��(2�,��o>���|�u�
ȳ*�5i�܍�	G�o�#=���灂���O^����nt���'�E��2#���u
�IH@��u�J�������ʇ�~_7��9��LP�ӧOC��c�t{����)�$zY�[-�u#�:����t�
B�KgF�A���Q�i�{8���$�J���{a�P����/^����R9�0P���3j,F��1#6�SY'P�С0�b�@e���L�P�/�L�J�x�����*F��t��5l�v�FL
�R1���Sg���E��g'�|��3�680���ruu��wvv2�,�n�I�b��% �J��-ǿv��+'U��s�3x,څ���2~�p\ �G�?�w�}|����4pu�XA'��.�ERg2��`��O�4���3�K���A���s-�R�H���{���4)��eee�W��kB#�#E�)*f��\l8���~���'����(��HN��OxƤ�Ә��'�U�f���aF���a��,�?���p;�uޓ+�'�������0`Q[B�������;@���ځ��w��+H�[��h�P�)�d���C���k/uUUЄt�P�p�AU���H�ӄ�J��c��H>��n��9ls�Q+�8נ	�B0aߦ��?������Tp�8��ǔ�75�nTP�-�C�kh(F1�ï��`��V�1w���3��Q9QUP$�N'��1ꙵ��%.L��x+f!��������:�i骶0;�Z�x0����tufv���.�	�$����K%ҁ�k�T*P����KE׶��J���A��,<����o��&6�����Ƕ�D���*��<�\�ݲ��@�P76�t]ePw�C���҇*j[*U��؈`9Y*�xJ�dc{�!*P�(�D5z��)I���R��U��J��$B��|"L7:�x����p,:o��e�|2�M"}'�D;IBF֥�����ƌt��?�q������������yG�A��K�siI�Pegg�!�����SE�.arh�)��rzk[`	8���tܖE����p|pФ�L
�����*�e:��d��3�KX��C�d(��2ǕrI	��u��t;��ftB�M86�P_��)�	[����^<EUZ�X2q:���1
�(0�%(�D"����d*�ɠO���9S[�&�A����Tz=뗾��3g΀tpL�ٳgc�$�7����"���g�6x��v��V���y������3��,�M��Ύ�+�(�Έ� ��N�xdO��[��76�%�����}xН;w�,0Y�z[㑅���V�}�ܹ��E�E!����G	�8F��699*"��G3hU���x4T
.�R��(*L#�^M#X�N�|-Y��³ �lo��b�T�X(@{=�yDw�Zق�������<i�v�o��!>Z���ߎa�O��w�cڢ���y�s��KA(j0ˊ�8A{{{���!�8��^� �#��<$T=�`������Q�nY����[�>q{eU�=�p�$`R)��2��o<������lr���fWhZ4\�����ur��#����Z�\�"�=�_E�� 2	"h��n�b.����k7	*I�A���@ͲY���H%�eff&�ߝ��Xo�<Cf>s����S*��,`S���\x�9�|jfH�
h��e2����
%�s(�E�f�hr� ��`T�5:��PA��]���pg�������f]�95X'���e�'lll�w��犖E{�$aK�)�;Flws�@�t(l�F�6��ΐR��Z�^��b�x<�9��'�#��t���uEN�Rϴ���T"�� ���'��)?"�'!b�d���*1�����I��ht`H'6����D%;sc<��G�NCA��m��1܏�*Q�L���� ���A��D�x�O�XH�IƢ\����I;#khۭv�'��z\"�qgg�C���2��!�l�N�́
���������D܈���6
J$�i*wà?�}Bڍ�񸾷��Jv��*9�S�w�\��V蹸�sM�Bwl������BF�����.���]5�%o<'�����P,�~)Tl4b����ܨ��m�M����1�����v�4���������抔laں0�փ	�A��	�V���1��N �@X' A?��'�� Mr��\,Q�+� ,����>�3C��	ݬ�������?�Q��R���ۡZ��a��:u*n踾����ٙ)Q䐌]1��(do����3"1��.5=��E�Eg�%����6�	���{���T�NB��z2���I�s�=p˅'�ޓ�� ����]��#ES�:/$�%�J�P�g
�=8��)����9<<��V�N�`�R^��.n����@^!��b�t��- ��Ҍ&�?qT�riT����m�Ӂh(,�@�S[�*�����+�=�ut#�tU�,q�29��庐@�zrDo344�*T[	'� ������P��6��@�D���T�	/"	|\*�T��E�M �1�Od�϶}�~�|�éHGێ��)_,��ӧ1e�.QC٤ZI�J�
� ���,�F�` H��T�T�2�����!x�L���N�|�l�ԯi�z�O܋�XXX�����A��H4(��J�"�^1v� ߗ�e�ێ9;;˘�plr�'*F�����AK��L&K&�;w�^���d%��4����'ܰ?>h�Z�a��;��uݳ5�<��DI$qa�+(�4O`���hG�$�"���´'�.ʃ����>�=);|V����E�ϓƥ��Ex��("�����W{�
��^p���U�O��+�ϙ�7�U�d���]�=z4rkȉ��aķR���\Ӻ��i����&k�� $��p�s�7U��{�逰�*�ޠ��s\4	�kyy'����ǐ�-vv:��ڸQ�nQ)����N0���#&����c���|�@A���P�(�&�-ԣ��U�b��h���/���)����m�j^OP��/�{��a�����Wo�v�^�}��P#�;	T*W�3�t!�*GS,��3��	F�s��"\��~��$�
T��4S(c9��{��\��A����%�  b`*q/�$7�8��5��p�K��R<��nE(�i�x�,p�|���7�\�
<�.Ɩ�e%�<�ި���;���*;����%ه�!*/���TJ6���b���vnS��Í�r�a��U�Ø�,��
VIBI%��&%*�b�8E��/>������8ۙ��x�pY���}l'l<��&��p܎�$����QwC%%����~:�C=�U�m�1�����c�0#�Ư�qF �p�m�Y
:��f�XA'�����?s�ܹs����.�G*�i&Ec�)�y����+(���l@�Go�%N%��R|<�f(��N���ˑ��b?pE1p�4/j����U�f�A���p�j2���D�n�O��^w���KX␤�/���!Y�6et[,!k*?E�܉�[�?����o��M���$惈����n�Z__Ǥ_8sj{{;�M2��vG
l9�t5Jd2�G���!��:݃ơ��no�|��]��Q8�H�	9�J�k����;G�(�^߀��=D�E0P���/��}#r;!A�a�`+���e����dm�t��sK�l�:wnސ��}AEU��ez�b%��	�=��R�d�H���g[�w�/�����~`���\?7�+�癔Q/8��NC�"�EfU=��(r�[)9��k
(�j�H`+sК�XIH�89�_���(G!�T����A',9��������d���^F��h.JNb�He|E+" )>�P��H���N�8���"��94Y�?���X6��Ӌ��nq�{��.N)��NG�'<
#׏e��A��yټ懣�m�$���c�	�Z����шY������W�g� ��L��0���D;$ᶍ(G�&���/F#�(
\ɧ���D2'	acU�3tz�[��P�Ia�����`9�\��_$����,8�L!�H�y�������{ԉ��Y5&S��ʭU��b�_�j�J��!b��q��NA(���+%dV���S�Cy�0�� օ�-�� E�F�-��0Y��l�EL��5�%2	%[M%
�r@1�˾� y�^��n޼IF�d#�xh&NI��� O�w0��U%�=(
�~�B�ף@�a�hB._���TxN�a[T����ed),2�9��8��cr$u:=H��t�)���+S�ΰۧ�/k%��v�V�Hǃ��ݼy����`�Rûvm���ɲ1i��"���=S�)�'9Zh�9���I������U�_����1Y�T��R��n�H*�c��'M��WR��Iu;O��G�gϞ��M9��`D�,�C�rA��K�.dkR"��f�<6's`U�N.\����K|"�:���.��1��'mܐ|b��~�p.	�N�̈��d*��X�vHl�M	�D��<���x4�L��N�/�'�-,ׁP�����n��R&���;6 ��i�ܡ�����v�f�ǰ�q��Ur\,��;]H:8c3�t�_)�KU�F����0�q�c���d�b�%���&�/?8�
��*9 �,�gd��W<��, %�I�e21􅡜��1l��t՘A��Hh¹èJ�O9�[���q%�":�.V����ۘI��(z��3�9� =P���b�1l'�+A;8:�,�rQbq���2�Օ�v}��7nH�|��1&z�����5���jZ��si`�c�sm.a�$�����'��˺��dMm��Q����i;�=��K_�\]�~]�,̥e�766p��B��q^�v,�Ãvvv��T|T����0d8M�\�����:|����������
Ayb��<�UUS�/]�OǙ���@ .ЉQa��>��u�ˀo �ӵ:zÃ�M<E3 �	���t�%�5�1�^:�qf�y�\\�ӟ���u�_�5궚$*	�R��� �W�*�X�l�`1�D+l�e�1��f�϶�Y>{+r��U|3�u�Vp[20��дx�q�(�W�6��"8�#s�nl$�!,[��u:������! �k%J�v�V1v1-�.]�����s���Q�Nw�R��>:���o?7�q�_�=�L�/�HٞB�Lgr� ��(�k�r�H*j�7����糒J)��@���.4ֻ�$@S�� (Ş{�9| *`96��p����Tfv��`���w�B�,GS$-f��[�� ��y�m��TdQ�X��H��7.����㡐ȡ}-~{�]���$le�p��h�	
�M�S�~o�ޕ�9� Ԟ�v<c��Kz�?ֵ�,Q��ȶ�=6́#KF�3I���Z@��f�ˇ`$�<;�l����x��L6S�́����#�6��J'Ӷ5lw;�Oḻ1F�(d_��B!�N�Z�`]�����D�m��pz񧨎I!�DJzh6AR�VS�Z�\%�dNU���>��WkSx��lD,�ۧ-ٜ�َ��{���\��\�3H����h�L�
"���h�����>�1�L�B�G�u�l5����Mܱ7�W�}id�CŰ�h`��\)�-n�5�y E���յ�ѐ�!D����dwg�M���@z�X��L���E1��y�*���p8¦�����d����
1q�N��;�êvR,YR��ųX�λ���V2���Jj���B;I���"�\�R�+2��03������T��R�/�>r�g��F�H�M�!�Ga+
%Z�j�1Eֱ)67v�&�$�I�c������M�~�j�tl��:����}8�=l����B=XP�����v[�T���b?;66v��ln��By� (��v�����vd������C��1�˥�,3$6�4b��"��{`�`���GK�I��s���-�3P�	�n�O������pX�I�3=�,l�n��7$��˹R5����E&��p4
������[dRicnn�V�r�N:���~:�Ȧ��:C2I�e�b��&�ԅ�P���^,_�?K�|��P���
�sc܎S��ͦ�	m[߈d�皭%���*����W�9/$a��55U�2���o�[\[ava�ՙ3g2���x�	7��vI0g�	�=�Y�TN2�DJ*��T�[��-
�B,��ρ؊�o�N@���т����bF(	+��
�rQblt�#��F�*n��!Q
M��8�Na�$2w�����T>�����7�{t�����	������� 
�����Q���h�(�%���$�%DO��bm�X)c$��)�%�
�"?�ȐEQꪬp.=�v�<"��i��k��v�Vc����!�0fff�@q����+AȎѤr�T(%8�{BD���$�q�y�9�i�4
J��|���,��6M�I#ac��֭[^ �)7o��.B���jX�ゆG�[I��4D����]�!�/�k�#l;���1
��E�@4����������	��7R�tM�uJd��{�F\΁�S�/�����`��Q����4Q��l�¬�3G��_o
F+�2'n�n	')@~�s�5�8���@��!�Y�S�$2�9L=�6�=Qe:�d�_a��vkkk7�]�g����O/�R���LW��mH�ވ��D
2�쓜�' +B=Q��e|��Ĕ!f!2�ܼ�:+�=��c�	q<�XC���B��x/��LS*,�1�]�i�e/&�f�������>W��\�j��si�s�,�b`]�v�x��2F�)��T�U'o� ��)CJ��eI9���*����'�8QY��N'\gf���/@3���wT�^�BX��^���T��xr� @�+��2A��9�	K��H�����o��G&�4���
0�>N�mA���Oc��&i��Odw<";��$��c�KKKv��>�Dc[д-/��PRhOC�,�K�V�r� ��#���>`_���[���G��z�ez�����L�pآ���&
4wc8��k,����y{#��c7��!k��4'���ʇ���ؠ��-��|�Eq��a���mo�m��ܧ� q2I�A?�Ts�6-le.Y�މ�x-"�Z�t�|Z��{8KxQ^%J�Ґ>��0�>R�b1�t�y��o�:�d��ho��Ӽ���m|ܛ����X�C9��Ö�c��h��!������-'s����>-�SYA�P [�rEU�{AmB�'y_ ٌ�n[���K݁�ŉ1 �y,����'v�4�}g�@80��iG�/�C"L�x�%�N
��.A��L'_��Y]9�UZ�l"��4���f�6H�5ض�gA�i�{$��c�c.u�ǹй����<8 9cw�%ݍ��=�6�����O�<Wn5l-$w��=�t�"�!G�IU¬i:�{&�J�*
_z����F������Z�����a�:]<�5�N{qJ(	t��l� ^$�9Y
��2�w�սy�6�$@�b���o���%c�N��i�L㱪b���Jfi�XV��+b�\���B�ɣӣ7b�0{t}uuU�d'>����K�.ᖝ���/0V Ykq�h6~ ���� �猻"���&ȩR��Q(�HڭD�~@�;]|=��F��0Í1#������,?��l6�JY��p�L�jr2������;�L��=J%R�b��;���,�'������B%�|}�ǀ3�!�G�"%v�x���
���&��nzzzscԃlM�',	>D�4�q4V���C�-B�@�е=�D(�"G��~�'HC\��TᘢXl܌1�L�ElB�fz6��W���0�W�c��
O�Zx�pZ�����*,M��S!����Ne�m��R��h0<.dї�ݕ��l�"�\##�ؑ�O࠲h�G��g&X�]�tD9���S�$a�@SX�!���
�����z6[�D�d��i�3�h\����nh�&Eϔs�1H��Di/h�N	Y
#6��;�0֨�&�c:7���P0~QO�ǁ(��ǐ/�땫&�Fd-L	��s�^��T���@ V����@�x_�O�x�-��N/�[�q�^t;��3�7L ��b$	B@�9��㒗����V�
�Nڷ�$/19	
ĭu[g���͇ò��8@��x�Pv��_�m�/�"�c��v�R�w���l8�X/�:6`l��,�-�cx�І�iidPȼVSH#1k��qb������`�XQƟ�b�'�6���?��5� {�R�Sl�V�S�j��0%d�n���U�@�¬S�ؖX��=�GD��8;3O�C��XP�B9��4���'�,'��_��$x*Q�emL����Ԁ�5��A�e4UJ2+��]�V�����VP��1L���I�!}ϕ>ض��[^&3���^Н�׬�s(j4�S�N7���@N�t@1v�4LMa]�^�
���X~�{��R�"+dr�����2�.坒iAq\;}�V��d�����_��8�$S�j6C��Cڢt?�T�#	$Ӌ�u�_��)=Ax!����&z ���)�VZYY��7Qx���f'�09��$D=(m���M^���	>꼭#2�{c��b�½�.�<Wo��M�f��&�Hh�2Y�(v�00A5��e�w$l��4ٵZ�6�� �Y��o��I2~!'���$,k#5;� ��
��I��d=v�;B��T�-�cTk��۔T%�|�3�q���!]�:
���6�]�T�Q�BJ�k˚&�3�-��lw����*��X��.��F<���&cI�/&ڇϡJ��=����>}�Z���l]ƨ?X�t"��ZpSb0�MQ��J>1�j�=��I�U�C�xq�|��Ɓ儲j�z܈��/�C����,,Y�S��$�$�r"���G"?�F�JM7�5Y�w�cl�L2�5�R�Q')@t� G�ͤ:t�W�x��^@�jD����gڎ�@+��G�J!	堎Pґ�dNJ�Aʨ ��b�/E����L1�H'����fK�H��tC�W!�e��1o�^`3!����F����9�8m�rx#|��~P�6���q}����g���xr8G�ڂap�#����;߰U���"��ޅq�5�����ҿ��["��`)����b�~h}��a{j�>/"*,�Oȶ��eS�H�B˼�.�<��=�����3��s�t*;;W��k���8�G�Gf���~a{�F*��3;�?�`�X�X!�J�
�)�+_"��F�E
/��_�4B��"���OUxJ�kl!���2�"t�.�#D]��9�Z$����0��c �� �I�
S���[p�u�X ��NB��Fr�Ν��-�O�ht������9���I�b��z��9�Uq>)���GXBgs?ƀw)g�)>�uE���l�� ��!� ��_2A���вt�5n>ay��:
+l���������C�BW|�YE�Ÿ�qx���H<�8��Eśa�H���Z���b��6�1l	r#Sb͑�����4³�=Df<�`	�!W�'���-��g��{�0R2��q�V9���c�4����XN�`�pM{�����"7�jPbiX��B��!f�C���p'3��ax����oD�C"m�ժ�N"����È�B}���Ѐ������̑�ٵX���,o�F�����2$*�����? ���=-9;������P(�2++u�=hl�rߓ�"ްc2:f�BV��\{�2��c��J����-�6��n##�/,��1���;	�)�_Q�MLG��\�\(\ͪe7Vw]N(@�9���؟�e�t�lԉ^SAF�r�Ce8T���;�� ���ʍ��iR�c�c\a��u?U�׭E����U�R�������g�����?w!Q�'��p4P&�p;D���|��c����a�51Y�r�Y;==���?�Nq)�T����e2����6����s�_`�������m�J����Aއc Wx:?�������|i6��w����B�~`����{�^����I������4֐�T�n=?�Z�Z�ɮ�v�;��eCoX���	l���	0�q��޲�v�t1W9�\iU6Hv{����R����Ô�w\��E&>�W�^���zu����.�铓�F���R}1̑Z�u�� � ��
���\·þ�6�V��o2���촰C�k��|�9a��j�"s�Ga�᭡����ᔟ���^�$L���X螛�ky�,e��`�@N_��yL�3Zӥj!"r���-F� �m�9^��L��~��2Y�,~��9�X��Z�A>�V+�}��=g�ݜ��א���F�׹���~�u�8��e[\�~R�g���\��J�����r�	^���n�*��g��%Q[����*�v��;8hὠ��vXŌo�.\�Ҁ�Q������I�����/!Xs��q=�F�˕��u� �T�bWe��Ϲ�f�Z�Ё�F�V�m��x��?�,����G�D�+���Y�s^�K3Xf�a���e�{;$����\��qB�X����T�7!���`�Xy~	6�
{���$۸��h�I>=��E�a:_L�J�
�5 '5���x$LȚ �x��
5U�`�����o�.�d���#C��o�K��s�fG
U�`b�lQ9�WL������$��r��ROֱ�[���:�p���;���%x��,N���7^sUi���Dx�뗯c�G�+ⷷw��!���a���+A�1��j]u.�!��b�dE�����������g���,�#���nU��V��Ӫ�R�7���޾E��Q�B�?����(���T��w�F��*���cL�8[`tcӞ�{��'#V�$%re�U�L*�W)�LW":��^�z���W�Ul6�r8���r�	��C`~ �6K��X��I��͘��<W\4X^_���>
+- ��*`�����D�C�c5����N�N�:ʻ�>�R~���P[J���n��".p:-�������^7�}���Tx�+PNjҮ��:��eU�*#Q���"͌���4 L�Q�l'�z�~9[�6^�Sff%�Ð���<�w�f۱�x�[�O1�xlU��j*��b`�+T�	��^���������͆$s�,A^�`T4xE�RJ�`H1�x5R0\_���J�ụrAΜ�!<?>4�A_���~,���PX3"W��Z[5�׸�됅�>��R�Ep>:Lf�2 �e^7g�5-i�cq�P�p�0=�Z&J�KW	����9WƓV�ҺZ�����	+{B���Jt�c9r1;HɪP��h-��O�=l��W�jW��B�6����$�ͽ�Rb��BEE6)��@��]�ew~��RF-g�d!��X�*�����e����9�	�kQE���-s3�i�^�xe ���Y��J��yuks��j�����o�կ�������վ���:�z�р�%(�!)���^�\����x�Һ�8^.�o����Wi���W�Uk�o����&������ŋR!t����6�gO�9�2��p0(X k��奢�8l�L������T��&�I�-x����햘��)�f0��P�Y> �-[���/q<���)��J�P����qw1+������ �d�%i��i�����s8�>#vk>�݃t�}:�7^�q�q��2ܨѬ�'�0O��f�/#��\�����&���B�j���x�ݛ�VaK���,j�4q����[�f��'�<j�h��97C@I�q�2c��q<�~� �g*��&3K��Ѝ~��	�m6�t�Gx��t4 �}l)G5����zQ����$�b��W��h4!~�Z��i����m��7^߈af����Ů��eP���eH�6L�N��[����ϯ7,�ݽ�B���]��Ul\�g:��Ń�Η�$�`�Xh��W��.��F����j�R�l�|��m�R�7�c��NT`�xE����yA�?:�E���kb��l0��ֳ �����Qߔ�#�s���"�_��p^|�2ãu,`��!���2�����&v�\'M��pD��>��t���a�sT���7œ0��������<��$.B��z���iJ�J����'N�s�l1Ÿ�W�Bq9�K�G�nJ�DxE�\�ά\�����|���aj���Q-�3��Y.ݽ��|��M��9��J�((F^0�^=������<���u��=V�33W����a�Y(���d�{u~���Nmd�#����C�r�ݻG��v,�ا�~:��az�m�����+�������
�Y�oݺ�ŌI*6>Ė5�}kA���^r�m��d���F�>3|���u�Րݰ���2P�˲1�F�V���Z�L1Y|]�[h
�򗘕���6;f�{�����jxl�MQ$��_��_a�������2�4>�C�d+���1 ��=V9A��e�G�������9�N�*0>9>����r��J���M���]�|��ơ@6������e6*/�T���p�erz^�>#�G��ދ����͌��E���2�`�%�ht|x�diF1��#�O6VϤ��5��u߾��&�&�@��Ky����5ǃ����hJ�`��O,J�vC���g���ٔ�XY7�	Kcxʝ�/Ĉ	���#�*���eo
 ��f*�	3Uk����������`{�N�	]xk<�U����&��o3��*^���\�IJ�r�Jba�.��ba���zrq�j��������%�O4��b�>����d,�J5=xB�������ղ�WDF@��r�obr^9}�$�0�j�'ԓ,:���xV^o),*-E�0r�筗̐c;�x0�U�f<򓔇c9m�+Uf�� �� �6�P�l�r�!K���{<σ�wH{^g��nY�F��`ƍ��^��;?��g�6���?;<C��q�����X���O�I��>>���>{�9����_c"�����bo<�� x	C�I�~��̚&5ݽ�9������l�º�S���f�;^�P
ܜ�C�i��� K���[�a�$�lJ�ŝ�� Rx��7W���]��B����~�z�(������d4�����Z�]S)�vw�U���ٳ��h�䮉K�I� ����5���s�^>��0��=�_�tpr�Eu5�L���錒1� ��`��	J��wU��l�UI+kw��Ex�65"6n}ttT����β0���Z��.-��s\��b�'>gD�^1N�x��5W����K��q��pllTai�N��a���� ���qB�o��z���gȈ�s�$�)0|HH�zՀ$�e��byN���]�CDn�B�b='+���q����N��?��`2�io�R|������[/K]Lt��T]^^ˏK�B�]���z�!�XM�z]��1,�J�Q�
f=�[�z��.V�f�R�"N�[Qx2�!��;>�!�,�S�[,B�q;����5n/H?�A�*���0T�6A9A��C�AS�{��]yS� ��~�c�]x�I�y"�
�k�>KS���1��6��7��ڽut��'Ϟ?	� "�~gSS��J��e)�#6S*��J��ӧ�i��.W��#h���\ �BO� g���Z�%r�A��pu:g	�<�����qV(�Q��)_�|�]�*�F#^Q�W+e�=�����냽]�
��v��&�ު��_��-�>Ƙ3���R1k�;���o�F�[�<�r�v�.`xi��F�4������㨈RQ�{�Z�޷�~_���Qi�?_��g�6�ۼ�IgT�������W�W/����I�����Ư8�t4���:0�r�@�����i��e�bB�&V��`���������D	v�}��Y>��7FC��-eV2�Et��\�јT�	�N��Y�lqy|vߝ;w ��^��"�{�>NVy���c�Օ�+E%��I
�_�z�ݞ�.VD{��g�>O d�J��L�"CޗS�w�=%��.���Jz%���͌.Ev�p�+E�-5���u�j%s��0�j�>�Bu��\�\,O%^P0�����"^h	��Uևu���fK�B���%��
��9jL]��(�PD��}<��F�P�IF��ro*r� ���Y�]
>w=�$�w?8$��I���ꈕ��>X����-�5�H��*QDO)~ey�*��P�F��\d����ge+� ��{�V�B��r�/"B��i��
��a��մ���+ ƭm���k�7����)�Q9�
��3��g���1x���o��m�D) ��d�՚շoD���M!��.v�Lq>$&�G~|絛)յ`��5�W���x^ wEnI�Q��sv�8&%�xD����ʣU��BakK���0�p�JkaQ���s�<�`����i�M�0jXِ�t|b��>?[��g�6��1>,�w�K<O�R��ѣG�@�O=7��iݿw��;�>��!����dVt�Y��{�����������z��K^oHlVg�}��˻�_-'�\�Z�bT���V�r����R�5(������,E��x��/^c��� J'M� a`��59ż.[���b�����7�c��!�ð 9o ��(ʋ*n���������G��p���R�7I2�p-��%$�[���&]��ԍ�T���܋8��['�-��B˨La;/!���������Űk�az,������a�_�i������Y�b�
pͦ�ba�}<��-����W����CT�7vvH�8��J�t8�)�+s��`�E���lxL�9Y��E��G��|ڿY3AY����vp���_��c��7u�m��n�χV_(��*Q�?���˗/�3�\��)�s�M������۹��D�R����Yk��b#�R>}���zr�!�;ҵǍ�đl�A"�2%�!�:W��L65$ސ��[L���Ap���E�<!���&o�F��>�h��'��v�����u��4��E��j�Ǚs�m�Q��Z�������B	w:WN�A�v:���E�~%N͋J^�z�u�[����~6
�f��/_<����.S�}?h�X��ƀ��4[����bjP�#&�ɳ��G�>v���B$�_*Gf����.c �P�mR��W��� 'X����z�J4T�����,�׽Y�$���WL�Vk�'???��y�,�熓~��m�+�+��B��e��>!3�'�fϺ����Aod��}'W�ҟ��S�:ƾ/���s,q�U8V�	+"6�l��>ǃ$���s3���[��+�4�֫�O�N�sE*e�3l=虬����]c��������Zb�A�^�(�����F~��Y�� o�&
H(�o~�/�g~�]Y��ܺ
��l��9�s�~ǂ�X����}�嗕J鷿�-N������J�*�̣
����l%�=?>{FV�(b�+c)��Ć�x�u+I+:���y*%vw��L�~��v\Օ�1.���[#�X���V�����#
)7�2���#s�J���cj�Ȩd]G�fSWp][N��r6�a>�_��*�Pl���?>9�Q���?@U�^��:�M���'� [��Ç�#�F����v�麷�����0�\�Ê���f	�1a1�U;+-Q/s��P"Gf>&vR������8q�'�% 4#Q/�޳�兵���Mv���v�e�o:}��w�R��z���?��3��
�q;r�T!0�&^��͋��=��Wx�d�RY���ɍc��Sȩ�U*Fh�ݐ�3�n�z��/�ü@7�^�~���'�)��(ܮT.(7f>���>��e<]
.;�:v�2L�W֒0w�IP+�`R[�<5�c\
V�c�4<��^���6-|����:_�e(�{�&��X��,WM������٩���}��V�k���W�F�A�*�B#����|���	�OZ횸1��3�s�j=ߋ���6�#���X(�O&�=w}�|�uㄯ,q�Rz+�Lpo���CR\[~��]�E��m�M�^�����7MֵJi<�X�3��R��]�E�����o_����;�Gp~��ONns���x����۷������c�W�H�;��\�������r�\��<���b�����؉=7���E�߼`?'aH�������WIJ9,L�y>4��,1������d:��]�͓�w6��F{m恆#��΍�pw�Y�}��V� �C�m0��#h)\�X.�x�V�����Jb%��170�sQ�tgw:�=y���iYb��^n<aZ1�߼�F���`6��*�V�����M�ӳ���v�C����\F;}t�y�a��'�U��*Q>���r>w1D�ْ�3e7`�u��3*$/��yK�=���Z�ǣ~�-W�f���`獑��q����'�s��97�I�;��<+�����I��9T���^m�+��,�E�����A��W3��e�J'[�p��}kԹ�ַO���Y��?���n�*M�Lg�V���~�q�s���[���j�	HĪRxҳ�X�&�Q�VmT��4��j6L�T(�}\���'��a�]^u0�{����Zv�Jܨ�*+o�ը�X��|���V1��x�M��c�B�E�Pf��&W,o,�~��%�b��n��
��Z�Gv�Ŵ��:�f:���<ET2�Dr����޾=��׍��~���';?��C��J��C ������no:���x�����3�� �s�����3/�%�zT)���W��-&��e����]e2����u�$�.R%����v��z������˪V���'��n�By:c9���!q��1IRV��P��/O��߾9#_��������Ha�p�a=��*p�c���Z��1K�����b���Zӱ��'�Z6�`E���F��>���Ƒ�r�M�h���b�)������PEoU&b7ڰ��g��׃�O~��,ep<6ʷ����6K�q��j�L<�[�P��3�d)#���� Ȫx��ɢ��PnJd�]x#�bV�ș N��2�k5��'U$�nKA�'��VJc2����;�^_��r�p�Z(�3U����V�WD\���V`�d����!>\�&y,װ"���h��J�B��r�y�V>�-ޞ���J��z�5
:a�G�`��'2��f��Y�fV���m�ִ�-�P����
K'�̜㍒�8���a��tSs.� ^S6�ZM�|yɖ�2>S�cު���z(p�D�ɱ?�o{Dh���	va�t�`V��d�r%�`���W�,k������
#4/�rS��Bӑ�4eM�֛^�V��1�����~��<`�k|��g_�o^�Ĝ���~B~+��Z/��3���a׳�L��`6��&s��'*j11�[�/�X:@��s��Tڭ#��2�\^��KJ҈	b�q��Ն�:L�b�����Y��O�W��V������YU���/�$빳�Ѻ��Ee;���T�$v��W���}�/_�.��U�.��ǖ��g�2�n�..:Xa�/��Ax�hŖ}��!�o�Ѯ�Q��:�d)a�9!1V.�>���o�b��Ç�a�X�X9??'?k�C�
�I�좵P2�J��V��zV�g��a� �5*�\?73�_�m�%��$VU�"��ƶ�7�O0»�%U��#�LK��WW�;jX��+����AH�7��Ѕ���^zC���{��f�rß�G�GǷ��3��h�\o��`<�̭3> �pE�I2��07*��6��Z+���r�Bӏ�\NNZe�-�6��{�_�z5����Y{����-�,�l.�X���:��k��l�_���0GO��8;{��4רV�$���������;���Qށ9?�xV��[7�����/��-��R��a@-���_k��Y�ǈh)����l�6uq5��� a�f�	�wf(�λ���$��Xz�0��n��b:��j6뮷�m[��H�0,;�6��hH"�%
���I �u�l4(�7�З�����eU�a>�z��:Nb�#k�مE���y+�hpH^�F	�N�5g�ш5qp���{W��p�1aN1
M�����CM\ϺZ��od�A�c�]^R���^!��8��XoU&��+2�5�'��U|:���.+؝��G#5+c*��O�*�}x�P!���n��vY�R���6k4n��:�Zٍ�-��Z����ڸ�A��'�����i��/��>�?�#>��K��j!/��Q����z��
~��>�B!i������a�j[��a��E�c,P�a�CECX�jGh�ْ(�i�w� �gx$|�����0<8���ٳgخ��bv�j���|1��X�gx����j�j���h��lTu�{ڟ���x`U,�L2c��˞z����@��	�AV2��zC�VmV�Օn�p#����l[w��J)y� ��W8M�/�(ƈ�։-��{w����?�z�9���Llnk��&FCE��X��w�m<���;x_�-�W��R87&�<�eQ�a��wzp\_����rA�4�]�}�"�F��^ߝ��%G,\G�L���r�@'\8��r{#Gб���&x�g�e���XkC����$��x��޽�'��O��I�RW&u�ht���7�Nu�Dp�@�kfm/)�.�M�ԋ2+��-����&�!�R�d^��C;x��j��L��ŉuN��˛�to��&�T*�*_�?x8����6����{��_��_�̛�"ɂ�$8A�0x#�$��\��̠S]�toh�,��E��]1�v�д���%|ܿMG$&.���Ȯ��,_'0��Ci|jC�FB[,��J��99��h�hҪWKt���Ï|��fm_pƍ��<���K���˔_�Y����� �2[�t����ϟ��  ��<\l+ܑ��Q��07�QW",k��I��~��߹�޷���Z�/��<�W��`���Ԝ}֚`c<~�h8�^\�3�m���ٔr�w=�ѝ�K�dSH�r��W�9\kz�S�f8�ʙ/��N��5&n>�Y�T0^ŭ��m<�@_�u��`�&�f{��Y����O!�z�A�Ӄ4���$i�guH�ɠ'��!|�	&:g�^�b��55ޔY�R�U�n�
_�\��G*y9:����a��0��2���xC��C�=:�P(���Ϊ�R1����5�Jcf��t8���s��/������ R��<2��2�Br��+a��fċ/�MR�W+�h�Z��6|X7u�Q�6�9��l]�T���}qy�06�;�r�� _�I�t)#L�~�j�٪�	��^������l�x���|\���!W,Dd8򳰘/�KN���=9����u/��P�xٶY��>9fl0��k��sa�������?��$|�p�7<�����c�rH�E֋y��C�!0��}u�����Xc��x<�\r����~|vq�4�E�c��ThMC�B���W�x&�
�W��o����.���	�x��(W�+�R��MV��x����O>�����uf�Ѡ?�2�UW������x<��k�O�s�t����a��:�h4�W��r��6p��sw:�1V�J�9�v�,F���? ���;G4,f��~�����ё
�I������|���|��W�3�qðE[���ܘ3Xg��V�-��W/_�O��~�+�~����XT*c�	_�z���;d�HX,�R��b�}�}�X����C�a&5�jh���+���sf�����d��$�,׉5eY�/<��L���T"��,�O~'�_f)G��U	�:j/!"ޜF�"��U&�JdpA����7V~���Z/J!(���.�V��$���t�zN(����w�.0��k�S��:8��l�˖Ԏ� �S{FD�j�����߬�Ȁ�\����c����WRG����l�8�Ǡu"t���-bs/W�xp�ێP��1����ҖA1b�����l��˧Mc�� \Y�`5�qB�.�'�'��l��+�f�����5�[ܫY���U�"?@	����b���Ș�\¬��sXLer0Y��R5��@��F���Pw�e���:Y�F��X]����l��g�@��8r�Pŏ�sr<�h<�}KHz�%K�F(�ᕽ��Y�����TL#h��&d��9[�) WL��j2h�Y�sy�����[���_�DD��e��8q_�~-L0񡶛�vNIY�!��#Q�����j����{x;qmiH	uX��t�����j�%���2���d���۷vwZo߾bo��B�>6�ް߁=5�W��W-�D�!C=�)
E
��hX.��.�Bʕ�l���Oാy���:�J�_/�py�V�$uJ��5����y�V���cɖ�l26��x4��V�l<�J��t~�0����W/Ɋ�w)��.�d��[�szz��r~��{X,��6.BC���ϱo�>0��vr�6����s���`bh�VGjr�{8���<>>ʲm��9��|�Ҁ­FRw�1�;��!�MN�l�~����p0fe/��&^t�8u���W������W�7�F���f#�v���ɜ�ԫ#Bu�CO���ƫi���釁�LRX��$�1��r)
�>�����ɓNgvz�`�����:>:L�\��@�R�{�D]�պ�d>�l��{QRd�^��4�F#L�%���^���&��4�� `d)ެ����=h�jL���󜘽r��&�$�?�ڌ���:��{�~p:���>?'�b�H��d��;��s�u�V���!�G����m��;�Vwg�����זn�ܹ��_���Bm$�2
s�S�Y���	�·��!�!cs�s|p���\^����ղ�!�^���>箖�J��F�Y�TV�X=D�nSr�H;V4@�И٠�.��-D1�t2����t6�V
,m�������>E�/r�16�45��۷o��}�P��yO�~���]�󃽝٠/�����ep�dk뾱�S��d���2NLIdN\(���~�Y�vwjQD��BTH3���J;�p��"������X��c9�ë�1���"��<x�]��=��>����`��������{b���V���|����],�7g�e�cY��"	W�m�zS�I��g0>�L�V�ZAE�տ̱��9��b>�W)�/��̘'�`�Y-]ն�PUKj�"�`lK�#^�4��\�/�fA+��?A4���+фCu��<��;��bg�)�z����q�f����NW����LC!�]/��Q/�M���2D��?>�u?>0ZC�8�F�+F�no��iXV֨J�թ�Y+���lQ��lO��ᴜu�}�����o�m�.��0&p�Qe0�e��T'���~]�{�	�� 4l�Fj�M!n�q!@�hh�Q}2e:&@p/\��n��
���vrr�S/<��ò�b���fl ���
��������1.W��e������0����_u�Q����ո��-}<*��V\���b7�L����M�����ZKd$��p}r�Û,2%�1p���RV8�}�t�*��
�d��vA�0�|�	X�Z����EB�j�/^(����ۿ��v\|��yc<T�a�8n�\����DP�4<�t�2>��j�m����݃{�e{Y���N��O?m6�q�쁛�Z�l�u͞�:�'���q���+����2�g����`w�Y�wJ�m����O¼wxp�����w����qi��J�V.���h���R{x�.��ۿ"���>��^��;wNo�����Rcž��G�l�IJ���.ߞ�}������˳�3/s�\P)���$���c���6�`��l<����_�&�7��^6�!��p؁R�l|l�ղ�e_bQ��F�Z)_���|!�%�n�#F^�R���C��b4�޽ß�x��Oom�!�p�f�Ms>{��!�A���dS�n��t|��}������ևA΅�X����f��-���`p�j�,20q���ށ��Ӟ��!��+3w�v�m��������C���G��Ţ_e����횩���`�`���g�r�nV��A�~�����c熑[*�aa�~����NN��[�����a)��4���F�|��-�],�Z��|ɚ5]�{S��>�OҺ*��Ә��ao<��Np�z�p�j͌4[>緛�;�O߽�|��Y�R�uBFwǁ��n6�������V�q�ֶQ�zb�d�x�%ĶŚ�>�F�:����Ʌޭ�#���~��|!��O�v�p����h��p;�5S�'��@�tY�0Z���һV�.�TT�Va[\x���ӹ�N�iCJ*�T$�	����M�j��ֳ�9{u������\�U�0��^-���;�v�b��fW6��ݾн�	��V"��kk��R#Vv�wv����֙���j���+���>�������zFh �}ܾs/x~��e"��R1�4��tx��[�R-Z/�m!����`�o�:aqeH�-Z�L��k����KcAJ�c��~j��� _�Z#q��^̰UXhm}/1R��R����9�h�(o��
��_J�:~U(��YF�:��p����7����x/��wE[�W��^j �5�v6p��cY�{9��a@�@���<��?���-�쥥�+W-��=�)��h@�OboW�&ZLVC �F�8���5�t	�(��=�����|�_��U)�B���V�a�j�i�w������+�*���(2�oz��j
m�Ԕ� L?=LH�d���9 m�S!ʙmzaz��T�W��a��j�& �W����q����O>�W�Eu�#�hK� �\�_{�����B����.���wW��r�ؐ'p������r���	�����9���-P�/5?W�DO�QA .q��� C��~����6��F�f^��x(R�^[�Ɗf\�"1!XV��I�#H�
��pk����E�@9��ve�w�#}��D���kȯ���^'Т���<����DE�Vi"p�R�`�ɔ���n)���N3x/e�p#e �ɳ��*�*Hf��|��=2I���t��=zxO�Xd>�Ǽ�A'Y������c�J����Wm� ��"�B�U(USV���=l�ϟ���a����	�z���rƨK�����.��q�Y�ɨ��M۬Z*^\��#����&��b^(Q�%醄�aXb������xe����e8 I����r1�lZ��ڶ�B�-��K��l�мD���!6�`�7�*�*H%@����j��i���K��ao���}쎷�΄��^�����q/޾��\f	�9?�nرA���.�s;�݃ý�`0�� ��n��v���w�\d
�\��&]/+�6R������zY-�i16q�QA�Ü�`�}��w�Vψ� V�h�U���S��ܹ3����]v`��F����3�޺��(�������!W`�8������!���nk2	F�N!�@m���2�M�����~n�\�;;��utT �	���r��jU��o�ś�;g�HWk�Q����-����2Q2�۸�b�
������/������f���^��GA_.I%@��}��lL#�L�"x
*Z���X��j�V�aX��l	y��n��w�޽O�ٲݨÅ5l-m��2,�d�X~ �?s�d��NJ7�ZOc�W��|>(��������6^-��D� W��P�)�m���e/�u�.�7��(ψ����7�M�H��.<�l�̧����ɦ��x�Ǉ�V#|t$��R	���LV��C�����%Ƨ�t�h}#Q` \���j5g��}l�2ڶ[�|�dɲ\*��L���L�am�Z�w�Y�^,[$ʓ�mY��X ��ᵯ���Q�:�������Q��
U�p1X��p�+�U�E6؂u�����,У�c�����V%�dQ�����{�����p�Z�'��b�N�:@\,�g���dX�0�e�F5�l>�1#r���z�.r��ˬS��[-�F0�<�,Jȇ���U2�*�����Һ��.7�jd��~�����X��7ų�Q�l� W(ARK��D�����}��w� �5ohN�Q�E���<��_��x�Թ��
O�a�+[Y�"���~�����!G̒�i<�r|�zί����pYu�T��R	C�֒/^7e�b���e�p����>�lpB�X7Y\�/2������l��a�����ᾨ��14Z��fK�>�<ȗ�P���r��Y�������M���b��9��[|�[e�
�����e����l"�����9�UD,��ڼ[�F#�R��cp[�yU�3�������[�*^���1���$]rF��+�[1	��k���j�U�I�P�w�C�>3F��:H���f�����V�^�6ǔ�C|���
px�.�(O�nT���[�e�y����W'>(��{��-3K�)\��������G��ͮ[�R�c�#�������f�u�֭��KHCŎ��p��)Pq�qwͦ�Y�6�<bI��rQ��*[�$��ce2oQ.��8�?�t�^Η� ���*�j��*�`���[�&.�%�^�\"i�hL�6,MHlgk���/p^�:����c���lB+lw��x8¯���K߽#�3�k��{��I�|t{sց��yl����}����|3���ö����A��i��2��n�V��o�w��1�j���	�P����"�6�������b��j�@>y��
�H���@�d:#�G>
���d|���=Vo��ˤ����IL�m�6+d��'*d��d��N#3���Re�=TJ�����$�n���:d�Y������y粧C�gݫ��!���ͶF��?>a�w��g;���3g���c��U���.��s�f�m�f�ۂ1�e��^]��ӽ�]��`�ԣ���o^��	�Y�ݙ��|ׁ���8y;8�Ӷ�5��L�XKp�`���|�z��`fLy�����/vZm���β��|����6f�tjt��a��d:`a$�9���|5x�j�wՁ������G�n�{��-	"Zg�I�m����\1�����l�V�+s�ht;��Ņ�l6[��{Y�^M�;��o�>9�a� ���+�`׌z]�f����>�uߖ	�Cpbi��$<��lG���J�v@�GP��h�Pݽw�{��dx��v�,��
a�u�ƪ�^�Z��1#�T�X�Ǉm�L
/����ޱ6�MR�Xd�c��(�&�2s�kH�V�d��C>���#P���M�?��uj�����(J!O����P1P5V���ꫯ�m-/U-�8����(�k^X;��vY�C���	���B� �B��ԇs��ح6II����IsCZD��T�	��D�?|�P%���_��.סH��[����
E#������ma
E�~�=�a��s9��[6]%f�&n�q�y�KU�O~��G�1'u�yN�Pb�%d�*��H�a��5���U��T����_~����i�{!/J�*�V:�X#c�*W�~Y�r[Z�]=�D�$��cBA�ѪX��Z��j���x����['G"V�U�T~Y�#�M�����}-����5�#\�Eu�d��k��<0C%F�5�f�/��^��,}�O&�`�^�T7*D��+� �`�)��YF8Ug����ĭ=ǽik�K��P�t~���hy��7?@�,Zn�CNo΄�xS`Q����W���:Q��i�sSc�=���ޱ �^3����%�cc6�0JM�X6w�03������W>���1bd�'�u��تX0��N����6y��J������?� xl~[/j�������:�y&�����C��Iﭚd�|�d��:>Z��GX}��	� s��[�}�H\'g	������c���|ֽ:�o�X�0�R�[�ۈW��h�k����uj�x:��9ڻ�7$]p��r��R6���.)��]�$�nt��ˎ��4لA����x�������^
x���G��	�V�X8���a�ՊN=nU+�+�ORW�nXP(1�^�װ%^�y!�@��!���^���\y���A��c���|�����2C5��0N`5�ƭ��ݗ��[��r�~/�[���\�A�z�BI��QXI7��|Ш�6���*��T(ϧ�mF0�-$*~�W7l�o��1�^;:�i2�^l��sE
�-�w��������q>(%����M�,�I�/�����jc�X�UN�ւ��Z��s&���S{:�¹�^v���R)V!�&��d4�R<�4�~p�%�Q*���e&�ݜ/foޜ���������d's�]6��m^�dm���q7�M����z�֛3�,�ш9��p��Qa:�����k�H�b�V�dI��C"�!RG�>��:�;���w�o��R��kӁd���rU���X�u�I���YP(�)q�o߾!	
���Z�W��RDe'��Nt2��1I�9�Ž�1��`���Z:d�fluy�:�J�ԍ���HXs�Ra����b!����Rb�fm.xQ�n�I*L/�'��3������m{�o��mU�2ۢW�6�p�WK���Z�R�I��"�a�-|����0!�	mk�y�r>��U������;��u�
*��އQ$ˢ�몌bh:��%~�V�L�C�8sd���D�Z8��'yI�*�F�肈@��� -��N�z������n'�Y�{�]��ap��/U��P'�6�Սs3�a�ы�zr̚�6�߯�^c��۷oC��^����wZm��ܜ�=-�誸�	�̗{�Xy�W����D�S�x�[��G�nZA1(�N�����׿�5N�߃1g��#�)�@A@��6��j*� C���L29������vTm<D@�����XQ���"�$?U�
����s>y�Dn���j��hNa��@�����g��	�Z1E>���{��K5V��"��RP¹��u�F,�tuS���%F�eA�IL��2:�� �+˚f�L�K�l�Lh"�I���G|W{���l�T���_Q��s����>F�_�
����xj-��6�0PN� nT[���x�ҳñ��MO@Q`#,�g���-��To�����˧��b�.2\>+3fs�.�fTA�A
�=��Y֭9��Ð��&��R�d����o���'�ݏ?�62��g��1�������_��Q�?��?}�W8�G�X�nW����V���ջM2�w�:�m���;�����seغp�'0B���������j�N��2s�1L׀\���mg�+��;�V���c���d���t�jeدp~<\�< ���~�Cp�EW�>"
�Z�
*�W�(&��߱m�X�{����^��ۦ~�jĜ�j�c%�G�{��L� _Z%�j�M�0)�s.��,�b5����$�m������߬g;�g�뇝��z�q��uc��n1)�c#��`�\$�y�J{�K_?|T(�������fq�m� r=ɇ��g��{�v��Ϲ�|�����s��[{��Y.g�Gߍ&3"~n��z���g�l�I7�ń�I_{���;���/�������QP�`:f3�̚�BV�̾6j]�'�6�;�-�Wk�m�13�m��v� �xO������Czl�z9[^fE�]b$7�v
��(doJx,x�˷oT���,���P)����m(��)llȶ�n',�?|��{����pU��p�9�K�f�s�[ͭ5ޗ��n��ًד!e�z:_NG��P~9�nZ-G0�	�"�g3l���5�b>����$^��%�<�������R���v�Z棠X.tz�.�o��b61�{�;�\FBN"�$aRz6�E�J��N���Uje����M�p��c{�M�Fy�X(��8]�OvZ|�{IVcC�r�Z�֓�z�Zt6����n>��qx�螵�##�]�F�Z��f�W�缏Jy~ Q��]��}�'�=��$�#;>�����pI�얅�;;'�;lT)��l.+�݌�8��b7�˫�HC�`﭅�`��riB����,l+� 9��2�w,��ȾwFͭU��SEυP�-R�a����Dd�L��K���7�aW$#,�A��b���j)�^��^�xqpx��իW֏�,!���1��r���f�ӪU�y�g1�k��_����!
��'Że��[��7��n!nWA��a�XߔZ�����6� CI��,4��G;�������'��М3����S텬c�ƛ"|�4Eo�믿��u�1|�؜T���y�������p�*���OK��*�5�ܔ��{�RQ�L(5���h��l[[Q"Ay,�W�%�`n��76��	jGQ�mb.��l.�M�$y-x��|5�?�3���R��Q���Y���$IE2&߅l�,H"� �o��ֳ��|ny0��m�j,�����d��^rUr�,�|&�t̩�ԃO��z�MV*js)$�t��l�5��1�1��:*�d��ke<�VJ�=��Z	����\%3DQ�*P������4p~9���Em\J0�g���K�ZQ�0�z�%�j�!*��� p�iY3U{�gJH��A�\���ϟ�x��9�B1|��)9�Hx��� m<Z��O�F~��<,&j�7,v5[L�ݻ��Z��XO&w�?:==�CP��.P���$ �z�![xƒ }��v��8	�qH���hش���el�M������!�`�Auzx�,	|��E��ſ��#z���j�z1d_�ٌ��ɦ׹���>C?���[K�j����U��@�(Rz8�B=,���r��+�v�������p���ZO'���V�ls����s�d=�����8^���潓�O��g����M�ɜx}���;'�v�x�Tz����A ��C|����-���׽mꦛB��"�\���v5�B!�|��A1�x�ӣӜ�K�i�����5���@�� �\Ԭ4��7�Ȗ�\��4�/;�!�+fC����갽�(Uަ�xПF�����z�I�y�m�v�j�٩i�����b��v����Q~�AR�L�+`��V�z2f�3��"����d:zN��'�^jըg�~����fnP,�=w5������n���`س̪��tu���t:��
��K�Lk����b�7�x�֔ޢC_&8���Q����44��Xt��R[��j6�G!�0���ծ���Ҫ����Ѕ�Q�UşF �_��t��6�鉛_����nC��(�T��K���OXD�kc�/�uE�að�����xDd$��̧�뒔t�� f�xk��}G+�ؖ<��~�)	2�w_�"���>|���|�����$b���oH��j5�⍕"V	�W��v��|��8�7�cc�s�{��z�o.	?~��G<��yp9xSQ�Ii4R
jgC�bzNU/E��'������56ג	�[�M��*'&�ؾ"�wǠA0�'����ׯ��24*iw-���{O�P�5��i��7��R��OK�Hx5`ǭ1Ԣ4�Y;n��e����'�D�!2~1�"���)9a����Sͫ@�G����Z�\���m8�A6;nF����F���ע�]y����;�MT�x�|9=1ۅ�DxM�Z)+�j�/Q�v�W��Y�� 
P�>4P�
�*�#b4��e|k��e)h��wĪ2le���l��߾�O�;�%Z�H=c��l:Q���`޾}�I��6�΍�Z
saT(95�v�	Fi�nx�~9��/j������M�k���ރa9����v��l
|ϐ�,��>9=ܫ6-m������;�v��\Ȭ�H��/[��t�Y_up������$iB��2-���I��F�O?�W؃���;�Cx z��U����P��x���\�$�P1{�N�6�LÖwr�B�;�)����d��P#�y���:>9��&dg��ˋw��Nռx�)�m!�Ǔ��Uw�ĭ�܅Y�Q.w���M�F��,ϟ_��6�U#6�@/7�{�K�
}�$`�I!�rRK��j��f����|̾0i���_LoWFR����:>"���k4ɶ��|[N*��oV^���4��݋��N��z�~�
�J��y>����br��F�^��_��Yv00��aw�6�<�0h��t�l���ڋ�����_}���_}~���!z����a�0�8c�;�ΞO�Ũ�o�y/�+������b���ċ�_-�ƘD��fp$+*���e16�ը�=?���1�\K\6iLp`��G���@���*
��J���u��{3:�cP+�޺ꢱ��3�Z�Zβ�BL�����&X{ۍ�ɒ��y�eۨj�vH��2dTb'�x���بְAf�	0�W��p(ŽF
��2��K��s���рy���81׹qo�>���jNv��ѱ>������!��{+a�y�55i(�~�7�52���1�*~9������v.�]� �� ��!�<ҋ���$Z�D9�VqX����w]�ŋPAϟ?�E}�T�*cJQWkY����w��~�E�>�Է��ē,��C���
��pX`�DB{oO}���zZ�𡳂�������2��L�$���/��"�	�b���կ~���|wo�i�P��|������ D /������堈,�ت7`�x��;��+��o�d�5Ox��s��K�#e5-z>P!�;�R*Ygb��i��c�b$�%�'��O�ja��
j���t�����P�����!�lg�QUk���bv:}�������G�*M�ߠRL��
p�f_�&�XnY�i����y��w�L��B�Z0p��h�ů���=���n�����͝*Z4�b��K���o	�GȲ�T�����:c �[��bB����:��R]��7tm��T���USHu�-tN�
]�!�����	1��Xe"xka����掦^�887����ᗿv��6�x�ي�q<u �Ü��$��P���?BX޹}c�6@'I�I�Y
ww��T����I��v[�����&���sy��#l9K�N�/�M��j�us�܅}���80
���eG!po����B�r9^M��r��*�RH:� ��q7n��mV篞wߝ�@ܟ�'�*���u����4^�x���O��ý�lb,�W��{�-��b>�Nz0�
���������-^<�����^o��v����)NN!.�F���4��j|9�1��j����К�$	�̙O�@���w!�,G^�<y���<�N�+�z��뜿�e�{G3?���쀼�U# �>8�쀏սz���ŨZ	�a��j���f�V��{�Oa�b�ڻ{���X,��ܽw��u����'���J�clK��N�����P�hV�����'��+报��m�\c�,N�Z�Z^��K�1�o޼����6K��;�}T���u<aIZ��׆��j�8��k��x6����\���,���6���j��x�G}��r�m�U�u^��Ƈ�-��b˺p���7��s�FV�SW����p��y�#?w�Ήp�A����~	�k���z��S�띛��d<��W.�򋘩8v�E����pI�0��QW8���f�l�����9	�g�n5�Q��ݗ;�����tgͱ����U�W��m�9�h��/�/j�/7�Hv�gl-N�Hյ�"��7�v|\��p�YS+�����jLJ�N�-T�[�F ,�+�!�_�~MH�u)�-,�ϯ���>�]�j~��.w�n�-�g�Z]��j��ꖌ'd�`y]�m��t�Ť+n���C������b��bZ��P䦽�@=��T�0�4�X�pq<�~�%��7�|������9#�bZ��:��!�h�X	�bt�=*��?��?ʍ�s�����e�ʪo��Q����㎸��O��3�7W�(��ݻw� S�!�@��d[�(��S� f���.�ݿ���{��q�|!���Wp/Qf�kK����W�,�5�h�����x�� ��L��kh�L6���������+��U�7���]Y�3��WɠƂQ�A�Q�jU�����wW�E��.fT�9x,�X�n���u���g�&��Hc�8�g�Th"�K�)x}��,�3�d������)�=�b�g���Ņu���[�+6�D�A��ť$�₻�YI�0o��6N�a�����q%/���e���`�_��t��6����!2K߻.��b����z�e)�`�Y�X�ySo4ae��-�Po6��*���4[�Z�8q��j�ޭWJ��>Aw�k��׿�u޾Y}��#�aR�SF' X��L��vH���Z���U�����w�}G�i�Q�;A�:٭���~��xZ�<=j�Ǥ%JW3��}�5����O�zW��v\�V�Tw��D���e�R�n}��ޫsu����k���;w8�8=��l���\ƞ�U��V��j�JV��r]�7�ή`����y��׹|��?\u^���_���@�sH����
�AΣG��H@��n�އДt��adCP���r�x��F�wp~�E�xF&���n�:�W �j������$o���������u�TyWw���E�Bo�?�u��2�s0&s�ڟ�?�u޾{-1WV��l�n��ň-��.�X����ߕ��BM��i���D~*A���$|��i�ܖ�6�0<�#OEJN�ز�qj�b���|�U��7�(�$��v�73�m)��R�c����wO����`��b��z�o��5R�jU-tn���L6v���?]|`��I&��ݯ~Xc*��ʮ��ʵ�Oì\����F�����o�"���������Mz����ŹE{���ٴ���5&/s�/H�Iy�޽{��%e���j�Tl\����ZA�?�x[�a�^����k����`����o�p�Y��>L2��3��`8	�?o'���m�7P7�E�����#gc&����7�y�P߯�\L-�R��gkY�yu�|�mCM��C�l�4b굦&�!�fc�>|@�b$N�9�#'W�k�&^��HJg��ę�n4GTB��?�񝕄\��!X�,Z�U3�� �nQ��D+�,_7���"�3����ܠ�j�t�2�1�tI�� n�֎D�M��VG���0|�v�8(�t��z~箜J��v$lC�����#5��O�>I�d�	��V�H)�SB�Hc��	Q����j�w�pߒc����-��� I'a�!|�-R[7��S.Rd�y��m�=�z�>����(�"��8�/�Z�Qa�����8�y�I�B� t�4d!d�V�����m��8�Q�FÈL�@�F4{�'6e&�b(�B}fn�9��9#��6�+���$6���}�`s����U}�:ɋETy�ٗ�Ua��5� &t�h^����-R�+UY�a/�C�Tq�����gmy�>��ͯ����jN�g;Uj
7����?~�Rq6����Y�/.�������as����Cw�Z��3�����;�nό���2-6�?�h��W�F�#35�Y�=K�k5Z��y���i���B i���j|�ZVa(��ͻ��ڶ�rD��k�_�zg���M����j}�j ��|u���H7(��L� ̀��5`G��*ݓfo|��2/�2<�+��'g�=.#;�U��R���B@��x�y��s��G*ۭ�7R|f��G�߶�T;"�G	����.~}�7�P�e�X%O����������$��}���m�3_�����ЪK�Ua��E*0���C\���P���e������Ӿ���Il<s��$ުx���D�f1P�|p��R�{+�g��@�|��_bl�A�Z.����= ���Ƥ9��#]5���x�XVx)H��>.�J>���#blۙ��ԉ{ ̟}��[g2w��Zm�R�!vyMs3L��}��GoIn`� �+.���]9�Jd_}cn�K9�C�Ƽr �-m�5P,���m�#�e�
�X?` �am���C�R���,l5 ŲZIڪZ5�9�ل�,n9���!��F�٠�E�'-W���:c��סY�38[W�����O����2�|�����0i)�o-[����3�[jŭ��J�s"��Z���'6/Di�A���R�j=�TيcY��Y��Il�E���q�!�"m����<F���[<���,���-�J;$RR�e�d��yOh9�^N���<�+�Y]�/c��=����A�,�C�\�8O�����ߪ����I��Ž�|�nw�+A��;�Y,Φә����n��P''�ưig�ћ�Z��r�fs��]ׅҧ�ö7����T'��6��!����|�~�XG�U�2̒Ca�p��FSOvF��jZs �Q�l({�dk4h�WDL/���e|-�.kc�,�L��<���I/�L.�.�a��S�P�ܡS�~6��̦�i�VƑՔ��;U�iS&������%�bR������JoU����L��u}ȯ�E�Y��*׃�u�%g�9��Ec��A�7G����r"��c� D`8�"��k�g��+m�4�&�L��/��"�ʟ\/�Nb�[���σ�$*�(\�O�)
<09k7+Ț��X�o.Gf��3�3�ȷ<𜊋`3q�n��K��TB&���< ���f������C��·w�崸��U�sz���hi�}UB"�ꠀb+��V+(jr�@��`��*'g���{�5�6��K�� SZ��^3
.Ǻ0�|�
)[̥=gN�L��g��
���S_G�[�:{�q�(E�m�N ���9ˋC8��n��@lq�i#��Q-ǺV/$ڈMRAݳhG���"������{H�;���_ք0L��I>��:�⫏�ߝ$�˶��x�6�����y��fc�k�����T)�υ)�Z#�A�5(ɛ�Gw���唌/�%V���N�ۮm#�Q�:{S`Xg&��3�hЧ�ڨ����ꨯj@S�k�l]Fn��x�0.Vx�^�A��X$�'���˰������*-�2�c��\1$�q�V�k�(�9o"�	�|B��B�hQ�c�p\����c����_��a81'��eꆲ�������fG5n�O-!W[i8�fH#�
.��7E]����x_*�8ɬ�>��Fᾤ�*i�">�*���ڠr:BD�ى�HS��kB�:�TYW`��g�9��ܛֻ"o�����
1�hۑ^�a#�Y�}�X���E�=���D��+���S�$6��=ef}J�h�7��,��#�9��Ȋ�7W���6����QS���T��r>�˛v���&6
ko��!j�6����m�p�΃�B�f]u���tR@&�5�"p���_	�y
�0���=Z�v@� u> p�$[�t��5?�'VĘ\ѻ8��-�w�	H��/Tf"7,F܎��I��n�S��`�_��{[;鵊���c�T�~�C9��~ʩ�2��W&�H��)U�<�f�bYl�d�qSb��k���z��%Y���w��e�47��T��"��~�ª�����Rو��Ij/���c�(���    IEND�B`�PK
     uK\�6�P�L  �L  /   images/8fef4bdb-224a-4a07-91a3-222e74c30575.png�PNG

   IHDR   d   i   C�   	pHYs  .#  .#x�?v  �eXIfII*         2       D   i�    O       NIKON CORPORATION NIKON D800  "�       '�    d    �    0230�       �        	�       ��    40  ��    40  �        �    <   �        	�        
�        ��    �  ��    �  �    �  �    �  �
    �  �    �  �
    �  �    �  
�    �  �    �  1�    �  4�    �         �         2016:09:27 09:37:50 2016:09:27 09:37:50 Тt @B O� @B            
   X  
         3064640 60.0 mm f/2.8 �/�  �iTXtXML:com.adobe.xmp     <?xpacket begin='﻿' id='W5M0MpCehiHzreSzNTczkc9d'?>
<x:xmpmeta xmlns:x="adobe:ns:meta/"><rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"><rdf:Description rdf:about="uuid:faf5bdd5-ba3d-11da-ad31-d33d75182f1b" xmlns:exifEX="http://cipa.jp/exif/1.0/"><exifEX:BodySerialNumber>3064640</exifEX:BodySerialNumber><exifEX:LensModel>60.0 mm f/2.8</exifEX:LensModel></rdf:Description><rdf:Description rdf:about="uuid:faf5bdd5-ba3d-11da-ad31-d33d75182f1b" xmlns:MicrosoftPhoto="http://ns.microsoft.com/photo/1.0/"><MicrosoftPhoto:CameraSerialNumber>3064640</MicrosoftPhoto:CameraSerialNumber><MicrosoftPhoto:LensModel>60.0 mm f/2.8</MicrosoftPhoto:LensModel></rdf:Description><rdf:Description rdf:about="uuid:faf5bdd5-ba3d-11da-ad31-d33d75182f1b" xmlns:exif="http://ns.adobe.com/exif/1.0/"><exif:DateTimeOriginal>2016-09-27T09:37:50.400</exif:DateTimeOriginal></rdf:Description></rdf:RDF></x:xmpmeta>
                                                                                                    
                                                                                                    
                                                      <?xpacket end='w'?>H��?  E�IDATx��i�%וÉy�S�YU�*�\��AEJ-�Ւ�0�ۀ���b<<���b�����?��v�%Xj��E���\E�\�s�c�#�ڑE�C&���n�p���2�g���^k�}�eM�p�׿���ן���>���$֘:�?����L�h�����jC��9������B���\EQp�9^�%k4�G��9A�������L��~���e� 
�򲄱��,"�BQ�E��M#�����!c�e	c�u�9���+���/�B��հ���0�(�ì��a��U�c.$�b�g|]~�����a��E���74,��U�O�L���� MSU�7Lb��Ԓv��-&��*
|�bA��Q �M�SEQp�{���?Tu}�����A���$���75�_�X�t������G��x2����k,��1�DU�4K`Ybu	k�i�y�1�c�	Y���)Y��6=w�1/\=3��}�Բ�,�
� �
�/�4S5=��
 'ҔT47�S���*/H��Ƒ p�a��������܂c9x��p�_�X��Ś�lr����]�y����^��5���O�5��}�n/�Q8��1��+��"c��N'SM�a>�+�2�f9�ō�Lb�_߶tu~i9��,Mj�L]3&��&�"�UUN�OS��$����84Mγ̟L�]��Tu�(Rǵs����ٳg��X,`z�����ͭ�+W�^~���h�aQT}�K�̒,oD&"���,)R�����B�ZPU*e�cTe�!���dY�3X��4Sٶ��,�i�T�@��%��4e΋�ך	��(I�ϳ���IX��G��Q�d�h�o�I{�篯�.�;w��K�<q�2��1c}*�l�n����?}��ݡ��Qrą�dAd�Φ�e�M�8�Df�.K�uI�S�9n�Wu&/Ve�ĉ�)yٔe��� ���i��slK�a�ቻ膖�YE�,&�fb�G`�jG��T%��0Y+k���2��FM��qu���[믿���_x�+O�?ah�߀�~e�(�.���_��x�FS�=(�����6tX�d���'��)L���$�Q������.�4h��aK����Լ�����|# ���1@�u;@7۶K�YcUi���	��ɒfXeY�3o��jZ&������b���Ta��LL��p����[��y��3O=����A�V�:��77~�����Hy����M�O��*�Q��1rY-d&y�'aN���t4B��@a��Wp��9�	�\5���ZU���U�1�(Q8�#XF�Q#������XNP��9�]���u'�����"����w�7b&I�6dF��,�WH�LL�������lܼ~�;����.*����x��?���z����A�Ҽ������1���������0L(��@�LSW���quE����/��NR��� 9�f���<�E��8��GC�1Q�� Ci�JL�ˌ���x<I�2P�F�GԼ�����*�Q��RlY&C`�\�0�@\g%#��Y���z��{x�o|c��/?�؝��XUS�����_���=QR i
�d�J$�I����좬�3+J&3ϛ�<���HJIV��e�l(�q0�,%Q����x%�j2�a��h8P1�כM��Q����0�O��TV �u\ �d:"^�<Qb]�;KbiD��1pO�2-r���<c�XD*��#KS�r���5���~��7�;��Π7�����O~���t��:P�=��ͣ��^����p2Sm6��)�ܒ$�(�x�����Ξ����LΒTKALS'd1F��P�d0�Cʇ���1-kw44E��S�V P���N'����t�B8WYC�&�Ț� ����Ɣ�~����Gԗ#�����Ԃ���� �Y��/��|�������`�7޼����'����B�v����~�DXB���1׊�O���A����́�e�8���qI�($��D$�x^p�8�e)�a%��J`R���?���D�0�'FRTI�UR�L
�#�Xd�skLd�|�� � I��^L�Hߠ�pu]��RP���3-�/��s�o����ݹ/d�w�\��ßn��"x����1����.�	��{w�Hf����0�d<�#Fj�&��I��Lcȳ�U��w�Π��J�"Ї�v{-&�Vղ���)C!��^Y�P/�<��;�8<\�X�����5U2-�%
�&�D�����>%s
!rp���0�4�~����L����,���667���1�%N��{���I���|y�,2m<��k�E�WT/�dO��GLBOQd�h�<KJ����@��*��aP]��*O਀m���W��b��$���)�e����a3� Љ�g��v��eV�m�$#�:�R��'����+�Is�0Ei���t�& od� 1
#���� �a����+�N���=G��(ca���W�v�v	��i!k��d���.\��5gZ:R~F�m�vB^ z���&#^�g�t���hWy��a�V�u�e�;��|���'���Y�!{�&
y]��ʶ���eS;�	���.��JA�eE��(��)�2IJ�K�jԊ$c�L�û<�ʩ��x�Ad��Y��ZP�v�g?�������?t���Yc]�����\�A�d�3b(
����>�@m��PQu�&4J"8m�G�U���Z���h�&ɺ�X6`l2�Y�2�� �2�ۃB܁��si���`��-2��1&`n`��0�^3t0N��AKa|b0HJUw3M��Q���-ɚ
*�@�8�z�RC�
�-@Ai��a	"XH2�*��歍W^}}yq����Y�����/o��D�� ~��H���1�%kT<	�Z�P�#��"���^����ϲ���,��:*�&3�vd/L ���@��A�"�R(�\CC@t�pj|�$KKC��1(b����T۶�~,�@��Y�� UD�Jd�(�_��A��*�eAs�p���F��=k�|E����gY
��z���K7�|������N���� /	B��A���CUVq�������d�<7�E����>U�W]C��-�����w]@�xD�(�5L�*����($2%)<$�,} \Q��G�E��ABi��h}@\�(H�8ઊ*�*�ZR�$�VH��$�ȷ���� �v� �j�����u�!UAȦ	�
�����}���O;����o��d����c�Y&x'fA)�,�0�C��@�c�0-���V��l7�(�^')A�4n�AT��'LB�6н�H�%>ן��0^�TbuQ7��?5 r �@���eG�4��t9��kd�l2u�d&��IĀ����@xڲ�2�_r-w���_¡iᣪ�k��T�)8#$R�� ��-��4������`^l�����ݼ���_TbF��0��A��"Pɨ����X��G�@6+���y�8K�p��\]lj�]׀��	��تHݟ��&MR�%:3)~�q��T����e��ku������(v�U*����r0*�
"�s����v)����	�%���|��a`&pC��)�������ĸ� ��1(8F�����<i�?�o,��k�o�pQ��6�h��m�c^W &�ͦ������ ���z�iڽ�a�ӛMa�A�gg��f~�Ӷ,�"1o�#�����<M�Ӂp�^��4���2�Lp
�#ܟÄ��:��.K�q>�M��Λ$.�� �a�L����y�8�7�D��Q` ��& +�r@�$�e}^�:E���/LG�:�n�om�n���xkgg���C��y�P�(2t.��8���̏a�k�o_[�*:����T�˼i�{�x�C-;r���e~T�j��K�c^7���K4�ȁYi�(��!�����R^-t�� E�&������<Ơ��	����'Tƒ�Џ0X*37<�E�fä�GrA܁�����U>�\H�a q�wB9�_����ݷ6�6�7Ν>��ë��w� t{�'��T�aM�HDU��C���1r<}p�.�,z`T���weMį���@�8᪬��8�Qhc~�A�x�Pr��ڊ]�� 0uǱ�WU�K}���o��oA��<����g��E���*�qI5[��"�v���	d�l0NX0	2 �������B���/�iD��������q��h}}݃��kP������t�Ts�$
��	4�Q�(44�?�,,u]�Z��8��,��	|��Ԅ���v���+���t[�<&J׮�&Rz��`0��_���h�I� �TTC���� H�r��8���k ��[��TJlcK�2��F�����d*/�����/����IS��l�
�,)�e�qLҲ,	UeE���w6�[�,���oՂ�
�Q�۶��i�k��μ)tg��?va�o>p|���S��.����:�ůi���/�w�}M(�,� e4M�(�"���Wb
r'\!��{D:��-[���Àv�Y=�������>���+6�(��~���@�����G�
�
x~���rױ��
cPVq:�!\�j�y�rD��1�v�>�YD^�-7L��;{����]Z��q��EɪcY��կ���WFcgg��f�;D�Y�W`}g覉9N@O�2M�*{�(J�8yJ�!�N_\~�҅GΜ�����Ce׀Sg�{�ʵ_���a��kBU�EQ���g{�CZ�U�;������(�D��poh�ZT�$]�8��sg�y�Q&ܯw�j��_�'O��~wggg��\5f���%&e�F��X��K{ۛ_�N�\* 礁��i�啥�'Np�Y��5���碑gW����y�҇W>��f	�+I�*׈MFI�@9��@6Q��/ :y�q�?�a�:�����3'מ~��/`���:x�\�k�+�&���{�? ��?�muyu9�
Z�&����s���LS�Uhc�]G=����r���}�o�%	앗_^�� �A$P�$
�2�u���<�*_s���! ?��ⅵ����#��tK.���;� ��,�Pz����cr�D�ChGa������8� �Ȓ��%Y@�'p ��>����M��^��-M���.�|x������6��l��NI*Q����=hE�rii�'���SF<��Z��?�ȥw>��xlu��:h� ��d���š?�@s�(�aHL�
��۶�|�(*�\Y��Ň��׈hVf�����/��Um{k#+R�*Ҽ�ȧ|𱧟9u~j����[{�[�'��@V�2��(�RID����:� `�=	}F��K �B�����n�s��:x����A���	��Ѕ���S%��^�|�_�l��C!�1�_���?�������..gSӵ�u��h#�@u	�L�:���^ZKˋ�����������0����/����{?�r�F$+�J�$�� �VË��O��C�k� ����{�s} D2'�qZ`$M��t;�a啐��v�����ʴ<�4M��ɀ���N���x"��� �7�u#�HC���9.5�����"�[��;�}�C�t�����oF!8B�GBB� ��uT{��ȼ�xue���;�l
�.����Ǐ������?���5��VUi\$�ФY�{��(�n�o�&^X�7x�tmrw:��8��C���pw:��&��Jm3@([ ���2�ԏ!S�2x%䪼2׹rk���i�z`����4^�D�K���+Ca��f@�0-������g�y���b���cKW�W���3�*MJ�%ic�2����APdeMNŇ9�1p�C-h��_����mYїO���sP�UiZA�9���x4�a]��EqO Ry�]�>%J$娺a@�5\���+���<�NC��Pi��=�y1�2U��������t��$��l�/� �` qK2C�����ӅFl� �$�Ӫ���?�����T��+s�~�*ԉ�q��-�Q #�B Ra���r� 0}Y�5��7oo�a�8�C�ı ���$�(���N�y�`6�!�0�QN�`�B((I䃢�2�:���8�ꂴ�����	QB�UE-�*�#��� $; mM��q�ׁQJ4`�>��omolj�ZQ_�dنZ��9�F�{���������ڰ�'/������y�膅��jL=���E�Ʀ�5�R���0I3|�,��?�_~e}k��~׶�K�O:��v�5;�[��o�/,=�_Zj������IJY*�Dd�4s�}�s�&�_����%��T�C�o���.
��J"�q�a��X)� l�&��m�S��'wn\�L�c�nǆ ��l��7��?��?���S�}�g��B� �`����x����\_����4�LS >]*T�8|������������_x���9�Xj�I��G����W�?u�Hp����m��E,ab���� �A��a�x�4r�&K@貎cC���ω��k�ճ���YrXjȡ��,"��P]1;�����\IC��/^���0/���${�@�^�ܹu��u_��_}��ov�ݏ��6�*��re������9x����0G�tu8��i�뺇++�k7�Y��W���㏚�J�,<� �"�tbu��c��K�6�,�R	hQ���;��a��i$�F>VC6��@��9&Xf�H�����:tRW�u%�f�\ -�^�{�+ZX�B�	M���y��o�;�"��� ��k�?L���+[���ݛ�]}���>�I�:�M&2���j����$��K5�"�dcz�0rue�;l3�hB�D_�p�ˏ=Jexؕ���+E�ܐr0݅�6˚�)����:1�jz�Պb�YqٚӺ�e�����3��0u>�rLtko�������2*��{x�z=��ͭ�=$�o>����5�S86�ZC��I�wN_�z��W�yV���j<ODރ�t;���_F�Rה�-q��on_�q����vG#�.�=�ڟ��d,ZO}׶���0�q��>�zcw� �����yI������>x� u�6��֫MU��Q�������u:�ZcSu�$߂�@\���TD��no�o>r�iX�\�O��)5�cb��s�~�!/�Ͽ����(4?��\���*�����*2���Sk>�����$YB�C�7 �5�l�^[���=�g� z��C<��q�kx:��-��k�"U�D�S1\�&�*�(�]XfiҴ����
���[�4ÐH��Q�ئ�|ZV���*�L���~�3�1*(FPi�dF����s;`2~bnH�6�8����)c)�S͚�2�_I�̀�W060ޚW:ݞ���n����_X\�H~�?�\T���/B�b�+�Kϧ���޾�Q�-"Oa�g
���ȉO�� Ծ"R���8�xrM3�B	p�Ӛ�~�\��H	��Dq��Q���� n��{�y��/�%F�E�.���A�u{]꤀3��z�;��1�g	9�2�C` �p�l�A*�\����,;��2Z��O��P�Q�<+0S
����f2�� cBQ�bC��h�0�i��R�/XY�6���ȸ,��S�Q��QUw�v�`Z1�x��80�
��0>�u��3$�����fS"�+O|��,D�)�HK�|���R���>u'JT��׮W�BL�ng���$����?5�$�1�@I�7�F塶*�y!YC2���Q��~�������G6̲�%��Ys4//.��iх�A�Xgn�}S+<���!#t]w����a-�TD��^�νutOG�`�H7sj?��|���ģ���R��j��S���j`��q�iP��i����Pd:*W���0�T�K�G4�kòiB�j��!a]���zL�)�VT>{��pӀë�ִ?��`8�'�]PK:��@+�:��"��)�^�����n)L��Ҹa|�)$�%?���Ǔ�x�.�Qz5�0M�����̾�ƛ�����LT5��)��"��a�d��<�[�M]���,�Z�I��xl�5���T4yX� �	� ȗT4�q�I��"8h5�<��2�n�WRj�4f!�w�>�H[K,Yi�4��w&S�2���d4�u�[�ɱ���*5d4�L_֕!K6�R�y�@K�s��q�
`�t�n�FHI ���d� _�DI#%��*�Ԣ!���(���㣐F�zp��h"��w�m�z]Ǧ<�0�������}�����$�Q��wQ�U.Q�M5#�hU��@Mx�?S{Чð]�ᣄC�]�νM�w�(]�����H�"6��Y�����(._��P�+<����@x�8�!㴬��J~��1�q��-��&3ݴ�1�n�O��>E�@V��1Pފj�zې&C�<���0�zY麹�;����!� {�k6mw}:�l�y���.�E�{MU^<�F=t��p�Kܹ����~^SGѡ�T�d���z�ݧ������������t{�[?p���*bd�F5aD�B	�ʓ(++��ᒍҦ�������H�p �ג	ô����.PC�tj�o �}8������.�����̤���b��i���[_���RQn���"s>SY�5]Q�(��(04=,� �H&,懧�2�J[�b�p2�P��g�A�;��&����C���ն��tvw�tbEZ��$�$Q��;�@�I�u-d�0D�@+�2�Y��9|��!x)b�1�Q��X�<P�H�Dh(Hb���:6HJ��D7�q-۹��{ݎ����-�������c�Șo����V�]�|�h}�u�e�c��,0��M���Z�6T�����vA��jw0�b�kY���;��폧;�a+780���&�9����^A=I��� �hLhy���~e�I�H�0`[M���'*@;)@P��ڕ`����LO+�$�)�R��ݰ��Š�w�m'��dL���<p[R$����+�ׯ}�����v�XaPhyW�����:&��z�a��a��1-}2���S�$�shj��ɹ~�n�0`�7"���LCsd�'�R7�l�xVP��:�l�Q��d��ꆭfY
2��#r�"GU��@m���PVi��!�H-0�m�"���`�
��� �@�����J-�8ʬ��b����R�o����p�s�]�~��������� DIH��` Pk�Ӧ��Q�IS/R-��	��5w؅胆����v��h%�T�Ѕ4񳬴M���I���[��H
-����~�7��*E� *�8�	�Mr��gD����#��v}���"��z�%Š� -��p_ה���o��w!��F��,J�0����صM��_vaa��K�XFB��N,>"	^��Ȧ�8?���h�9�L͜�]�Ǟ���I�W(�(h��5^RgqQ@!����@��Z]&�Sh۳��ZT ��|7͒1H�E ��$iO��VTqC��%�0L2�%QDW�ڐO��v!��S�L�P��)�ƛ�ݒDnei��ӧ?��V��q�4��ؖZ��ـ4�\��;��	�m&y���a2?{#
%��� S��TI`����e�6�D��D#��|��p�y�݇�������qX��B?��p�*�SjgЅ|�V��򄀅k����ƃn� �P�Y羿�,�{�%E˳=P
����M<8x#p5��"u8qlaa�Po 6�(���َ7��;;+�]*�ᾰ75�4�x�YV/(���@0*m���z^^� ���i�!���	v�[I���1��m�K�Q� �Q_ЈJ������h8#�L�yR�3-�Y4���\�TU�dH 8}�Q�&�=
T��-
Uy_�K��7h�OR��]bv�0��WU)���C8���@&) 0����'�  ����c�W@v��H��Q�#7�"��bd8�*H���t۶:�I,�+$�2LsE7i$UCٽ�2'�	9HS�Z�tM����N�P'�E��TZ��/�k�?5�K�H5&���� ]��㪲�H�^$��&?d@��?��:�>�� ��M�#W^P5\C
2���c�0y��n�� c���nZS�"L��c��x
�&+ PBU�Q�~D�}\�2�6-s}k=�F��N���YJ�a�A�:���#��s=sPqd�c�y
���iI"��M&pE�cK0�p9��bk�Wq�z0�9��`�F���~4Ol��c�7r���/���m�dVU}Ō�<G�iqa�%��7K�4��l�[U��t� ���g�F���L���s�mooH[��⃫W=�7Sj+��뽎Y9\�JU�LF|fy
cW%����I�P�I��HS&)��I;|�8Nj�pԚ.�"^�u�J�$�i�&L*��v�4��pE`{#��a1&�Gw���:��`���,�}�����H+I����nI�S�ҿ���Nw8E�':r71�C*�hRV�������-�c����Z���� �
��֝͂vC;jӵ5�7E\TE>�{�
�
~9��(%"႔�m�u����筮���m�	0�AZGqPӞ�b2ɺ��������3N��Q�$Myd� �(�ADx���FH*���]Y��(�jM���>�����}0� �����$��(ȭ���ئy�'>���tr�ʵ$�tM�ģ  ��EY�(U�@#II�Qt*D�N>P�`2��ty���>��מ<�#��G?��2�Ԍ6 !��@�T/�`|�4�x�h|\�i�9 5�Zǘ��BQ��e��?Ҽ�E�2�#=�&�L12L��ݤ�bˢ������k�;s��ӟxc��襗׷�+:k@�/��5
আO��_�$Nk1�&L�A�ۢ;�2&�DIb`�?{���Ϟ\���?�o�����}�dM�R�4L�cC3A&*��*��i���� lZJ���&�ъkw7P��t��/�<�2��kŇ�UZʉuPBPK��MR�a���q;u����{��?x��yU���_x饫�#m���Rd�	i�8!dU�R��ZlrhÆ�����psF�2r�\KV4�1������מy��.Y��������O~�D��WQ@6Դ�K�/W�v3�y��5kXd���2"��jډͱ� 
�(<ME���4CT ��H�*�ر���9�tm�::�\���TAՄ��n������_��Xi�eI���"#�#�6̘(pRڅ_v;Dw{Z���p�|2ױ|�k\խ$�U�vh
�������aQ{=-�5�m��̣�g���~[�@mx���s�W+i�Tb���*�n*aW�����s������Wj���xcD����]#��w�Y�3�<4�e��%��ͨ�� �h;�$5�]!�5�0��Ai�͠c���d�U�2!0~����8�%��M�� e��"�UÚM�4�j:a#�Dzl�v�aL�����$i0��%��
�t� O���i�����I�A���4P+uy��@����߮�"_EQ(�4H
�9�E��PW�tA�c�%�8`!�aN���C贊�	 E���5��j:4p�a�U��&�" �0K릢
j�>͟�S!7M)U�<��t�[�*RE�k: �,���8���o����K�KEW��I8�m96t����Q������0�q$��|π�hO�,M���tG�q-����.u�5r�v��d%�b &�ZD e�!�3�jd�Vh�� �d����"��mPV��'5O��aL�
4�1��9�B�10� 	�j3�����
G�M�K��hci�
�JS"�
�H�*�4��q��܀
�IB���(�m�k�e�]@ٝѿ�cQ ��,2�f@�@�����I����<:���\VT��?����\�Z:���J�&�0�mg3m�iK`i��^����Y�n�J�3K�Uf`R��1*@9�PY2��<tyy��E�m���i"��qLȃL3��<
W�q�v�G]�D[���h�����;����L|ϣ��8�㗴cF���"��1�o��RQq��2�Ad��&����#�MS��xn���
P�#�vi
�J�:KR��� ��g&ۆCY�Pނ�ʔvrt�(���@0�/-��:�!�6��e�p���6PB�9菢Cv:.~U��wEa M߲ۨ�3�X�w}4N8�9��% oiq���-���I�wMmJ�Y8����6fҽ�	F%1<
�R�B$	�H����b�6�j���ʤ@Sڗ�7�߇W���66�
�F��o�tF`	dP�D��}ZǥMy��:���s�遜b2�IݤD>�6G��tI���kQ�)0;��j?=�(@��*�Y�`f9��e�\A+�u�J\��c�(�<��$=O[�,�KA�����"��f��¼�س�hg�2�N��*'T�Ff��P�0���P/\�2��7E톤.�D��癶�̰����o,|���FG5e�ēt;]:����$�h�%q\��I���r��j��G�#���$��ݠ6c��#f �b��X�|R��� 7((8l��qJ�é	a��Øzm-4�<I�6a��������L�P�M�VS�טּ�6��j�
V%x�H��!W�Ѳ�F\�i�YN\��7叮�ma�-���@��d�lÿ�s _�ԟѨ$vОB��ƥ}�E6??�����U�&	&ɾ��%�n�n��Y�)QU�!7�R�:��ȯ0>xu���l<�3/��M���	�5�Vh�y����3��H5peo�jB�N�1��eQ]Y��4"���X����JO.Z�;�����76d����sо�4
 ��D`��jlo���G�'�(���xh]7��đ�V�9Ͱ�?��ݎ�?�LI�aB���^��L���F�)�-~���F~�yAg�I���3pk۱:p+�#o2֝xEÉ�dJKa�;�V�FZ	m��`�&R'@m�:��'�0�$ W*q�Dd�uq�<�ȩU�𴱂�b�U�@� ǵfA�U���(*�cJ�X͡�����2{�Y���c���O}1�l[�8*x�QS�$�\���$@/E�ɩA�[��)p����æI�-PNہ��tUQ�3� I��'Pa�y�2�=��ʳA��sv�}��D
4Mj���C�A�3{#����7m�8(Pd:g�Զ��ե�Wߠ漢�{�Aʦ�_�)9��K�^�]�itF���;
g3d��-HȔ��Ƴ(���Q�B�0�4O�($�-����J��L'` ~e����yA�J�1����!=q�G
UHu��hm�7�ZG(kQF����
:�AlJ���,
���vv���4��\;\;�Xx�h�A���1�v��a�Ӥ=v�ъ%`��ӂx	���8#�?�X�����!(i��̓!�r��l	������F��"�D���9m!�tz3~&I\%m����؇&�A�<�E���Z]Q��m4ܷ ��
k����Rb(�*���˥�=j��S�D[�VV��O�x��fy:�4�]O�P^�še��(L���hJ=�ee;5��9(LS����8v��[�g��V	rV'��2\Wǘm8ZI['0��r;�WS�nV���ؖE��b(	�,0���t��m�M��!lu�F8��$�i1�/��Ӧ��5�$�:��j��Ͷ�=Q)�3 �M��I�v���.�ݾ�����M�yF��	�,��dR��b���c�ڸ�� 'H�H���w߾sr�ĩ��_^�`;�i�*%P�SZ� ��\���-��t�J�N��Ǐ��c�E@d9��L�tS���:'#��0�u���NP7M��\����EoD|�*����A� �i��U�y�G�_(JBˎ�L���3������b���d<Qڳ�������]Z<���?��x�D�	�P��퍷v�N�1L������{��a�kL�`\��ʏCS���Zqݲ�)>��7#O�oB�S��� �#�7yj�0���-�Y{Z�Bj��0ڮe�%���t
^J� ā@��2�����l�A�k�p:�X֎��{�K�eb(j��no�LF��ť8����Z��vm�Y��,Wl���ۧ�Kmؤ�GÙ�AY��g��<q�O?��/���5Т�g<HQ�����s$pk:I*��z��
c��z_h�0X22r��p�@�U ���D�������]�N ��z$�	�СW�.�=܈����Z��aJ�8�HC�Y�,�o���c'>;�GMg��{������1x�A��4���.|���'O{�ʍ��mǶ��kRy���tsg���5R��^���^}�j{~5�+Ǘ��,�[��'�c�i�48R��B}�&Mf>���N�F�t�D{����{E>�����T_- {ZE{},Ӡ��y��G�V��Vg�zG������XQL)�J������G~���ׇ7nݻ{WSYT�rd���6?�?�ģs���Y4�~��ڐ��I�j�P��ݸ��}`uE�ߺ�����<5�����o߸��7L������[�yۤMHj)4?���Ҫ�a�U�d��(>��gt�F-��+��B�" ϯ�<;�uE�UY)m�_�\�I�6[�j>S5�T��Y{�k�\<j�(Km�߽r}<jT��j�W�[Y]r�n2�i�'O�sP�)XYW����k߼q��'VV.�=s�g����%<��r���-ZL��J|����Q�t�V���J��������Kگ�5�&��݀���ڃ�R:0KP�iO2�� م�O�CU�l���Gnl�l�k-.t�|�ҥ��V��5	|�olnoVy�!�6�-.��\��c�V�d,� �r���n�	C*cB�h�����[�y�����y�q��$��K>��ཌྷ�������!-
��XvqE���?���{����I�Q�7��q�����,@J��Ü
#��US�O�鈌��!̦f��=C���7:��<���Pfwqaaan�q��{~>�[�|�����W-{g�	��I����ז��gc�1���O������@1��h� Lƣ��[���7�yV9bc������3gΝ9Mͪ�t i{��A+��Vď��S���I�`�m��-߮��.��߈r���ݽ�zA����@�[4��~́�~��򫛛�SQ��Y�����ib���s��{�G�!�9���;�w��G�	�TTI9�?�z�i���׾�9������Ф��h���O����_�d{}H�i�U��+3��.�Sk�=#}t �}caJN��8y|yI�M�8��3�&�������]]��7�y��_�B���?z������A$��RZs���$Z��>��W�;j��I?��{to�`WI�j�[��:�?�z��r��/^���.;_��_�QU}!TV���x�:#�e�eZy�AE��h6~����_`��L��-,.�?w���{S�w:�Hy�5� �*+�^������K.���Oe)��y�r����|��w������P^��T� �����_���n�g�|�Xt���3gF��_��%�h2�t_����p�Eɺ��i>�yO^��s�̏��WVV�߿��+��l�[�BK\E�Q��hZG�η�̙�z�ǍEFG�}�K��lo���͆�Mt�8��#Ww{�a\�5���6w�|�������.�7�5�����[�/_~����M����mFq� 2dx�v��!����W��StV�'�C�U�����$_�z��D�������	����ݭ���[�gϜz����V]���=]��uiӄIr����^�u{���-)�G��c�n��N��qh�r=J�~���u���h8�X �'8I�o )�]~7�s��:�}� ���Qjq�Ɲ�8x��w֎/=p|yuuia0pM�6�[����hG,mKn���]��v�mY9�u�.H�ͯ�����UP<Z�*+�����6״}>~��&��;�����.�PT��@k`�b1�����$U�,��W��?��n��v�e�8w��"��+�,k���P����f�`�tlU�����[
�� ,���:ԍ�~)H�@���nC�\bF!M��64�$�y��N��2��y�Ck��ƥ<O�DH?��,栙��Ɍج��~@Uj���Ђ��Ry����hOz�]HSY3�9�У�S�E�v�D��$��=����?���_���k��ϞViAN|��M(F�2���ЁK����:f�Yx��vsf7C˲�i���[:���Y۳�J2
UJg�A����h�����4N=u�6\o0?��!��H�f��5�Vm%S�=�������E��Ty�ѷ4P���xq.Ȭ�mY�����4+$I�Ø�M�Q������oZ�QG`}��ZX[������'/O'c���l*���J���&�Ш�f)E�]�i'��aB�
�2 &2-��WS���`�rZ��#��m�����*�f����,��tC��e��Yե��tP*�r�w��!���B�ʲ@��S�˃�n)��Sf��uV4ԛ����x�)D(���_��;��J�n�ş�lo�G�P{�J�8�et�Gg\�$��Ң�uI��E�a��,���Q��N�6<\)KK jܞ�#��t Z+����-t\��aU����E0IY�
׶�i��7��B0�$E-��{�ڼM_E?�
:sZ��vu�V�����j	a 3~~`�:���oc��)�\_��4M���O_]|��^{��;�{U�u\7�S;�b�1�:�OV�)&�0t�T�t[�3���E��v��iD�;�j��nXy�^@�óB:ɋZ�lK��O��q=O�(�桮�S55�
C;(����Я�,5��K�g�"���Q58ϒ^�M}gk;���y둇N?����_ �5�>���X�P�W�-..>|��[���;W6w�����!/�+E��Zi��-�R�$2W&a\+�c�kkǪ��fA]5@M��,5l���-�>	�+�2+�1,�*k��
I�g�e�����n�H�~��$j�c�H���ϧ�s�<�u]���J��ХsgW��O<�ؙ���_�_L�|Acݿ� J˫'����î\���k7�G>�}6����I[=�^Tu0�
M-�u�F�������e�QSX�5�s�,��2�D�x���Tn�1�,��(�ﯪ�Z�:�b��\Q��sE��&Jՙ�(�π�g	�����./-?~������+���|Q���|s&2���2�}��g���h<����~g}��� tdtY�� n��`���9xTTY*K0��V������z1�L�穝�6]+YJ��<�~���(�"��h�m�o�kӶBY���vS�B]gԛ���BS$d�ť���\��Ud��-���kF��9<��sKZ�N�`hgDC��UQ�}�g����e}j��i��G��Ay:��?�%~P�;`�T�k[@���(��(�������=��ZޮW�9GP���Yˍ�Ƥ����jG���    IEND�B`�PK
     uK\c0��T� T� /   images/2b856d38-88e4-4759-8ee8-6b01c1d6fb9d.png�PNG

   IHDR  5  8   ��e�   	pHYs     ��  ��IDATx���$7v'��83���*6E��>$���#ٮ��E��?0����خZ-���:Xwޑq��; 8�#"�Ud��ϊ�w8����!��R)���RE
��RkG������#QB
����:<�+���q�2FI%L�?���4Q$�2#�ئ�ߌ�H��Z��H��f��sOK)�����.N_��NlJXR�ot"�X�$5,��R�[�ͻx�&:/���R�(
XU�����?M�C!"S"��E�A8������5�B�\~�T�_�e�I�i��X�8>y�f����T�l�Qe�\.5��0�ME���yZ���7��{J^%�*�$��<�?�}�Ϻݮ)�צ��������pE�<ϓ$�#BgYvyz��ŋ4�g�YQ.����	��Y��K'pv��#�1F{����] �j��'���}Dd���0��(�u��_����*6�~v�R��4v�GYd�>C�Kͷ+}W����0A� 	�	���B`���J�|ʂ��Z���c)���7閴�UY'���W^5�'�g���2�$Z�~��Xe���;�#ฆd"����RKk���b��L&"�a�W��3�t0����wL���� �tmE0�#h����RK�[��	0��^@��%S�^X5R��L��o����K� s
��B�>T �qm�8�|6�^� �-�e Ɗ��D���Y�F �H�Wr���i��hi g�Ӌ;]�Z8i4vI�����&Zi��,���U�w^c����ۄC��W�\'�KҺ	^@^iqz�J�r7�Di*Q�\
�;[j)$�Q��
�W����M���H�@OC���)JS���B�p<j܍�S <��J&��jR*K!���
-}߈g{Q�0{K#`�����>�}6�2�{�EZB6A�t��w�+n�e0���W/^@�.//�g��2N"3�d����Gi�}���{�C.�i#5���磑�$]��4R3�U���l����WDkO� �)\�4��E+���&��W�����3!�Lr③Bl�t��8��|6�#�ζ�5�t5Y%.�&�o��,�K�ٮp�x�u�C8Ѣ�R� ��U�p ����J�-}��o���NNOf��dV1����v���f��Ud&�.��X��¬���hݴ� �����5�ű��v}Ԅ)���ă���?�Q���H+#:I�|�O���x{��^���t�)�v�l9OK�'��-8��2c݄&k�!}C)�q��D��Pq�˔���X�3�g)��1K+�bqyy�;؅�R�z"%�h��H�J �S�.�2ڊ�[��Γ�SClp����;��j��8����`��	ŵ����τ�4�I�6���U�� (Eg�&{H$pݠ�I�X�@�\8!�
!��[0C�&��.j�?.&������m���/����w����K�~�Nf�?+D�3�5֫�6�3Jol���ɲl:�j=�_�ݮt��Vq�����T?�����0{+\�	g�u�I�jd�2<��#�ߙ#X��K@�Q���cڻ��5��-���J�4���i/?���z��U;��ț�NŊ-���Z��C0��(`�2�L&���/��a��F1[�d<l��J�Pɚ�L�����wb6ދ�_+�"o�u��������h��:�(PŽѢ�+ŬiC�n����H?�
�މ-� WEq��]�e�"3��L��V�����h�!�%�R���ϲ�Hg-�E�)̪�(�3m�|<�D7Uc"�����ba�Oc�����l:��:��c�U��#�M�%�7�M��"e�a���9�Z&�敾����vCo��H���,].�G�^H���d��1H�FYZpf4l�sT(�Ŕ�CVk~s<A�5���O��(�܈��"�裏vvv���B��b%}�o��J-I-�dx'�b>>[,���"�*G�]Ԣ���Zj�;��f?3"k�q?	J�3��$u-I��������힬c�9e+X�$g�Ҵk���Z�� S�4xN�F� ��O�GW��sƴ�EBj�I�[��RK�k��
!��ryzz:�x'�.��	aB噷���	�BF��s�D}=�]�q�ӝOѩ��t�t��\�%���r� �p_`}��I�/��� �N����pk�A������i'��n��x���U���mR}���1F���'��`g�Ȥ���eD2M�Q�h�<���ƞ�kk�[�����z�$����7�= ji������iY$�AN�5��E^�D�*%[;{C���A7�>V��Sw���'�rA^��T�p�H���R`�Kr�$�^>�~��wE����_ȀY������峧��A^,a��͈1O�$��P��À�F%q'�)b��H�V��6v�#����?���5����@�������}Rci U�g*����.���3C���퓱�Wl��܊S��A�6�M���Ë���w�pV=�U�'т���/�e��E��ҏ9Y}�J�&���Nc��F��[����l����7�c��1��mҨ]�`K-}'�\�j��x?�ϦZl�ٯʎn«���<�c�m���1���쁳�	'���̩�l^�޴c"&J(����!#�6_�A�z����2[Lg��.0�8����#�/�h���8��Z�d-�r�̗���
s�I���Z���r����~
��&lⳈ��R�7��&Z�Q�����;#׍�6�=��=|��?��\�'�	�`!���ZX�[Zj��'/]�sUEh��^^L��*y�'I���@�`�d���A�F�M���0A%����teچDQ�Y����̹"�g^�W3|��@�n�fرf2��(ܸq�֨�q���˗Yav��V�,A�����B�Y�e��!*��֜/��z�ゃ�Kx�m(Ϥ��k�m-��i���p.�xh�7��Jx�*���w�k�Zj�)L<i�|��|6���b?���R}����}�֒�N���K�Ÿr�李h�#�A�G����1���Z�!�k��K��v�*
̋�՚�
`Lwpk�\9�F;�N�����l<�w��^�����=-�����kN�O�]r6���.����B��~Г��FD�ҏZjXb�n㎵9-���!�䔶�&G��bC�:MX����N�P�p�;��CA��¹Hk'~؁������\�%�u�,{��Y��PV꘼'1�$ղ$
DJ�<'m���#l�ۛ����!M����T#�3����]�<�isYgV��X���L�UްA$:�`��t
�,I��h�5������Ǐ?��Gl ��m�wK���F��2_�/z�����%��[���!3Ƭ��������[�*�����b���jn�j�V}m��7D�)�bJ�"MS��E^?�/��XRY��F��k��b��p�!V	�k��)�Ќ ����l?�m49�8n"�|���L�&�e%2�eV��#�.
����W�����ph#&L��h�CK�2m�EW�N'�t�����|W�ۆZԗ��J7�j�W��բ�T��-�%�	�0����|��9�[^1�V�k�!�/�$=S���u�mZj�OM5��G(�7�@f3JF7s�r!l��}����Re�\�W�իΠ�?/����A�xQ�l�7�P��D�(,g����n!���pd(��b�����燇�{{{�~��WK���*�cIRf�e&Q_�b��]]Y��q��~��a�ي%=C1�����Ph�B��}&�ҷFu�3�`c>����moo_^NA��&A�������gv)d
�:��r`>q�ߙ\Lʬ��$˲$�ԴRy����9�#P���Ez����w&�@G�Tt��yA�q��F�
b0�i���<|�����W����`P���
@պ�?~���қ��j����1���ك'+u)�.0߲��@�����d���|'|��V�r�-Qwm`ŕ�6:�ձXL;�8J����C%���W�V�����\�͂!X	�
4b�X��R�X�H��V��,����sI
j��/�KX�ƮJ��F�)u��f� n��A��]����u�����WuxQp�Z�����4��6в�^`��?�%_7���X���ϻi"l4d��V�z�8���(w�D/�^�<O�*�J�y�=΅�8�v�����
���C�蝆�ð�g2�ue��V�T�<N&���ϓQbY��Rk�F��F&�L�X�3���aEI�%��gX\2�<L��+ho����u賥S�A�3����[���g�}�����[TcA��H��6Z�^�u��qP\E�m�ҵ���hm��@))U��[�_�4�Cnd%���`���>���R8=�Gʋ���H+4{%����7�3ZPd���4mk�al���A�_�y�^k�!�r��Gn^m�Y{׵��J[] 7�(f|������`:GGǣ���[i�Ӂ�a)�T�MK��N`~�|�6��8��5S��ҵI��e: �p?o�, �5�����TXP�1%
\�U�.u���^�EWj�ָ�eB��;��M�5.�{�ƒ�����՜����VW��?7���k�,��.b�^�M|�w��7�g��F
*>~u�n��8LSU�0ӥ�
c�1*R� �Q��X��%�����0D@�z��%�'h��>U��E^"kນ�ן5�q
�3���N�a|s������/^�y���W���7[��ɯ�:�9	�?WC�g-�����g'~�z5ޓ��7R҆[�Z�'�+�à�e��u�����`��9,�$r*��pሺ����冨|�5���q!����z[�y̽�e��2.�Zh�_�L�4׉b>'H���φ�������ыagg�JS���Z��i��@�ʔ�O��g�a�:4KluSQK-�>��,R��1�ZmY8WM��e�3d��ضPb�@JU�kFy��7��ߔ?�W���['�Jb_Ý�H�Z x�IWi����m�?��˯+ܳQ�vu���[�.m���Vs29�CWH-��&o�$�ZX�ł3�by��_l���*��ni�I�D*T�l�k�X, �I��b�l�º��֫��V^�V}u�
���f[[[���'O���h4-��� ϓ�5���y��y�uK-y2���y�m�r���̆�7q�+f��M�n����x�h� ��W�F5�NO� W�"_���x��b)��4�����ٓ����_!�3�Ÿ>�1����<O�����?k���o&�W�A=�?�<D��rI5��|>��8��n}�'B�y����<>ӡ#
���l/�������rc�Z�����u)І�HyF�ɹV�*��E����]M�?���&j�����?�z��	U�Wk�VF �-��4�@��>pը�e��1��(7�P�9V}\�}�-b��u^ȕ��5yt��w�GY3n�7k����r:��.fc%�8J��d<�`ڳ"7�ĕ�+]KtQ�O��)�x�4�:,�s�3�����z�I����
ά�Ne�s�{'��9�W.���q'ĵ�Z�WjB�.;Ep4y�%I�QFQ��;>>>88�������kZ�4��Bx�I���EK-]�jR;M�F���p���O��AoDK-}�Ė��d2�K]`���0�|>' �5�J�K"C}�p>ǜYI��*�+�B+VD��	�B@���1�]Pus�h�l����+�6��Y�EU�A:��tJa�DB�����7��~)�<�;Є�44-�j�[$Ju�s8�2�[@�Ȋү"t�i�'�rZ2���x}V���jJe��hQ�1u~���%Zj�RS�a�^c����|cD���m���QT(��ֽ�d�}��ϸ�|<����0[�0�bN%���:r�Z��%l<�e���'�c��@�a���59�T���X�Qn|�j���WDo���h��ʲd�/�X+2G�t(>�E�+ۅ��Em?�\p�F��-�\��H��+��N�e��zUY��W,6+/�ƿ,<J�.���|�����8;D�$���œ�_�:�Ӓ(Ɯ��L.'���&�tb��S"� 3��9Nv
&�[[��=���އt���W�AS�ZW���g��� �aS(���cc���Ъ��x��:l�U�zܣ�W�����2/۠���e2���&���r������U3"X�Ѕ6r��M$i+gg�"���{�77��]�woa+�X;��B�URu��Y���M�G�gW��Sa��lBP�F���6Y�k�5j5�lķc��᭚C���LP<�)J� PA��b�Ai��S���4�hu��O��c���J)��"��Aƺ�eP���m��@�Ĉ�(>�2�}y���d����'�O�r�c�)l�q��f��b9�[�1�������B .n��4��5u��V_8h���~���ڤǻN��]Ó�����m�L7�Nb�fL�@k���z������!�|�ݬq�i����"� �G���sŤ�*	J���\U�j)���T^��N�-��ջ���XCυ���a#�ưgqs��ěL,�"	���.�+&ײT��#C!��y�DՎU�l��j������wm�He���
��0H;J����i��B�*A4� Z5nkG̺*����	QR-\Ǒ�U/��h�⇌�cRy#<'V��#4 ��{҂K�(�%�ޔ��=\�x��s]�f����:��R1�5��m'��k<�|^Z7�z�q��O��N��	�ѳ�����@� ?O�S�g�r����'�+� ;y�Y���9ø2/4��$�K���t:��ȣ4�opA�5�H���62�lO8��b^��gv�<>�~c�_�BT�`9���ϡ�ֈ=�`4<x���F�9��!���$[��ҟ��t�u���53���^��;�M�8�"e�(����Ҧ��� ��
vnk���4vu�M(��6��La�W���A	R��%�Lp�l�!���� C��|��Z��r�MWKlE�jd�G��R�>�:�U~)1�!N�S�C��^I8�:C��v)���T��}n$�"�Z�'x|��Z~T�$��V��<N�;j�|&���}���}���	�͸�d�TX�$���:ZV�q�0N�O�{��1�g������	ͱ���?���6���N��uV�Z���q�5�KVZ�&�x�+�#n�����F�'�9妧�ǝ�����{NK�U���Y��S~m�z��K�XQ_��Gls��-�xi��O��%FL�dl�?�b��5�І�1�,�%�k/q�[;�T��z�������,�sK�}s��i�)�����LHE}�5LqQ�.�����a�!1x�@�A-J��Ͼ0C�����cb���s��Im��oېN�gH��zp�1cW-U�)Q�t�.��T��X+��ҫ�W����\��Wx�=øM,�C/�ʁ����2/��|�.��Ϗߋ�����C��J���4a9)���N��[�v�~Yb%u���R0>�.�Ɣ6=8�<tw&ϳ(�����`M�yF�Q7�x�ݯ�	o{������A�Qܐ�s��ԸĄ>�� �?⧚}�u;��x<N��[�o�K��g�&������t��Td,~}#T��V��@��J��`r-��d�3儖��^�����yO�?����U#"��hrUVXE�T�
����"
f�q��OQ�/�Ց��n	a!����|��A��ϲl��,Y�����˓�
�?���Ux�X҅����U"�`cc��5�0�G��;?��3ɢ�u9x4��p��1�ߑ�FP��[9q�Te�e�`E���+��g�7�{��k}�oIFe��x# �t/��2�y"��e�ҼƋ�|;��e����.�%�,����@��n����;�3���PΩ�4�W~���]]���k~�`ъ�U�4*跶Y��BI��d�v�0j�����7�~Ϧ���P;?6�4n�����<&Q��'��8vB_��F�?��ɇ&�j���h���D�!#y[��^C�ϥ��5�#���Fbk��%9񤍈�Q�g>�����/*�W���,@�xd�\,�gEL$�o�*+�w%"kAŚ$��Z�e&�h�"�V��t��5%��J%�80�**��q� \�Q)R���7R �K;�.���0��hޞ���Z%�;Ն��D �Bj2T��%C�N�5MSzl��љ��˰O?�x�ҿo��n��,��V����@���Fo	R�U�`4c5F�SQ����!3��g����I�� �:tIfS[�L> �P2��Jt�f��&Dd�Z}�W=�M�+����C�'*+c��+_�� �(�U��BYʿW��),��lq||���^�Bk��o�x~FQ�={
S�o(�J��8&�(�OKԆ����XU��,���4���J����~]��p�[N�ـ'(��_��	"63���\x�F��[P��aT0�&]�Q�<AE���_h2�.וP��syy��`N~�lp\�Y0bU�s#�Ym��{���1%���5��{ªgHd�!b�����tS智��"зa�pqv.� }�p��"9�i:��f!gB�jH��w����y�=��N����ܰZ=��g�l��������g����SCFW�YzHE�N%=�(9�W��J��;e�z�v��W��[�B���pj �(��������`��h���Ǩ3���qG2V��.p���HU.,�QN�`mg������?>y� /�������(T��Ddܪ�</-�l���J���,m��Ɓ��lB��O�A����f���q�An��ܭf-�U�3��L�����])N·�C�W���)/a		�"vEX.�N'
�Ǣ&ln��PM��+�t�B�p�k��f��&�>A(t�)ɭ7MS��;�#׎/�\c�3�I#	�@Fb�d��e�?�x�h�D����v�R�"�w^{:�?���um:�S�NrL|��"�$-m�t�JB��T��c�5Y����;j�c�{1�bRfY�zE��;JKŶ���1ʆ��ib��Gv��P_��t��b�
'�Y�Jm9Y<]vL���" X���d���W\��ie��$IX�5]�)Ԯ��XJ��[{`�dӘ�� "!X�ż,t������<�L�V��l<�0ܸq��z�����v1C�- ��ɣ�(�$���]��e��8��d
���}��Q�.JlM� ﺝ��^���F]�Se��t{���,py�����F[��Hf��No1[�c"LTq�Ħ4��Ҁ8���tK)!�l��|Zȴ酢����4�D�G��	����wV?�~���{9ƨdbN��u�Rh�XQ��<Bk,�Sl�ls���<�x����N����蓏��y�sU:1��Hj�U��L��ə&?B����^��aąC���p3��T�N|�+�@	�5i[���ޯU��"'���k�g�Q�����X��\���q�e���������Z�3��c@������SHRb�f3!#X?�J�=yr��]��:�N�vj��$�8�����6�ۆ�0��$j�՘:�P�ʠ�]*Q�#.҄��U$#�|G�-�*s��*�65ASY�A����!��	�O�=�� ��<q�A�Z�������6�j��%܇L!������`�=���U���ͽ�=|�����ib���"�ƵU��O�A�̋��r�����,WGr���G��>���6�5�gK?���m�<��Gn�,d�����ĐWh�z,ŕq�OH3�!up����z�&��tN9Ea��f�BFd�99����c��3��Z���}ˉ�ZΌ� $�s�{^dp#� �L�#459����5��'�Oiځ}�|�"I�C����+���f���5'��n�u��2��$���� xp5w��0C[ȇ4>˗gj��~`���v��B��$��
:��ui�_"��-�*<�P�܎�ΕU���5@B�q��s��ɬR�7����#%	��s9�y�a�++`u]�4�>ѫ��g[�S���\|~S����8�1Сc�����!�f
X�l!��?����X��7n��B��]Kޅ«ǼU1Q [��	&���s��b0鮍���|���o��W٬��W؝Ҧ�1���$��4�Z�Dc��Z���V�1"x"%k:�P]Q
l�nlo�p�^Ҙw\R�/JJGnI�嚟V�^i��t�5� ����~�um&��2և��F�1"MPq&LF�!9&c�
���*��6,�λV%f�����R����F��:^���3�A��3|��]�9�}��9�j�Z2͙o�Ar͖N��'���� �(	x�jC������s=�W4���U�����R��t"�<�GQZ�YQ't�]��9�$�2�ʋ��hv�&�Ż;�L$�� i���%�eN���&.�*3���6/.����t��E�whGk
O7�޽{w{��j|y	 ����u|��7AY�#��ڕQ�9=�'����Q�����0Nwv��Ds���M�:79��̊$�3jD���1��Z�Rc�A)H))x���}Bot�稐Y�#��T� ̣E���l��cjy���-�B~M�*?%9
a�"���vu��Oz���&)��*4�kQ����~⌔U���(d��Å�hu�
,���ƪ1uD�|:Yk<�~�o�y� 83n��MwZ3�+S��d�%{���Z�0P��1P#y��������������t{�"G�vzb]�����W^�����\����I�P��u�5�3��aYb7���,2r�c���Rq�ڜ�6c��y!���Fç�Y�����U�J-c}�۰���+U� c�w&t�ܤ������w�
�1����|;��!���E��]����u�.�~!Z��U�?p���"��bY_���h�������D�r��]��E�u��0�?H\3h�9���?�����v��C������VM`y���_�~�gNIv@��ǣ0g:�����X_Η������l����v;�www�UJ�E�2���09^������e� �qe���K��)�y99��z�ap&kڠ�~�� Ց����������+�g��_8	Z�h����G�Q��ynl�blr=�m���{�`nq���ngx���$e܀�Mbc� 4��l�%k/���V�N8�lz�K���d'-�}�_�0�YR�14ޯ�j��'c��o~��M-v�}��՛u$��9�����
W��l��

�,]܉r���v�}k���L���%fl"��
o��ԟ�2�Mw]{������g�;Qz�(hd���)�`0d��,&0M��bq���²���>_d�ɨ�;�EXYfY��}Ϭ�u��TD�Sl��KR��j���G��,���4�T�N��iLVy�����?xj�h����.D�`���K^��j�c�2��N��(�9�}�A[g�ÚM�z^~�W/8�`әLƚ�.����Cvz�X>(��{�W��+jN6��g�w�E�U�p����yu=�p+��s�j���I�3mE[N��� ���7�ݍ���v!����{(��/f$$����]��h�Ê�t��#�ތ֮�Κ@�9b��iEK-m 㲍��D���ˆj6r��V.�fO����q8���2;DpC6?�n��%����$���Y�� �tU�N'!�B�G_>K��;��~��p8�s_�z�q����/is��`Y	��D�Q`�3*�r�`�G`E�^�����O���.1��U�l��4Mи9���rqqF��?��1 �I��k6�c���� �dV�����Ҕh8�����?O�[����~vpppzr!�lv�if�'�@W�D��Ng+�®;��2�ν3nq'�_���7�}q�.s�|��U"˰
���q����p�L!:Pd�l�t`�`?ؔ�V4�)���i�t���HKB�א�Y�U�q[E����?�ϨQ��ѹ�~�?Z����_�+5�?�Z�,8�;~�🫻������*�7n�&;I�ߔ��� ㅡ;��^�S5�zmY�g,а��� �9�@��>�#<.�r��� R��<89�yx������H�.V@+=e>�8�p_��c�)�)�7TK �bM���۪|�aK���'�� xm�l�5v�>i�X�Yr!���4����S��v���?|�ȊAʕS�e/3r��w�t1X�,�nXSt�������3D��z|���i�k�F�L�dK�[�D��ٿ�l���z$�_9�hӔ�y�l�hW
�y��C�s�x��F��S��u�����}J��2b�B9G+�y_��t��>��^�>ヾ�+���Z��Kx�Ц�]��x�=��{���5O,��$������l�w�(*ȓ��?a��;���;��'�9��K�r�b�W=)g	"੼�1����6�!�����X���;`��}�k��"��(�����(
]�~�j6A�����x
>�D���zl�c��Ͼx��_�9�}6�p-`{�qA`?�"����v�p����i��p��M��i,B/u������#�F8�2#�A,Z��o9܅���o�$�,9~S��%Sᡐ�Q�o�!D��!�p�5�m��ոv��6nᯒuMd����h���go�rsI"
_���]�!��9�քa�W���8��B�� P�3���˱z�@̄e�c�p�������_|��?�.mS�0hP.]7.G�s����\����/CV ��c7棁��y"����0J�;��T��#XT ads�zl���=d�kr���~�ĎHh͗�A�@��8v�T��D����mLe���b��V�"5�
p6�w/A��3p���w��y8ih[�
%����G*�y�@f�9��e�vz����cg�v�UDJ���R+�!����� ��X�ȳ�#IL�[O/�	Nܶ۴��rA{�5��R+N���Q���5��zDJTF-8�f�D^ ���^�Si\��7f�-�H�T���W��>kT�X�Um��I�Kci�����0�!����MBQ�v��(��"�X\��w����x���w~��_��Q�a��\�E�ӝM�4����1,O�'@X���P�-���ј�t�ggg��`����zu9�)��C��$��N,Y*��~�t� <I�������	�q"�
uCBQ�wi`!YQ�8�E���-;����"�����1�|~���O���ӿ��9���κ������_������>:��(F�8��i�QZ��@%:J�(���H�C���J}�a���F�^ ;F<�R�E�k�u����([;x�n�ѻ&߲�n	s���}B �ї���z����b�E\nn2g��V�MبI, @��W��j�ы*p2��P%�z2�+�B�$���WK�e�`��ܨ�pưB�vTM�"��<��ᳫY�1k��kN�k�(�Ao`
�����G8����m��f�9�u����F[��?~ǝ;wp)��
i�i�l_�B%��m~�R����.�J���	YóӚ�T��h���\(�@�A�s�PH�D,�j0�O�qƗ
�3��$۾˼�6�z�,$��؜�/?  O$7�9�-�S�@y��.?>|fAMQ�XI�s*[����W����C��Xu�q��A΢�̿�u�����5��������;]�~��:a/�YD>�9�Ō(�s��� �%�b�&�z��	/ב7W�&l,�h��+��rr�:Q�)h��|Û�����&p� �ĸ�V���!ذ;�[w����S�p|뭷x�+�d���������J���׬��i{�|#ԁI�f�W�^-Qq�a�U���^wȗ�����3��f�r����&�8)��I���%ɰ�{c��87�4��aiJ��!ʗ/_�կ~��
)MԐ�:==��m��ŋp��h�2�����r&��S��E�Ѿ�l.�bR[ⳗ���eT����gT�p�{��6+���ù�WU�ae?t-�f����x���j�p�е �S�ld�s�|��Aa����T7�О��Y� D���M#\��~,�X��Z��}��ڪ*�U�0Xu���c[Mӄ/Ԥ����|6�O^8�%�Pd���4c./N�n-��O���C2��f4�����VQY�NF��{�[���[^�e����҄�'���..|������E5�b��4z�Ϥ��W�Ў�\�%g�v~f�zO���|Ԃ�!Z�@�̍��L�;�v\%������Fq�\f來8OE X�o�M�NtoNV�Y��r�7pU5e��0��-.+� �CFP#���o��җ���Ԇ\� -��_���Ǯ��2GA#�+�$Ei*ta�eץ)��N�����@~�R؋��E1qA΅k;۴�`�k0E��G���j��y����7��ٴ^h-�)e��8��x|�g�~�"���0�@�6X?'_C���%'PEo��Ɨ$#�П�#���@� �m�TRq!����ſ��,�������7@?~u����S\L/F�Q����1d�À9\������ӧ ���흟��..T�:Sq���BG����$�r��_�B� �,�v�ݼy �0@<���������۷���++�[G'ǥ�ż�l9_꥞Χq��7_f�^���"������t�%�#WK��5�N'���[[�������l ����G���dF4�){x	gi��5��K���� X֓'O�8F�)�/w0G���l����g�N�+�9���}"�?�&�v�b{�F���
a����ЀbQ	������1��D2�W>��܀�pS���X��$p6ƞ�e����j��i O��A��ӆ�ElI+�b(ok�キ%�� js��8}�cCGqrZ��0�/�,�YM��RQ��H;C{�Y>'��@�hhm�T�Mz�8�^�V#^G�Jǲ��+��_66�������)s,�?�#_�+�W��T��K){9C7�*�i$Iw�z�v$�>ޔ���@�S��#�ޤrY쒵T|yQ�߲ү�em��wS�g��=�*e�Qpr�a�'>��QX��M)�)55oվ+6>l�M����5����@�>r�N�,�9�M~�{�J�z���\���y}b8�Ď��9�x��,�M�x�����A�ZjiI!.�^�]B�M�o>3˪�!��k�XDt?�%!��1�EG��� �6��_�
EK@�����c�?�����lgg'�d0ﴡ� �ͩ ��D �P��pd��T.���I1_���.�����#�-@6p;�B�ӟ����?����K���-��!s����ǰۮ��gƉp����GGG�c�+9S��;��a����*�G������ZFIr���ˋS
}�a�\������;w�@?�^����ͥ�[,r�e�~#�v �r0����`�Y�g�Y�Xp-� �z9� ����x"؏Qa)ЦAu���K8����x�SeY�D�����Q�<�nxK}[����ҁ� {������]���|���* ����
7jQ_T���6>{B��0OMV��7�3�N�g��K|���wa�*�6a�wh���o�I�뽤�]N��?�j$�s[M0Q9��G0.��pU�<��k��&#��:3���h��8⣧(�m���P�M����]B��k%׍s�f�+%�Q�2����3���`A�N����U��l��Etנئy쒟y��5s��΍�	@/��T�3�S���9MoI.!�si��� OB���J~��E
�G���$�U|ڴ�}'�B.�RK!qvr?�B���ٙ�Q��<c��)�,K'�P�EM�j%)�칸�"�ɳޠ�s�/�x\����G���2,�����#t�xV�UQ�)?�˗/w�v#�@{��0��r:Drqq�a�ݿ̭=�drriR3P*Q�)3���d�yz6�xp��r6��_���_�9���?���k������-3' ��z4��BQ4+&JT,�bJ%�����b����:]�,c�0��l>���k�"�b�6����E>_.{��4�\��:<؁�O�^�� ���O&����Uw���g��;NEX�x�jWx8�f���ra�` �~�_<y��	���ӧ�{;��s�6����1��{cPkbJ�pr�����0yQ�������>�C���b���r�J[�.42d�&6L���b���F�'�`�K@�����R�������Ԏh�P2�>����b����^�q�ܫ��#+x>�ʞ�۽B%�fѮSDU�o���>0,��3<U�C���(\{�U��5KX�B�a:Pb�5AU��s�~��E�?Q�犺��pͩ�z.Ml���#w҇�
�'����6�ǫ7� ����֐QV�t��7��3�P�+[K'k/BgI�M���4�b���B�H�禐����8_�r���j<Wx|ݸ��RE,�J_�P*�9���	h��}�}��풶3m%ƭ�	�^�*49¦�?� �p�����(:;;{��;����f������dgg��b9��er�<�͠ر�w0E}b%�,����
�����Y�)	���	Zߨ���Ǐ��p �������:Oq��G��\�m>e=��?�g�{�n�
B�v�K�s.T�x������R������]�E[�g������=�	��UTǑ��}�B���0B� H�w8������� �ߺ{���ZxY0\���1&���eh�t#��^nmm���uII}�oܸ���4O����řg�~.���tcf����Ǝ~UQ��gr؎\�?b�X�Lׇ5:�յ�z�_mYz+��*���,q_�6��O���P��`b3��ǥ�Υ�f�*�7T��ܠ�Q�fA0'���=
F�1�j�si�m�F�)�q��fq̙f%9�w:=J@�4�!Jh1�	�K&��|�խ4�U�ܫ��N�5#`�ge<����#� $�B
-�B��O*E��RQDJcRj�Uc˯Ս������d���q�U�kV���Ɋ��0����h���0"���� t֥IY�(�s㥓dh��kO�#7�ȷ��>�8����eؿ둻�F�fcG0W
j-��)dT��X����.c�O�1�{5P�8�t>,�z�PɄ�$���"����ىJ;�����;����v�c��K��A(�e-�.���^�{y1fXN��K���i�����D��� �k��f��T�)�M"P
�Ĉ*E
*9M^�֧``���tv����>�I����V�6������x'	g��/�r>[ w����S�y��P���?��?`(��!<<V�1���0��lGrowy��i�b_&*C���a���V���LtQ�Ɠ��㴓ܻ�Γ/ c�}������	'�g�'X�TP\-�g��.�ǜ��FΥ����x����..O��FYa����~���N �>}���� ޺u��t|���c@�Ϟ?�1���̸�}�����֠��}�d0�N�Q2��p#�\f&J�������3��<+_���W̹g���\���c	S�2��C ��j 1�y��dCҐ.[����	V�8�Uy�ݚ5����K��l�[����77���y�_�MC�����Z0�.jծ����:nn���
e�L�Jc�~����Y�v1v:B' X~]�>L5����^�<>�K���sҐ�%I �?�����4*��i�T�evF���x@�M�X�+x���^_��ϔ�*(�� ��r؇�v�3�W���mmִ\�f�Dp�D3U'���W��:/�G^{����e4��"[j�I:���~1�'�?���w+��OZ��]��&�'椑�U.���J����݃&z�~^dI�|��'������^�����ŋ�b���+(����a׀��1&�?88���\���<�3��Hɕ�+��'�'��O�'�G����ɓ��{ ����I
'\���0����Yu A�i��o~��?�/RTS��e�v�������Jg��Ϙ4����dp/,�@��D,E �m�Q)�!c�/����+�.�bG>�{�p�͛7a����E ����O�={Ǝ}�c���	O�M.�'���/��/[�Ìr��z��l>78��5s�TO�;)�}����Vor�J8Q< ��5��8� ��w�C��Y�������M���v��v��z& �Jy���&�Q�=��Ӹ�z�3��%x�hh$
�P��*jY˰������+�\0%y�ٜ16^��86K�Pى:���k�u�UE�� hgX)(L<!]� G(��΀!.1���y�xG��,��lw��+��L8M�����]OU&-�"E!%�&��ɋ9�$%ylX4c|�5�Ѭ��PU|/�<�� ���b�߄7�2�>�E�Z3+'#J�3cҔ��6}]t��s�̲S���6�B��+h��oi��I��K���Zy��#�{^��aB�Q�X?���.�&�����q��7�\[���@��G�SQ�&?�W߫�63BTb���9킷����%9��
�F����g?U����\Σ.
�ǧ�>��c�g7n�0Ey���|��/�7vF���ŅXU�P�L���ZN��|�����#-2���sd��FF�%��@\ѳ�[��p������:�;��;�wޝ�%uA����Mٟm^JF����"�ý�����<8 �V&��,f�N�є��GU�ı����Gh�q{{{�_<���� ?]\�T6Bes^bX��0U;�fBd\�q�OFf�<�U����ls2����?��_|���#��m�ϋrytv
��|%I���� �h��w�;99�����N�>�����@E�v:�)�G�p��t{б^���h|k?������ƴ&�en����ߵt��.^͏�r�3� �ԍ�>Ư�9�_)�>�7k+)�~��ۮ�n�P�U�\z^2�kU�"~��_��OB���L`�ض�{��Mw��x��8ŉ�8^�L�!�:�����+LeX�Br����R*��j68N�A�0�!y���R2
�����$�;���N�2�.����͑5�T����6b�De"�bml��I���r�1��l��w�.2�X�sm���㫧�@�1+��m�:�_��Mw�F
���Ǩ���Hk�s5h-�
�[��_[j�
���k0k�x���ډ
 �;���lLW�JpV�����"L���;	��ak��_������/�y���r���>|����g,��y~0b4��j�^oݽ�������O�>�r�l����/?���b��^���D8^@�d����V�4hi�ܾ}��GjAr�#��࿘.O���l���ف�z2��9THW#.�������G�=���'�n���N������.�E;���\�x/�t���Ś3h:3�bS0�pz^����@��LF#C��
��	�.1����%���`O�6�$o�����9�6��p�iI���4���0h�1�<���A?~����������D!zS���*���9>t	�^"��O�r�*����D�fet�,nl�@͍'�����J�g�*h����,��cg��� N�kز	uf�X_�c5>���+fs�pP�.�`s
���*)���":�!s��[�RY��wj��q�	�S�����Q�a�����"+ �#p�.6���K3�`�!0R:��*N(�qX������c�w�G���z�u��������2X��#e��Nw���uv����V��m��.��\Q�WX?\��h_\�T.��!Xc��x��OpoVYs���+�t-�8�����cu�������[�����g���X�=�5O�HJR)�6���ꢶ8�9h��*i������VyI�v0��qpp`��
�,�Y=�_��)�7�vSZ#G5�i:(���ȍ�)48�Y�Xi|��БLY��D-+.NWƈ2���
̠I؎�Q�~
جԊ�Ք��u��9@�Y0��Qo�G�%`vRNo�2�^q1A�Ez�q�͚n-�Љg](��"WQ,[�\.:�D�=��V�`�Ul��Q���"��*|���_��c�y��ҠG9�3 2\�7���2�eur���mB�2��������;=��z�����j1�ܿ�V"Ͱ;�\;;��c2�_Φq������ӓ����_`�m�H��vE9�LE�`�B�
yT����j���}d �0�����q�v@څ]� ��ޠ��h���;��e^,
ܨa{�� Pl�8���e���v����<��=��'<��=4��Mn�uK���������u�>�M�P����4�l1�J��N�Fv�<~����>�h{4|���֠?��띸�	�M�
�@�x2�O�y��,�C>��?y�R��n:t..F�[[ۯ^���;�a�����������#����Kƿ��_�����xk|z|<��޽�t;�������N^o��'�e��*�'��|l�7ߺ(��?��_|���7��|�gT�4*Zd���#��[��,��8Pr�s�\�m���:�1��4�5�>W���Ɩ*Y)4Ӡ�S�&T��T���2bytdZU�]pS*v�����S�R*bw�[1�0+�0k�G�0z$�+���?[��X{���V,�$�	���ϸJ>N�F�M.�S �"'��(B�H�np�D��*��١a^�mC������1l4�E�t`�T�`lx/_>x��b�ΣG�@N������wAL�p�n͹L�p�%�� L;�Q�.�?�r;�9��kµ���XK�S�� �i�!x����B��s��/����w'�|���JC��ƥ���8���a�dS����'FHJ���Ŀ�+f���vy�V���O�*"F�V?���$oS�v�+I^C	���Ճ�ʾ-��ē9I�''1f����a|w��}Z�"�������r�H�y��h�o@��6�*_cQ�]�k�YR޿�~l�:�3���t:e0d��hDY�	�j(��imC;�M����Ռ3i��F�R̺7�Y���^P����\{yy	R9g �F��*�`�!�6�͊�v�׽{��e���3�(�h���
b���人D�^�T�ڬǏ��G�j�
� ���>��@�qs� 4�K��1|��sT}k<�zu��M��w�� 5�5�b�<�����ܺ����Ϸn����v�у��s��[�~���׼�H8Ԋ�p8�{�.H���Ύ���ܻ���d��GJA8mHp�g�����cY�Ʉ�k�R8��<��1U�3�UV1Is�eecS|#z��JL���	:���M?f\�xx����&�HWE��]7��	�d��9����e���z�$��X�� z��Qv�t`���C����8����m�B�J��O�k�T�N��Cn+J������ϟ߼�-�2���X� ��/��9���p��5]a�g\�1�J6T�	e�n�W^��A)�q:"*�J��|N��8q�����>�3�l������� ��t�����(JYe��l��XV�l�o("�Y�*�nMɢdt7ݻu>_���Ǐ���%K�d�՟/y{�&�T���3!��8_vp~E$����X�Q���Y�m�jUo�5^Gik7�o��)�%��;Y��;S:�DS�y��-�@�uܥ�} vx`Q��bQA%]�e7��UQ������N���T�"x~�`q4/���F2�A�9f������K`���ļ�h��W���N��K��֙Ρ�K8i<���ON�s������B�TEi<R��Ԝu�9�D`���X������ݒ�x-aSu��a`Q�8��AH�$�u�-6|x�n'9��89?�u��orɯv,.�X/��+%b�䟃�`��yYfd����	l��2�L���ٞ%I��� p��>,�XvB%x�9�'��+��[�R
0����] �����������7}�<>>��{?��������e�/�����z�w�zE�/�5�	8R���N�w�N kww������P�Dʩt�U�3��u�e9�.΢bH��e���JUP�.O0 � !*��x������5�ay<Xr��f�'#U�^��L9ZS�����X�q�_3�z�sjJ�l��t��|ܐ[��Ì�<���6��1(��kc��FO��Mkŵ7��n�|����O����%�/�b��I8�4eԟ�1��Xs0��YL������b�ǁ�`�p��<y�A4�.�5[��X`�_9�3�loa%8*ndJWtwɘk�V��$p8��6�SCF���{Yj�l��1I�-J {z�N��-�Dy���l�u��w�1���+����U���Ц'�	���+S��3o�M=���4�����=N�ED��R�xKR���xS,
����v�o������Kk�����Č`�h��m�J�հQ��3����?�ӧ�~z��ͭ�m��"z���<��Pfd(K�zd0 �3b/1�c��ׯ�[!��k���R�~C��)�354]��Hs����6s���Iɿ��4�*��"��IiX���π+8���n���G>���_��_�4X�� �*9�@s�N�gƱ~�#W�9Mb��`�xR�I*Ʌ�����s`I���+4���s`[|��[�����/��z����o��)|�裏>���=x C1�B��eTi��?"��`g�F	��JmQ&�vd#�Ias��(}tt����ߊu�a�+Y�`���<2i2�����p���|�*Vk�� 8�sɍ��K�����u&!?(aWV�	�H�Ŭp��#�_I�1~��药�lX�N���zaI4��v��aw:iO�]D��2R�V2L�4�SR�Z�8n�?2kH�g"R�jr���>��G������/@J`8�݆9ʦ7_���!JLo�X�X�SP�bJ�B� �)?�c��R
�KQ�34�S}�&��\��� t���߽{w8��,���<C�&¬?���UJ{��kt��!k�c�'ak��`�U�!���lO&B�����h��~�hIb��)c�𼯴w�0o���v^��q�]��
��]8U�ߏ������W�NUn�I��+���`� \f;R��X��5Zj�|�e�5�D.&�ū}��I#�E���'��8��x^%�� 9��Y9�d||t��t:�8:X&:����gO_�}���?\�%�L��C�G�Am
��j�z�>�WT��s	p�,u������P�D7 �yd)ܾᵀ��A�Pu��eUT�@Y<Wrv~���;{{BŚ�z�g��i�����IE�hD��Vj�<�V_����%'	�6�S�?�``����޽{O�~		N�b��S&�@�-}�)[i�i�/rk��rrr�	vpp�F[8n���CxA�|�k��g������_���/���?{���#�w��� o���DD�VD!h���/�$Qi��͗Y�JhJ����`>M��b�JS�2͢O�a������Y�^��J[f���d��!(? 9hW�i���;�mZJ�Z�3E��g�W"�@Ƴ��<4��ʯ���Y���kU`�2h���»��R���ƩOB�W��W{c{���T�uZ����Щ��ޥX�#Q���{��1M��=a�����	̕��$C~cp$ �4���̅�X^��Ǐ�:�떣�X&�v�R3g�2�R${K���Kh�ca^0���	�Gh:�)56#���]�Z@��l��%����u�ȳ���^a6"�@\�v�Jॱȵ�L�n��$|9�{e9�íЯVe+GQ�8|!~���)w���E�'��!!������&@T~.���:dU��'�N?bMӚ6[Z!E[Ђ�JTڢ��;�e0�*,�u&Q8�Fe�/%�Y���w�����Zg�e9���{�߅�D����?��S@�A�юB�����a��*�e��	p!o}��ὂ%@�v޾i��,�����.J^Vd.㽓���UN�u�߂mp� �Ν;�^VY�8�3�i�����;��ћ9IYy�x$פv9�ۼu]��������H��p��?�v x)�ɗl�QY/++J^�p���)�_�1���!t�aw4h
`���>a78��^���^������w��]�����{�l������ ����	<��r~��52
Y����hCWafcL�;�l�)�Fn=A��܂��c�
&j@���ћ�:�u���A�sF��J�ov��3�8E ��s�/rP,L�&QTXӊ!J\˙�8�`f���&V�*�J�]U�38-'7*�I+*��}j�i��lY(yvrrv���Fhba��	����4�(\����,B���h`Nlu<4i��dz�Ī��E���3��0�n�F�����l[t�����	��ރI���|�t�������&���=[aϳ9l=7�wF[۽� 3S�q�Dxl]r�2�����ɗ�nݺ؅����y�Ȗ6t�R2� �����b�nZ��ǓKFZ �n�[ۣ�,T��K�VG�E	����rknf�4�����}����E�=27�Ɣ�E�+��^�xS�m��'��J����6�p�^��%��4�6US�r�=kL�_"�Zś\��k�M�"vi��01��u��t1�S����>Q��y�\���&}x�J��R(+�����b���d;�ы���w�tQ>}�x���I�j�&p_hd��\;�M��x<15+J
���LE�m���f(���`�6��|����Sc�{�a��kɞ��Ay7���z̢`8 qw�,y�H����Љ��l69z�� @Lg 4:����g��w|J��T�e���j�����}�1=�saܾ{���h �n�VBB*^�Ey;�z�F'�xW4�@���a�{ǹw��/v��7��?�p�y���mw���ݷ��~qt��h@�Ы��3x}0!1"���w|q��уW�ǻ;[��(q0LA*�=_L����4ž@���&j7M���'�7��{�ݓ(��f�,�!����CW;\�
�/'��P�:@�_җI!k����#E?*/��+H���z�]�H�8�|�i6���T�`�n�e=M�y��grEo�d@��SW}�����n��<>�	�<G�i��IR|%��U���}�k��(A�v@E�Q�A�My����W[�������o��oe��i�hf�m�@{{{0�����l���������I��<<<d;�+��X���p!,ί�B,	*.;姃���g���ȝ�wa �҂Z1�{�6i��i�\@#܂��t�J���o^�r�q�a��=�HeA��J���~�{���̿8��
�9x>p#�
�������T����*�h
!%%�n��TTu����4�Ɣ^�|���:Po���׊:-���pj��y���Hi{��@'$�����"���_�0�	�$v�?� +(*���qL�?rI�dk��g�}��#�Uص��s^��p�s�I�U�Sok�0�x�W	���g�*F,��>��B��hn��b�u��M�|�&�rY9�+*�5n�����}��?~��ƈ�0f�#t����'���ˋ\��iH�u����^,rA#|��v~~���%�����a^No��8m�Ju�@���ڣ��<����ϟ��3PVjC�����<|��Ν;[�4��/�H�S xwO�}�t�/��C8����O������|W{7��c� )��������B��i7�ڋ�����6��=���IK#�@ 0�񮻧�}wu�Mw��>�_eU�@ج�J�e�k����x�+OV��/nJ��������k��R �D|Y�K"���M���,���CJ�A���< 3�@���ɾ�<�q��uZI!����z�r�K/���?��Ir���7�J��d��=]�ʅf�,b�O�ɯ5��S�'f�_�䢴����(_��q`�%��)_�i�71�إ��I�(8^A[*�r6���)X�5AK|�@�F�{i?��+��Tp�����������nD�d�+�����`G��qo��6h���ߧ��3�fdV`�������%9�ؔ�ӕJ���ܺugrr\/-sm�Mc{[b����5 �F��f���2�B^^�v� ����9y��G��ML��x�:~�(�a�\�ȩ�,��(���������۔nj������\z����Ȩ_(��=04�t{�Z��&��R���1�Vgrr�ĉ��奕Xk58K���$���g͑?DWG}������\���Q��1ݾ�(+{{Mm�(��O��B|���R�% ��lw��2���a����gjzF��V�݉@�:��Ɋ+Mf6Xj7�.%�RX�zL�aN���q⪼?}��'�xچ���é|��ϥs!|\琊�C��@���/��~'��s�Dƻ��uHyi�~檷ֈyJl=��9%������O�fP��e��TV�Q�� �M���
�*�č��C@  }a��W6�֓8�vZ�Ϭd���^�H���Q�-���`�z=�E��}��ZmTy�Eb���U�82"S���?q`3N�0���Sإp�����h~0H�Q�o(�����Dd��ġ�� ����?~�Q�x~s߯����͉�Ѱ����>m���C���I�ˋ_(1�ꮃ��(���������������իWp��� i{���[�I����%V5�H򴶶� !�@�m�2Di���x;�z�֭[�	+ǋ�ُ��۷o�={"qwwyyy�Ϝ93>Z���ND�ٚ���ދ/���˯��g?�w���y���˗gggq�����������Ϥ�[h���+�����:'a}�Vp%������u�2b)���P���7 U�/��>Á ����Qpg�%���ͦ��7�X8�S�8ϒw��t��Oe�G2��ʛT�ï���x%#Pg��P5�*e���?{��k��ҟ	��{ ?�)��S��?s�����sE7�6��
G<b�
�0>��?�$Gy�m+7�f�uj0R�(�Zɇ[��B=!�mJ) s'A"��V|���'@��?��'ڐF�g-$��u�sAa/^d!|>w��-+\��4��(_p�ѱɴ��6���ƙ5{��^?d%�N2"��QdN>7�� �f ��	���Z�b�D{�b��6����%?�-Z\�ˀ#���=6n'�fGw���Kˢ�
ur��9�N;n��G�4��~և�XzH��_Faċ�zlL'(����9�x����Dn�;O�y��و�P�i2�;_�`d|�ۯYɪ����s��T����ߡ<h��~w�������kz��.#�ȧ����p��L��U�&6��V�������Սmh�(�$�jM�%�e��{i��)GYգ��[fW���)�Ԃ�Ŭ��9aX.
)��׮]ct�z=�P"ԣ?)�*�g��̶�'Z�6Փ@Ȉ��w�d5�Xn�!7<7;%�&u㨼p��#�����,���<W�z}���O =�#�?��>-<�S�N��l3D�Y��`�Ɉ$�Y�x�l��_���Oǎ�°û����x� S2e��:�Þ�޿��	%T��J��S������K/}���89�0NP����3SӸ��N\eC�ё���*%i����� *��6��f��f[��mP��IemS�,�(�eB�q���j}�A'�T���Avx�6�E{�C_�.:3������,���p0��hK��-bH��sp�G��Y�������S(]�\&�{"WN�ST=�I&��Q+�*j�T��ft�V1�����BQ�w|.�����2��h/wp|O޼�%;��w�n�nm������3ŕ�*^�b�\�7
���;��͛�O�r����TCf� �fyV �8������>�o���8��loo�e�3� 019�0;����۝�S����(V��Ӑ���KU_���wZ�O;��>>�n���	'G�<�"1���n�+F'��=�)c�
�8�;�^J����׊�5�2�����l�S%�謢fy
��4��u�)�I�*w��i�QynA0��{�"JgCa��JG�������v��C�xb��!��l��䓑�Rm��mV�de ��X�æq:;Y$�$�[��*�� ����T`&���7������P|(��ڙ��h����nC^��_�����{`[Z�B�'T����A�ª���E�#��D��U#؁�5`�N��hO�{EmI�WH�U֍#�v?% ���+/�t���	dA��_}�o���sz�ܬ>������1cB�i�`ŝB7N��.k�|Exs�GN�<�Nf�	!����N/���q5J��O���|ȱNk1a�cN񝗊�>��VV�{;�M��c���;XU��W�����DL����$wEѻF�TZ�B��s�.�l�zn7��#G��~�ӟ^�t��W_}��	�t(@�~h:\qmm��ѣ8�������!��'N@��'i�2�z��ŋ��f��i�,/Ý<sfzb����P^3㓀��Q�[�T�_E�I�NK f Cz
 ��n+�ח���C'}��eE�������gҡ�����n*�I ���t��:�?qy����E���D��2��]��E�3����4S���YHsUpp�����fȃ�y��uR�g�s�ɗ���sQL�y���ԉ�L6��qs���zv1<���B���������/�*jX˛�r�����\bg�I[�@�X���������[^^�����@ǀP e����4��J������
P6-�4��ͬ�x�9!�]ò>|��7r�ՠ���HM-Rj�(F��Ǟ��J>=�0oC�X��A���Z?s��+%�%b��lU!ij�W��1��#ΰ.%�T$ĩY)�M"��͒�P<��Mǧ�d�,�BѳfztIl,����R�5��=�#7BM�M�i���df�ey�ah;�}�|����$�)��dIA �����܁���n�����[����s�$�塱�����G
���`~��U+���|g�#̦��$!�K1���"�f�� �$��/N�}�̓����ﳈJ�\(��������;\�x��Wn^)Z�W<W�oJ�2,g���`���T7��1O��/x�\[l������Lur�����.$�dmդ/�K�"�����O�ߜ�ˇN4�
�ZK��<�kkt�aP���˕"�Zoff&���n��K��i�-@�5����k�O���9<�o���_?� �o�isZ�0��^tPm���Ǐ�ܺu��#���
t���ױ�˗/cO`;��ʏ?����g����G��gV>y����Cр-i��~�N�rK�FcC��b�2���)�8����8�#�"䝔���į�-���q))9�M�v�x�匓g�e�f'���.b6[����<�e�69#�.zhe�{�ʳ�&��k9U�?�}�}��~E����\^z�X�K!�4`��JO��ǟk�t�Ѹ$�\e4\{m}�\��ϟ>~����H�������b�ٚ���zښX�������" ,��g���
2���r�Z�������T&<j:�î3D����A=HPJG�q`�,��&�ji��F�ǥ�jK:A�{N��ѫk�� �
��M��L��
�'�|O:�/�cqZi�Q�w��=Y�����Zu��R��(-���,�?���Mo EWߑ��.����*I%Q� ^r��ׂ�T=x�$�P�����h�;0���h�/�ɳ&W�����!}`��J�'#lb,V�&�S�	�Fa��J �j�B��F%���ʩ<��9�� �7��x�3|֧@nB������v�e������v��/ݬa2�a`�y#V��e(��pt�=��^itt��侻���"�La��l�M�^��b(� ��H2�ӂ͔ΥG`����N�T��������ki�q9qbڟ�
em3+v����<u��L)� !qH�@;�sbڟ;H���I���F�jaz2&8j��7vvw��")h�d*i&0��*s��'-j��-iE� J���5�O���������T�/2ƍK�ON�M�KʥEJ6h�ڝ�-�7�wjj�/���Mߗ<�J�oOcye�hnn�ԩS�o�&���Ű'5)[��B���L����-�����Ѐt����n����D�~�99)����5y�A|��]�H�uW�y��.��SǏQㄬ����T�b�HK���&z��a\Iր�V��Z�I���O��\?=�}rr�B'DzG��OQN��y}~�؈_��i��ͭr���3���*";Ԁ��+�YB��չH��s����7'��}�SMLL����pP��ibr�g�&+����}��I�Ut~���r��O~�Z� ^P�SSgϞ��O�@fƁ���ѣG /�?�k���±���jO۞P
`��������q$e����uڠ8�}�z��qQ�Jja�na��j�5{�m����J���/�s�*p2�2�O/�HU)�,�u4��S�lGGZ�����'^��LK'(������[�o���D��׭�����.L�B��6���T�]�9���y����8�aW���:��d��`��f�E��կ0X3yn�D�3i��$���q|���I����m�S�T��w�>�p�)0+��78�wnK��@m��ʲX�c�g���>?a�Y��Y��hҤA"�Ȫj社� ���bm&�VX�t_0��Y���=�:P�a�t��.+C �����%Ū��z��JC�;Β���1}�X`?�IU2�S�q�,��˚�ӫ���t�U{�қW�	4n��u��H�y��*W.1˕x53�IZ��ִ`�0sq�a����%�UJ̨c�#�ő#G��;c���!� � R����*K�jc�ƂM_YR
|v���sff�رckkR�x��]�}$����pq�I���|饗p�{��1o/���Ve���o���C8Ր���U�E�Y��L��f��(�q	:_l!g١��$ff�H'�8-��Ԟg$�e�i8�=����a)�|�L��խ�˺��ҵӪ�p� >39�d��G�J1����^/�R�e2`k=%�%rM�۞�e̖�ɒ�B�s:��<��A�l�qu�5�)�&�1�.qr�I��A�<�2�Ӊ�ݻ������onnFFgT�#����k6�g�X4�r5��0<Âa �X��1�GcNs��2f-AJ�φ�i9�Z�U�e �P���&ȓF��ptH@���yp��ZJ�, ,�Z-�mm�]!]��/9A�jv��M��M�DR��J�8�!�&ZBJ��^2�ef�SwZL�e7��S��@�o!K�$�hv��G�w�1�����$�^��'����~�#,��g^�@Ҥ !IKO��r/��IN�̲ wH�%�a��z�-��1�	�&R"SPd��&k;��8�h�4��%�u\P;�w��Cˠ"�����瀛�l���k;$�Ռ�ӱNQص���1��pB�f�d��my}f�S��愭p�洱��`����`f@y�����R	˄��!훺�ה��a�1�h��t�Ju�� ��Օ���H+�T<�H�
��qQV2�:$�Ĺ��K](��K�cch;��<�%6�,�)s��9ma�u4L ���Hr�#=�!����=�8��2ԕQ/ݸ׉��vL��M9�̤L|�I��Vq������D����Dc������|�7�X2u� @����f�Z�b	Zo�ɓە���d���#�����yh4|u�8/N�q���'O��8�yϜ9��oܸ��'�۟}~���ё:�$�;N��RY\\~�՗����g�6|���D*��V.W�,��v��/SKM�K~!�Hf|r2��Hg38�Pur�m��:���9i��¯X{�)�K����ɬJ��?|pr��)�ixN��ʔNz
qŉ��Ʋ���H\/u�螚Е��S�?�*j y9�mfPO�w�<0���t��:���z�~M�_ˠZ�3l�%y�5a���&�ъ���Y��K��X}�Wp�K�.޼yP �>+�v+�N�ވx���g�0�����
�3��bMD ��Zc n|�S-.>����8ȝ榀��O�p���1��P|I��C��������=�ݓ���������-)h&:��2�W���D,�2�?,�B�4�Ry��r &�}���p�ܬ��� �u������g|�{�Q@��Jx�O,�Ζ�z�Hg���]~���{�g�c�|��(H��T�#�#�����
}xIh�P�,6�9|L��;�_aДg6ɡ�"�H;�z�%�� ~�T�m�Rax �C�.v�F����ZB<ynZƃ���t��-�$�i��ͪ�8�|sn&�ݻ�p# �f��C��СE(��	�m�5IAP 3�]��N��n�2�d��
�w��-���0 e��5Oòad���g���J�ݬW�Q��M����R��,�nR� qF�-n��+O�u�*v:�0��H�|7�X����q;������!������}��d�h�H�V��!������6c j��ѣǢ1�RJ���oǚ O��^�+++@i�����kװ~���������l�|�M�<���@%v���X�6�v����Q�S����ySom�*�����
Ѣ���Qr�:��������eSS�[���53x=&P��g�Ri��$�k��2s=��r�'5x�*-�cW/]�Wki�7��P�M,4�Gu�� I[��o��yگ=Q�b�D=1L�����d��{(��Dh�?�	z��k$�����Yݾ��"9��ש�Ԙ�Y���ڭ՝���O &�^���֑�f:/<O�M�e��G?�ϓ�c�9���/����ۓZ�&��h+�Z8[��OMM���%ˈ����5,�����s�WV׊����c�::.7ɂ^]-��T*���x�ۖN3���[#��T��h[z���cG�S:tۭ��ܓq����G###w�V�������j��M����v��� ��f��n��J�T�6��B&��f�{L��K-��J�"�ߔ�"rz�jJ�Sv�sh�ڕJU+l�E~�0?s���rud�xF]}8g�� /R^��2�P��dh��}�U�P��d��e��t��yh��Nd�z�h���O�4��G����k�������)���vX0�D����o�ش���Q�Xl7[%P���o��6_$֬D'\-w"�!K#�}*��\��I}��f�/��$�!+y�� ���:����2�V��nbS-�;{�n��?~vf������רJ�^�U8��|�������g�Ad����8��MH�X�O������r��Q,��� 6G,u7gi�G�i�ƤFI�͏`Z�{�$�vb0�+&�����������5;7�����oJ�_�t�q�57;�Ǐ���O��O���>���B����'뻻1Pr,�ޖ�f�bt�q�Xҵ3$��?������ޞ�D������R=Mr!�a�{���4-놞+0�9�@37n� �+�ŋ��~t�+��=iU�6n\
!9�R`Y�f��n��_u����A���Z�$�m�>�L�!魛������Qk�+�P�(
�	�ݿ���w�?y�f����u6q�}Y� 굷�k�:^=Mq���?�����xfbJЁ���G�Ց��<0R��<?�ml��I���wޑt���������3�sR�V[|�P����~v��Q���L8u���#G�H<tz�V��E�_�i��%<���x� ���ޣ%`h��������/_�x���+�?��?�����?a��ĥ�ƞƔ�xskmrbg��Q6Ru\��H�_h/�E���_W\��R��{]}&��C�1A����]υ�O?_%]��Mf�ԳJ�S!�O+Įu�8i�A�5��8l(Cr֞��[!�12:2����\܂I�n�p�$�t�vP�}�dͫ�ٜ\ ˪�8����Xf]&�S�Y��H��<N��a}��=6r�
��ɪm�SҥDp�g�Ӧ-mr��]g�V��s��e�<?+��>|���6f�"|	\��ĉ8-m�T�.}�~�j��b6᭿��K�'H�.Xt��T �>$�S-T{��Vj�#�^�ɡi��|z�Lyxl��1Mt��0��h�tv��0��T}�ͩ�N� �'�}�UR��v!�
�Z��O����X���W"���V������#'o�$�*��Ӯ�Gq?g]���29ɲA��b�̢aD�#LR-p3ک����B$
��v<�
j�YN�\/��gy6���c��7�->���ӼSz��m�Zd���_�yO$>⡩�-m7��o��o��4y���k-�HW:����T�*4����^� aX�$u	w��I�j]"� ����x�5�Ǫp�!`>ܾ}{iiI��+k��h���mb�8J�^ĵ���0UuZ*��h�I�TL�x�J�*+�rb7H`HrM��Œ �!�m��}���D�i�7�ϔn?���l׉�Q�C�'&G{���߭��ז�!��z��g�4���-c��ݖ�uI;}�4V�HW��Y	Π�$���$�E&��z���o�k^�r�
���޽�ڛoM#��|��G��6\�[�� ����H�B>@�����
^�9;��_��3D+�����2wn�x���N�s޹sGF����z�c�h�33%�8�N�ŵk�pN��ve�����}�V��\:V�U�&�*h�#"�$��d�^�)�oI�˺o&����8k���z��s�Ϳ,��<Gn��&��w��$����*��?��� ���YgԤ���ߧ����N���G�X����W+���Ƥ5��T�M���� �a��5v�߿�z�N�u���	�#�W������^�:+�+@B++B� ӿ��N�ݪ�$
c�X�λ|�2� v��5���Q`/fu��e
*cp��� �1Gۮ������'ƘEnTM\���'�'w������'I�r���̩S�6�l��H�A�l\��
����%��>-��s+H7�z�3��?X�`��ݞ-;�ɛbvKߘ��7���V'h��%�T�Kpf}T,I�l3����CK?6�גM^�0�*+٧�
{�l���m>���r/
�4'�1e'^�#��^.�:L�� � �<ߖ���w;�X�MG� ��.��Ly�O5�+�����c[�U��)��3��0���Ķq�šਚs3)�����<��R}Z�������)�l�H�X�i���I.G��W�V���f���;T՝^ww��ji��R�9����0	.���*��n��<<�Fcǚ17fp���$���Kp �� �S��R�~����+��ζ �9%�� I��m5����8�Ȉg���5߸���㉩ɹ#���=�^;{l��]{�����.�/BR�����+��K�&�S�m��,f15��NW����p���߇4`含�b�'4n����A������^�z�;���x�\����YXXx�w��R�'��믿�7�8�o�y�ƍ��E\��ٳ�Ν�ـsba0�_~�򨎨���4vv��?����P}%�Teɧ�d��c$\�dħ�	[���w�f�_һ�W��DJ:��D!Fc�q�a�lc��}�_�s����E�e����Ch�K/f����t�,7"M`�2^m��d���9��؉���*o���1 ��R�$y��8>�S?KH�՚�3�$׾�3Kpo�>"�Σ�#�����$�����~��1� �a��PXz��	� n^4������t�� �[_� -�1�	&�V@���RW��� sLit�I&Ss��T[��'��{�"���u���{{���5Z�8�Yb�
�(m�aB��H�Y:�.5@q~�%�&�˔V��:�yi�N>��X����-,�_�_9Q@lJRA�'	���%yXp��ZB��*�!wi7��i�n�$��e�%�"I���-��xZ|��3���cj��Y\��f��в]���O�0d�?�'���Y��V���r��������~%�[���k�P�~�$��X�R�э��CI���vlv�&���~[����@۸Y�.f�f���=���źo��eg�7`��H��C��	��AM#�T��6H6�hz6>U�m��&�~?;f&��2e�/ʛ\V�f�z�SzMN��$!�.��(@
&�p\�m̄�X�e�iY.Mu�%a:N�(�zw�N���a�K��uW����.]���ݻG�d5�惾������ ;�)ћ���$	J5
u����ߺu�Yh�zc�p���5�{@��f<x�lHz>��|p��u(/���tX*�-tn'��P:X�p�ȑ��%�q�WC|����������4�H|�����w���s��)3f�Cf:kƲ�@�I�>N=% �D�x"�(�n�A���,��L���5+n�IS?�ge��'�K�o�W����m^��	�K�3���	�>�A�eo5�m$�^��y~g�����l}|f�i�7u�zF�@��iY�tU�IgW�#����晅���7w�xa���k�Z8{��!��h`.�X��@m���*��X�&ǯ>��Lg4���;Wb���d��_��VGagH(�M���]_��ښ��Ao���fa	��u���oo�	��@x�Dǎi6v�����@�ǎ��no°ZY~<7;!d	PX�������j7�w�JQg�-Y�S�(��ʱ�6o��p(aOB���,�ih����Kfk�׎�^��*���i�lZ�هn:Z�P:N��y��$�p�B�8�[����YlBzW2�`rj\=�m�� �	��eh#Q��d�D�N�髄!��:�����<;�9� n)YC�����U;�N��ɣ`v���f�b~�OLL�&�u�����O������m��;5�,��<��4�A� %o��w!��E����+�v}ʗQ��m�\�t�ݤ'����+�����j�Y
�q����[[;�ݦ��	���,ʸ����^H8�e��NK�TCQ�6�&�����{\�h<'I�k�Y��sQ�2��P�,-W`n�21�pDG��srFK�X���¦�pc�zq{s2��Ҳ�O�q�"�P��G�hI�1�Z����n�}�s�<}������wv7��<����]1�w���zajf���*{���W�|��ޓ'O�}N�>���q�¹��U|3?;���W��N�<}����v�3��٩im�	x5�@�'\��?�1��c�$`)�����3g�`<I�+�/T$�g�P:X`"���Vj:Z����6gP�<�{�&�1���C7�յϙ����=UI������2�z���ݴ줕V;��fr���P�U+y�mi�OT&M͊?��i����aω̸��=�9PGjr�m�]�7�����YJ&M��~5�$��zɹR�~�oa����Lqr�4&�h��B�X�W�HV��c� ]�B�p ���Ĕ�G���g�a����wa
�$ztl{���B�$ڏ;���y����ӧ�t�|����n"@u7n� <b�YV��:��X'�΂;�m1��X�b�5���s3��`����x�8�＃�OT�Ë�ìl�=�Z, ֞jǏ�d���u�y�����.��f"�QrD�E�swW�v�8&>K��Y6����ƫ�rK^Z�di�dQ�$��4�E�Cē�a���ƹd�$�Z�Y�cK���o9:��M��5��Tl���)�YOc��і29^�L�S�O�7z�s���G{-1�_*6M��y"�
ænP-�ۚ��`2
�Ǡ�����7�o���ה�{gl�$]��+�����r<��Ē�'>M1�2�%�r2�czZfi��k��嫷�\��?1�K�ڝ4�H������^���y!M�g���<���|I]�kOˤy�kLj�q� x:����H;�3��V�QPP��n'�^�uP�xʭ��t��=���b��woC�����+.����^/P��v��x����;S��c����f��8S���Z�/M��*����>�������o޼	��/�ybf���qǎ���ŋPj,,��ΜZ ���B�1������?��O��P������׿�5V��+�@�\�vmqq&�}��0�n
�3i��_.||���{<"�
��1qmjإ\�H|�����җ[[ ��_�4gF�1�|�9�a#�tLg^��~Hr0�h�Y�����/EV�с_�B��+�Gwc7��<�����s�ֲq�\�����w���\�7IL��MNuz�^h+�%+�O=�mA 8{����U��f赥p��&g�������������\
{2�r��ʥK���� ��w�r�%����S��;�<МR.�0K�5}�r����ok��9E}ɮ`@oX?���
d����I4g�sf�<:�V�|��uV}�Á��{�ryfn L�`^�kk����Tؖ&ц��;��`g^Q=�f&��%q uza�-���q�T�̌����L-�T�p_܂�c\�\�|�ZsG�8������L�rK<�h�R�j�$m[O&��
_�'���J��Ό�������D
�ap7]�n6q*p:'�HG��$�1��u�|�,Y濷���"9�������̧H�a�ـ٧��mC	�*�^�YUK>��&��k�s�TPj��:|F�4
i��gY��~�:	3m���&�c<P���Z�eI3�#����������GHT���ц;&�uZ��7�q��ړ�43�����$���>�8�	�h^_��`^���*a:P�c�hU���9ͺr�Dv�`
%6��� (8�/�.�4~WS��@��Q�"T������b� `H�#�J���߾s������''`����{vvQo<y"n�J�!^o�x��J�ʩ��;�����-L��hW����3T������]�������[o���7�Z{%����_�ځ4���J����տ҂�T������M���*�ә�8�����|��y�#`�՟����i@c`Ꭾ\��������ŁX����N��������?@��w����N�<��s��]v�N])״6��]���,J�n��Q�\,�e�ako���P�����-^����v{�maP4�FQ�9xs���6�g�u���$�������zv�x|���*4�*��p΅`r��~69?����Ȳ������g�kj��[e�s�I;�L�>�ss��)��[�:���"ݭɭ[�z�������������
4'-��� ;[/�����h�~�)�-�? ._���J�*O�C#.Z����7�x��ƍ�Ҟ�͹�|�	��㊌vs�X�`A��Y�	K�F�/��^���S.h#��}�{���t ԍSG�㼁D�`� iam`���	+a�
���\��i��hiz,���+��Xm�������'y0b�j����fS��̤�+�g��yz5f���K��fۤ�^b�ɢ��.����#c�_l�@F$K6�ax��(�Tmmw��&�Mr	CN�CN޹�P�����6.Jh��x�-�1�� 
ٽ�e�4��A�vy�07�!����7��ws��uKO2w��(�>��c�5	��g%o���P��H�O?�Ꮰ���g!	u�[J~���O��T�dh��(p_�^�� �Y3-7K�w�uB�\s�:+]�K:P.�S'vr��[E��2����6}όl�1ɌX�.��P�Z-�KMW�L5�:����ŋq/��^���HK�{~�����>E��'�[��XP.\�aG���OLY�4M�ٱ�	g�>j<K�/�����P
g����/O��������@���/�����_�nm?��`�B��Ѓa��@�1�������=!�	��]������;��������Â{:��:���k׺�ֱ��8��Ӿz�*�}IT�^��:��Y츳�C���ʊ&)�����8���I.�f��(��3�hܒ̨��ٜ(�uz��M�}pr�����;e�u8�r�I6��S �D�\�|�Rqێ���{�����=��阵<� ����R?�d� �\K��Ǆ؁��Mj5o���)L3���ʲ��lnL�>>?w����D+���>u
����?�t钌�6��ѣ�:��ʕO���۵�|��Ӭ���_���X����r��9֪�W ���-��Ըt�`r ���{�p,��RL��3S�ℝ���8�za��ݻ����+��Ц?�����P]���սW������*�/��I�#�G���ֺ�	㨐�ZEZ149>.��;=���5B�mx�9��8�Hs�D�,%�����\�Ӗ��$Q%"��:�� ��T%��A���i�FKФ�L!3�D2W�i�H:zX��Iw4��x�R���E~\����x�@LY����r��e���و�]W��@/�1�7Ѣ�|�5�`��-��K)��s�7Z� 1�N�:R������k�x�|�A�Ge�5��k� t<?�ۯ��`k�b��q^��ᧀ�AO�K������KN�?�A�c����7rѧ��~~.7g~�nC4���s^�ҕ�تB�|�H=���	^zЭ�*�J���ڀ�J�,�-� �����dR~�Ϛ�)�6��y���ېf�Ν�����ޕ&dmPZ9�_ͼ�(�Vk��O�����n��ۛ;��$���&X�c���R��3�$�=�&-�O�4��n�  �mQ�V����L�sp0��f;niR�;3W���J��7e���P��J�"3"�B �-ܩ��O��k�WǙq������^c��fblJ�p����t�����f�E�ή>Y�\���I�-LO�..=�Fh�e����(����sDΜ��֞<�x�v����_ ��}�נ��|����� ᢧO���?�����q��*�h~~Z�����v~+ذ���~
4�5���EX6�����C�} 3��;w�@E��D�5�$�9h=@�7^{���[P.��/�b]�<�����$��3�Z$���>LJ?�Ea����#E�k@��š�-`݀��%����n��`�"@����3em�B�+���٩陙���岴�1a����M,Ss*�q����i�* �җM�qβem���'%'���Դ��^��)��Q�X�98ٔ8,��r<�?�P�S��^�r��i���Y�� H"^�g��:AX�#f֣G��ܿ��#m /,�>�i��@s�n�±�	j��_�3(�]��ʮ�i�tbQ���ַ@�F89H��I�f	�X����s��l���
 Ұ����Y��JIN)w]x��2x@'�� "����N�H�r���$�})��ظ�

�
���ta���L�|L;�D2���,��f��R1'D<F�:%�_��7o^K�B�N6&�PI��� �%Y��8i����:
h'+�dT���NkK��k�,�3�W��>��XДd�*Yw�AL6�}�� m�@^�����U�����o����9���2i�r�xֱ�ݨ�c��n��j9�s2h7�O�U��l�"�!����9a~�!7��^!i +���,@Ar��4t�jO���O�H���/_V���� ��.6˗��'r7�H@m�K��m�>M�ء�K{}���q��;�������ش���'�|is5����{�O���5;{��1��m�|��N��JvCu��,��e�����p�A؅=\(I�o�]�p��i��sZ�;M+9�:E�&���܄Ue���p�@����������b�Bs=�{��sG����XZ�\ǹ7���Ϸ�z���  s��>���Ox7o��	�P��ز
��YPj���w���v�R�}�4����������͵kװT�KX�8�pB��u��ږ�sI\�i�mm_�j?����B��奬�s�n�@������u#���Y�s;��{���n�0�<�=��:�u��A�7�P��(��s�4���)�}�r����,_
@|���o^9�p
�u�>n�"���[��hS--=�!��5�{�}T�����FS�s���#8�~{?�$a߇Q#�rԓl�Z�
ej��1F	���O���= qi��-�u�t�c��%��S�^����)0>��p���i�a�tۓS�������xbbL[vE�u��taiaO����{-��p*�616v�����*�8I=MEJ�R��yjxVr������:�qX:8�~1��$�ڈN���T=�?��6�I��S�gx�e�k*@
5�[�m1s:�)EL� N}f�$�W��r2k��`"b�	#9>g����""��N�z�P�w
��n�M����J�S�>�M�`��#��j!&۴%�Y��<��yE��gr��(�SuR������¿Җ�)&�~��N�7���ZQ�����˼u�?�o|����JW�#K����/}��`+H�<l:&+7�Zg��nqZ���9��Ǽ{-�#1r��f$x�ʕ+��Vh�P��7}�R�?15561����V�Ef��)R��q�$Y-Qn=q6�|����L�;K5_d����J!��!���=�Vv��P2���Qq�����Jx�mM8�SZ�&�s&f�/]z�!��u�{p\���������޽���&�H"�~����Hｖ�S�ЉM ���4���B�A���ǁipw =|��ψZ��1G]w��l��7:V�:	�Օ�w�y��ѣ2�|v�Ȧ:�؎��1y:�����/���+�������_��Ȍ�)�ڢ� ��v�ţG��x�ٛ]ZV��PL_|�@�Y�����Uvw�J��V���Շ�����_����y��գ��W\�Z���QV)._�B3K-Ec�鸾�"��]�HA���A��|��R��û�^$OS�0��jj���q�d�$7�Ւ2�eg%Ba�X������D�pL�̜	)7���Pvv����9ۺ_U���{<uK+X�#3�`ey��3�f�ٜ�8�\����5����Y����e#y�΁��e4�s�R_XX AK�䲬�fR=gc���K���@U�R�Ѥn����.�E��3g�`�Օ'|�83Ϙn�р8��Yp��)�a%[Tc�0J��U*�`\�eM�>K���X�)��v�g~��]'K�L��y�'X��
nvC�]�Um��Z�<Z�F!�柁�qf�N( -zE����Ni!X���4ً�Ɋ��<�^8�%ƗE/T���O��Ӹ�B3��t�:}������\<�|�AZivp��&\+���"���ܖ�X�I���V�[����2�A�q�w�a
��9�v�ɡ�8�Vt�x�c�t��6a�D�萕0�� Θ��� ����(��z~������_-�7ג���3���~�OϿȧ=s'�h$�iݺa��t�����ni��o"�v�H��4�®�1h�Hs
�?|�k`��_����zjP��F:���T�D�=�t�z�l�����8��؀8�l֍��Nx�"0��K����)���nl�cI�U5g&��߆{)Wı�('&�I��juK���d�r�W�c�³��q�RQ���ʥ~B0���~��{�LGA�����8�n}��<:�]���J�����n����{ᅑ�%>=��ƍ�Ԍ�Ӂ"mz����}�F�ҹs�>��S<��^{-�.w���?���ӧq_SSS?��O�����p���Q|y��<j�K�8�|��;. _޺u�a�۷o�AO��itCi��t ���Juܠ�W��ª�OҼh�$��Hæ�:��ҏ��đXh �2���n��'\�dx�+���CP�r� ���f~�gp����k�8Y^O�eMiұ��r�J36G��8	��}0P�s���O��UiU�+Y|�Ȑ�ڨ�������X��'�O�ɒ�T�"���ɑ�q��%;��lnq�]P!l��������  qP��� �Xml�׿�5��M�쥳sM2-`U0�|OM\x��'O8����xV�>-��,���S�g`N�C?<����_�7F�G��3��X��3�%SD����:ч�	��L�Hy�H^j�2HV���8�+��^�H��i����M�pL��������$]�0���1�����X#���"5\��J�mf ����n6,B2���i�$X��c<���b�5�2�O*�|�6�p9=�E`�n�jv(�p����<;�h�/�~�ʃ?{�''v��9}��7�|�Kvf���@IW�PK\c(�8�H�4�ů�`�v�����də����36���>��!y���~�͂�8�(O���N�=υ�����g��́W���R��0>��L�Hԣl}i�K eZ�168���8�g������t�|��7�di|;�Ap��I��������o�Q�ח�z�Õ�Aݖ\G���� r<�(�N���!�k�a�%�D��8q�X�g�W��r
Z�*5���#i�f�l$ļR���*֎�4i�c�2�Y����1y4R�g��|�p����:q�������W�^-Wj@2�8tΕ���/��펍����,�ԟW)yN�JI�#��H�� Ę�˒��xyqjb��%VtϠ
n�6"}��'*��$^ZZ|pO�C[��֛l��_�����/]z��W@���lq0O�e�-���o��ɓ׮];{�,�O�S��ȑ#?��ϱ�?��?�t���;�t��	gP�y�* �uƱ�_ln��a�^��	 K�
���^�/�d�l(E��R�*�	5	wJ����f�Ō 1SE�\7�5N�k+����-8��XJ���LD���)�g�>��!���$I��T����oZ|�/<:W�%������l���|&Cf6[h��Q�Ϫ�9��t��@pƖ�QV�_94�v��NW�1��D��e���� J�г��i�8����x`9��|g2m#�[�Jd���9f ���1l����q8'��'�
��fK[��q�3��1A���--�:�wqN���։3�w&�I�F5FS�v�/����-�5�B�i�{+i�7pf:@[�-$w�-�1)8OS=7a9丼ق����+��59i_by�:��1離�m�J�d�K�d�#���!r��Ң�B�?�;����(k��N�\I�w���vF���F,3l�X͚����x����.5��#L����>����.���`�c�
~!1Y����o&-����͢ϡo잖��a��k��9�i�(ٔ��G;�/�g�lP2�����g2XP��Qy��DBmg� 1�Vƚ62��4��<��p��4C���Y�P��L���69���F B+���+�*�1B6��C��N�e���~���CN��|dB.ʫ|C�`A�AJԒq(X�Ɠة3\���J�騕1�E�b�>�3�O�׽{�.�'�c�v���i_I����>bn1e~�\�����8.�G�A���.^�h��k��w����O�:�O�����<&iaj�cg��įP
X�!X�L��>X��4���}�>�����q��+W�%��駟�#~�dg <���~��pr������Ν��`f6�ɽ{��.�ט��q��Ֆ�6(\�F�-�BK�Տ�m��HBL��y�����͠�p��g�W����s+��1�O�7�ܵ��H�eI�����*����-[�S3Ғܜ�/�g�o�똼�bl�<̊�����gg����Y�%��G�6YZ�̪�!t9��GO '�Ș�0�;�o�b �d=bwj}(����$(�I��*z�ΦLyr�����HĴw�(���=���O8��#�h�~V��T���S��?�c�d~6�`�3�\���X�Cm�<���7=9�A�5�aeeY@���5 ���ɝ�{:��6�V/�X؁ 充�W�����$�� ��hM���/T��Q�T�����3��K$-��n�<����J�R�i�-r䅔�l"�a3�\"K�����d�4�(2Y2?i �9qnfͧ�F7�Cz��Zr2��l?�*��Ԓ�)bL;�d.[��ZY�z� �䷃������}R%�l𨜜O'qr�(;��L�&�ʲ�g:]/�p�	@����5y�ܱ񣯁����>~�	�V�W[�m[�Du����/9��a&'�i���h���b�;آ%yz�%��!�&�B�p�$�Q�(�k wZ�|�7j�������^K�T��&M�t�FL�/*:uJH`�e&�������c���%%4J $���ShQ۞��g�J�����򲀒$�3�l��(۞����Ɇg̻��
a�C���G��cRo��cgg%F�%�Z-H~����G�P
�W��#��[7���lD咤�v;�B1�!��oh��и��w�v�|��u��n�X��]��Z_{���#o�=�8z�����WW�pl��o��Nc�J��nzZ<O�q 0( �����H�J�������o��*l��c�ho6l�`=�T���S s�/�^�\����Z�.`�$��R��������!������:3vL��
.���c�J4�Kާ6�6׌#��T����[�A��L��a�ӄ�\#�6a|7N}M:��>2y��^���9��iqn�!{������p��3D���!%ݬp&ʶ<3�?�8�kŷ��3k��Ya�1�L�Ȏ�����p'r'�q�h}����iXd��Lo��:sf|�����D��8'h�����aJ\�����G?���QhD�x�l$f4�Je(2
��G�UgL���`=lx��}SǱ U8'K��5������Ǐ����a�C�8&���T9$A,��Έ�u��qM��NSp-���"��ie3�@��K�RJ�b>ą�j�3O%-�V�'"X���M ��ܪ"7W�hr��$ˤq�qoV39�n����"�H��M+��O4=���K�q�ay�����|�4ck�@>�@,�ȥC��~�'�A�lR�-bM�Yr�X��q���*ȯ����\��� �T�f>PjӍ�f�r2�K^�v�ۧ�3�[�ZV�>M�}�� bf*�Q���n��q��s����,�S����@�[~��a�j�OZq���X���3c�J�GFz��Z�h�����1����c@c	wJ٢��.�5S���Q�PƝ{���Q�4�ޖg��
0�f}�������)�P��m�y^>9��0pE�G�Y�K������FIes�pE��Z���� �1J�����q����9X����Q=]UI�V(b�$S
��́TR�V*m�o1@����5`t�����������_l6���/��cǎ�Ґ� L4�^���_ �a=��N���FFGK�"������p^{�5@�����K�p�_|�a"�#�t��5���1G��w��\�芖?  @{mHxjw_B�&ZZ��/_�:WWW=����XZZ�Tr�-�Js.�M��B�^��E�A�ͷ�����nO�	������+��AC��{�-P����g���$��z�(��2�|��%���1��d��|�nZ� {I�*&��� ���vݢ��d|��yv����R�������,l����ב^B뽮$��qԝأG1�VO슦ƏL�5L�ĸ�Ncl��Ny�&��ZYlʰ�i6{8m���vfk?q��9�"3F��'B@EKK�ą{d�R�=z�T�[ۍ닸Iq�j8d�R?z����������M��I�[ۻ���k�6�Ϝ=����@����^�;�p���c������߾�; �#'����6���W>���[�Sӷ��TJ�ӧNPܿ��w��/^~w�Ua%`!6K��XYYL�C!�W�˜ǥ�'/����̑0L���L��h�k�G,;i¸�ߦ���ݓT9X#�NS�x��Z�d���Q�U�0�y����:$Wul|}cM�
��j��k��/LRpa�®�V��.�\/�c �#Ӭd,CO��*m��N/ 95Z�FI²�8�w�;���ĉku�AQ�"�O�J�+¶D\�8h�!p!���b�t�
v
A$q/��TO�Q$�]L�`��9��F��Rh{i��\�M8���!�M�O�&�y�����^k}�$
>�r�,Ş�*w���%%������8L�
!�ww��z�����o=�6�=X��@��Ҟ�k�g̮K�n�S,�h]LS��������85��P{78n��Ļ���Ipu!�^obr�byi�FՏ#K
U���c�q*Α�|�k�t�����'+�{���AKALMNu��vG���|�D`��G2���"��0���,�+��I%����E9҃�*\Q���I�3�֑T�fJ�s=
�hNUKz>�lI^A�*���J�����+���#�R�ӓ�yKDŚ-�=q℁�tK����ͽ݇w�A`�J�vg���D�l�<^����r�yҚb3]�i
���r�rz���|��@Vq��i���D)_��S���v�(�������ɍ_(6[�ȕ����H��j����_z���ؤ�<*����<R�z�f�P6I�nJ?mP��$aR����d�����CeK(\Ȗ��9���9���@	C����hKڢ�r٘��&	�irK/耏@��.��xG��QpD=��)�L�u��Z��Ki��8��e���[+zc��::~�@���' ��])-�P1U��e�6[���b>is�ş��_�S��a?sIz�o��l��F+�ju��"n����aWomo�w��`�(�կ����>�g�s���':���~(��9'�W�Wq���Ƕ׶k�+xA�[;QO��W0~q�-���Ry�6:������V� s�cc�Ϝ���T��k�ՒDo~q��7ސ�I���G``<\�37���?ƚ<x ��z �pwgΜ���o��pW�-o��:�z}lss��k�%h ��E�'󻄧4> �\|����!�P���t�{�S�O�Wk�J'��y�Z&	��;^I���k�p��qTX$��&��
�\�Mt����r"Sft�Q�
r/���Z �5܃F�<���%h�	�Da�C5D��� �
�WLU��<����&ol�tf�ו&IP�NLLȓ5�����lG�Д�O۬����DG[SIj��!�g�r�T$:Z��"�!�lM8��]�D1�� /HU^����a:�����0й&X�8{���<��Yf�F5L/���f*+جT���l����X�=j�@�89L�z��y&1��gfd����:yd�(�k	��ׅV����N���6�[�u�_���	ˠ���%��G��V�[����G�Fъ�Q�g�Md<���~ut�Ȇ ,b�#�����	2@b)��r��]eR�0��MSr�xBks�])T���M/�[�q֫�&ٳyY��ө�:Ps(�|�-�T6^qԚg����gԲ�ؖ>W�i������2mM.����O�V���	=p�w.��Ka�1�+���@c�H�1�#���j�x�0�;�h%;��eq�V���# -(�^�\{q�Τ#��������Z��'#Nhu~3��o���\
?Y?(o��.�Mk��r�]�l޽Q�j���KվJ"�0, ��&�p���y�4C����4�����G�l&͈� i�A�tZj��^r`O��T�^�;�6��9sF8%�܀���a��f''$��h�$CNLj6Yڥޫ�`���y��V�����g�:�踅v`(�a~�>}l�C�0��C�Eh.i�5F|'&�CȘ*7rNS/W=�w�Y�:�u����I皈l�&B�q��tf��k�,�?�05%	�O��~�]P>g���`���wd���G��+�k�X��]�G���վ���Ua4 X�n���vT�C�R�C��g�}��+����KXh��~�^8{�,�����0�_{��i<������)�)d>v��kk++X��W/��sǎ���~����1���~�+�t,;u
��G��W�G����t8�ܔ�q�2�	�DB��8���h�,h��|��	v��q!"2Kc;�wcUF�yi����eT������xq��2ӆ��D��&��%0^DMg���(�L|��͚��W��ܔWO��W�"9���.~���xhO��%���)��Ȍ�F���i��t�{L�a5u#�2�Ϩ0
;���Am���2�lҀf/LҴ$�.z�ݬ�������a�e�0�xJ���b	���\�\�ʥV�s���f�C4����.��d�2��gĚ����M��8v�o�ҋ/����M�Ӥ>f�=p ���1����Μ��8;�-ϝ� ↡F<���{�2�)m5<QT/��2VEi��ٰZ,�'��W�gV<��`�������)���7n\������@Ǹ.0���+DI�5mT.����-���,4i���
,��9�ɀ��%�>�C.c7+��FY�H!N��AXt�ǹ��<�����%�,���LzSI�����5}�*��=��]�����|��u��.,,��q�3 @%���M�M������]	ag񥸞̲�qXqI����N�Ν;%-�gJ��	�K��핋�F���O<$q�Z ��n��RB�hi1�
퉼~�¬�^�����e�����c(����<��|e�C�;�5'�6S�2# ��2�ƭ,��D�QZ
@������{M����Ű�iK�e�4:.���0��ƭ�x�[;�ݠG�.BO%K��\kc�vÉ=�ո�)]�]A�-��>tzS߯�}V�L��>Û�oԕFE�/^���%�$����쌯�| �n;-+%�6W:�%�W���aYptr�_"x���yn��`��r(����\[�x��1iO	+��k�O�"{j�W�Yr&�e�����J!����d>A�g�X{"đ��lu�d/�6z
ĥ�a�A,mQ@ՒĶ�%�0_N�<23?MI�f�Rڥ����E����GW��A3�_z����������tY9�x�r�&ވ�	R6���ݻ���1d���7o��ޒ������\ų�E���O�;�8=9����^�r�ŗ^~���/>�Z1��	�u�67�#���@X�n~��^~���O927::2Z--//C��5���n�^��ӓ�����2ޅ�x��;�P� 3<%(�W_}���O>�|����o��e��ӧ�2��)��s�����z�/���2�D���������������ʨU٤g [0CA먒4�@���%G�_�3'
��v�6I-��&R�k�6������ٰ/��5!�o�3�Jޅv诮�wW0'��M�f����0����"�b5^*��+��c�%����Z9L�@9E/�>O�k����������Ŵ �tT�I�'Pc�~�J�H���(�̤WH^|��a� � 
�]t�)���c����l[�\8��/4���a�%(������a���Ν�?�?�3���
�z���@d��y�7������ڨ�kJ�D����x�fx뭷~���qu�<ϑ�1��,k�qk���;q$І�PZ�S��˷���((��k���c)�p��-aJ��*��9Lq�%Y��<��N.ֶv�45{EE�1v���$��:�2�<ȁCӕ8_9%��N4DI>��B�%�"�p"x��o�Ӂ�
V�C�Y�b����,�dE<������T	 E��(A���1.-I�s��$��1���Bzy�r��a�=�츯s�7���if�3	#(�"%Q"iK�ӓlKڵ-U��*�����koy]�l�e?�+K���e��(1�$A" � `0�gnNݽ�9_w�� ؒ|5�s�o���wr�NY-&����h�Y:�a?R�R�KDc4@Y�̨3�X0��:����W�t��H�Ŋ�G�t霌8�J6]ẑ&��� bMG�Z�1��Zx�G���@�b��;"�28Aթ���
��<G�ق�ԁ]�:��J�NK�6�I������-[pG2�$'����j��\�V/�!�^x᭷�ڹs'����T�|6K�g�!�R�v���$��칛i;d^;��ƍ�g���C*��i"��� z���,�K
�nu6[�+��v� ����Q�c���������ਫ� cze���v�:���U"��w씙�����eM�F�+A�ݿ��o�d�����g- �Y�g�)�}�{�MUv,���Fϯg��>� Z���4NΉ�\���$���3�/�߿�D�g�����o}k����X'qe!�[[�qGlh�}����8�+in}aX���~Еd�<��<���m==�u�aX��o�Z�N�����i�X�����7^��%�8n�СCxO>�$��Sc�`�`���%3���xJ7&H!���a�t7
"����1�M9F���O�\2��֙��  7Q(%1!\�`<�s9���-b������Y����u��vW2n��^}��Y��f��!À�BpK�F��A����3��x-�yrP,3��p5��H�&���,�!��lk��-�3Y�ռnMg}����}�,�9U�f�����75�p�E3m�|I\�ޞ\� ����hk�t,�]��S*+��Y��a�R�,",X���J���y���n�
���^� ���nj��G�Y����޹�����σ'O�:�QQ�9{�,$,|c$�a�R���q�I=,{N�ǭ1ۅp!�<��@ʛ
�)��I������ܺ�p��a��lgΜ!����V �J�̸E0r9�$3��2*�L$�c}X!٘AC�kD�t@�mB!��$a��@HE:�s��?4�2Q��Li�%-Tr�F�F�����~�7 ������@��-�/��8��z��:H{�T�E�����I�=�	���Ɇ5�:�]�6c��$D�܋��-�{������Y���������BF*PK�%b����=� �2�bj�f�@,.f͂DUE�-�n��tc̀���YU+Ii��룚�s.\��SA�������x�(��_����R�M�#cdRq�a�B��3�ǌ�$cqμ��GH�L'R��K36L\%��qN,1���C�d2��O*ak��x#�4���I�zR��b��VQ��d$NPs���kB*�:��\&_r�&gǯ���|V=�1�Ӓ���c������1P��������ť�\1�]\�oo�����I;|�2��5Es�v5�d��0=�?zy���	?�Y,��d���2-�"y�V���N�� r��ŋ����Z��tR-�9�Z�"NH4&(W8u�>�b`9����_�`Ei�x1��}E uA��8�{$�����s�mئ���|���u�d��t	2��[��#��߈'��F$�A��ROē�yk,��T�����zG�l��QQ{d���f��\���S��5���tZJkp��V��D�dJ�B��֮�زi��5��&� �Ԇ�.v�Yu��;����A�=wf���6���l-\f���{��z�ȑ����zG�a��ޞ�uم�'N���V����M���V��^�����������t�2��U��44������[V[�����vd�3EC�������b&c�:`�$��س-E�&��|���36�Z7��ȉ�4#v��~ ��0�8��tZŭ9�D$�k�e��.)�텨aH%��O͸�Wc��>��\��N6�qc���Y�W��v^�Y��S�ƍ�H���~=A4]�ZP�B�z��'؟��K�!��\��O'��0TH��j���9ST{ѯ���a3\�]�tQ2%R"�H���+䮀.aKq.,΃�pji��rb������t8��Xl��Uʗ.]���{��G��.^�sCY�m�6Ɗϟ���K_�s�C�h��,Ü³��� l�o�í1�	2�fM���	�j��|�8���IaV��t�"me�z.\���6�op�*{<�ѽ��p	*-��޲A����4��3�iK�Z��kh�qפ�B�/t���P#h4�l;V4x��P����0�J��5(=����	tl`.A�e��&_���;0Ԋ_��K�O*��xo���(�o�f7/쎚P~	<V>11������������2㏑W�nZOMi�����fR�E�ğ��@x�t6 3�%�9�G��1$��8���#�8��N	�1�q��լ��w�Wd}$���X<i� �;�R&�i��%�@ߓ�)��B{:f0K
��g�X*aB\8Z�����s%���vVu�"/J�uTx�L캊k*3|fd�MC�ߥ������Pim-mXj���ܹs��.�}�k|�}N�r�d�����=BP����J��T���0p��rh�f	��?Y��l] ��_�����HBe���WäC.N�#~%<Ѷ�o#��f�ܦA#_	�)N-`2�	�t�y$QE�����PV���)�i��A�1C}4�]�`��%�5<̆d�'�x����9n;5<<,v|<�TK�?�O�+G�yrU,�U�)iC-�y���`|P��ɂڣ0��x?)
�a�����>ߺu+�2t;���
�DKn�ؑ;v쀙�H7�>v�#�8��c'�������=�쳳�3 ׶���^y_��qr���6l�ʔWs3VyE�g�U߳g��g?��s�=�kA����z�`��H���ѣ�)S��ա!������&�#N��k��W�I��g5[[S���3bQ�/G��D��䉘
8X�<?�/b_ZY�q�-��L�$Lԏ�
�T�f(�K��d@+��,�n����]}�F��P=y�)9X���Ϙh!�{a�@��A�%�VÖ�ry2Aq��`�6��S���XM��5Ċ�/�7�~u��=T��h+iFӽ�i�7�Ie�jh�q�%��h���tZ�@��Z�$(8�-褦D����F�Z�uy���X��s�l�����i�8v�̄2��ORX�n�v�����qx! q�V���i��d%�'b�g>���a�A���?s�l*����� X�/s�g�j:�Tw�&��LNN�d̊�bpH��p���o�A��4��n��R-�iӦdL�!��ZƔ�=w��х��_��_߼m����#���J%�Ձo��:k:�/�/$A>mC�i([�m
)�	 ���1�F �A��f�t����]���M_�u���_�y�E�M�󡖤�	���	�lnǥ!�+���lߎ�n>�U0�X�e<�xSKMh��
E��5�e
��D[�f�"4cG��a;}����5kԃ�.�+
�rMJ��v�� ��KC�ҞE�π�^,�e���z��h�2R���%2��%ђ����.�
K<𹅥rA�������Ĉ�sS�~��ؽ5�$U��
CM����B��Z0�7�ّ��TAd�Y����B��ĩ��LN]�ty��	p@gGGA!.B�c�)��5䵟~q��$�e�B����A�J���C��5���W`8j�˗��*e9la!;2B��Klq/�\v![�ʧ�C����A�
�tG+a�qNa�l���#�]�t샣ݽ]�\�9;���+%A�j���@��;�5�Ap�VMķ|�<@'p*d@C+��	{����2Y���.���aDD���T�Z#��eɉZ�h1�D:���եg� �S
�
B�VT8�iok�~��CPCE�FP	.��*�.�<{������o�l�v���gA���F�	��d�����j�ډ'e��=L��..f�M�ɏM� ̙2�.��sD�����YCÅh�R���Z�����̢80�����\�ģ��v�ܑhh�r�ܿ|��M	{w���]<u��C�zWu��_��}�n��cG����<p��]�.�b,���Ց�1==��:s�̱c�}�Qxw0��ɩS��w�@�~Æ��xJr �<6���k���N������a�utv[v�1�O�@4�B	��{��]�{�re,%�I�b�?�K}̭U]�!5�Zh�ٖ�d�\�f�+J��B�	�7<?9#\���r�b6���̽�Vj����(�*���H�s�>5��B3?H��9th�F搕�y��m�#̫�Ŵ�Aa�%��v��
�aܮ���$d��[o��$ex궊j��;:�a׮�8�<Im��&��pn�Jh���:���Y�ЯU��K�J�A[��H8
]H����� �t��[,�d�XV�9�9)W$����� ;)���KC����FK�@��"1�Ac���x�F�[�l��~�;߁�޼y�{������*�g�y�D�g�5�!��{�÷y���ȑ#���Y<U,��
���]�X`l�AwtJ�u��/°;a���9���7lذs�N�g���*���  } ����o�����޽{q��g��'����g����!��2Ȱo?9A����
z�B��b�j�#gF09le)$<OX���`g�_Cre���/D4�2庢��v/�.����śL�㵘�
�^,!l�Q?�h����ic�)[�>lx
������v,~|ސd�
KB���g��c� �dҜ�	:�z�*C#R�U�L+A1p�`k�j��.���[��~���Dߺux� �Ǔ1n��<��4k4[�q/�3���}#]���s�b��E��Y��ˁ8�x_,��x��~���đ�y��#Ց;��g8\kkQ�J�p�.�HsGG�5�KHɀ{g�Yb�ZgɸZA��ĺt�SF%k\� 	kbXgmj5^�X"�Qi~�[��1`RN�ł��/^����ɓ��%�sy���^P7�ݐ����6~�`����T�C�b�RsҘ$�Vn
�FCIZj$����lMYmMf`CB�����cZ㯈������H���"����`���3Y���G#���}p�̇�s�n�H�ض������j��u(��9�d����D#�hޡ��J��4�p'&���jY��g��w	���bӥjS;�YT R����/_�M�g�>蹿�������$w�m۶/~��"�P�"�X��Xn����٠�o��/�<?��ى�,,��<��@�Va�@w|����1����ԧ>������B[�o����@>`y�z�K<����C{R�2h��%�-4��[o�e�8D�tշ\�{<E)S��m׾�&��*K�6�&�e?(�5�er:�R��ۚ)�OUKZ�[,����̵e�&���܌��.F]���^w����
Y�^	���H}�ɸ1�����蟨�l�FYu�x`�p]�f�P��m*������K�l&/�1���7��-ϵ�\xl&��CL�I�$j�rW*VS�����&�Z��eq��%:��oQ �\�}�X\�h$)�ɔ�
xfSSK�ڵ�O�.�K�mQՑ��K%�䑡U�O�Ƈ0V@��tc���b>�u�R�b�p��E|���}<x���V�ŢׯO�)���lo߶eKfq靃o?��C�/�"��Ӯ��pqPf}����㩔}�8T.
��;���,�`�g]�Z������-w�u>����&�>�/}�K/��NE���E�wM�;#`���%��s�=�G����8�D�;�5��~ݜ�����J8(	G FM�	cK
��f���5���HN� o����_�R�w\ԏ�n�m,'��3j��N03��zE.���n3�uꄑ��]&��9�pyZm����ĺSk�Y���'+��Ȩ��r�������f�缘T�g�����ўH&d0C��U�&������V�:�d���4����9|��}��>p��5�z��)�����N�A�xz�Gg�Igּ�ݩd#dϠ�~�|���LslbB񊣓ׇ��2pa
��߸62�(9xC���,UR�K�\!�ϕ��bA
_�� Ru�$ӈ���م���ؑ` �`����-�{��
���J����>F�����~bJ�bnbF�}ëU�ؐjA�21����\����ݳjq)[�:`J�HTKf�Ŷ��p�q��,{�#1�څ�L,�h��b*�POvQ�ì�4��2���M�*�����N+���mi�(��LDF����n�J��.	��)�չ�����(X��s,�J��zժ�t���&��&�b2��E��[��{7��R��;Q�����B}�U�SS3�ώ��3��`�p j�����
E�σ�\
O?�#����%��q��RF�<d�d-*�u�1�������<W��]m���d[��'h������Ë�/
�}&�nH�ʳO��8l߳'���==]0n:��2�#��.]��{z�_�x�+���䋐�M����pV&�?���($P*#5����L�������r�a���O�kq�γ}�v�v���G�+
'�EgH�u�~;��]�v�x������cǏ��jjh\��1=���������u�{���������&4|�?��?{�8������X�N����{�ӳ����w��|�w�}��o�&�s��>��s?�����}���ruhz�:�U+��[�n)�p��;�y�܅M�6�[�Ξ93<<�j�*������7�^H�k�:5��ff6$���+�!����b�
��G�pjj����+TK8CEKQq	횒 *�\���XMk�A�BѽV��P%�C������� n.1�[��N ��S���[~H�f���k(�d�i�_�x�_t�r1�X"$�|�v�����rY��Y�^`�o>m��Oo���B�~ǁ�A�%;z1�������0��7�-�lZ��P�z}qv�lnmav�H*���0!�����56☦�t>�i�,'4%��s��u�����S��^��ǎ;{��$��ݷ�9{�,{�qE�-hٽ{����{�7hF�;�jy[f��g���cp?���s�έ�ׇ~�{�!/pN�:`9Wᦨ�a;�@��3gΰ���3Ǆ3t���Ν<��J�=f�.�������0��V��q!�<�i��
�`E�v��[��������¹�0� ��0��5n]���*%��cޒS~^��n��A*QL��^�A���I9|���D�AX���#�+��M��jkk��x��������$RR��XWcS�:�,��z/�,����q��<>���h���ш�Oq�e1_<j��2"��N��\X^{����4$���g�­4{�
��ѣ��?NQ΢I���K~kN�b�Ax�a|K��	R�YsX��"m�H0����I8�Y�5nԙ2��,若���߭���Y�
�Fↄ��x�eF'���J��()cuժ�vm,���#_ᚇ6u��E��+� .��C�A�IHc~N;y#2��q@u�L�M_�ʀ�V�y��t�;A�7�MAk�nC�$�D\r�,h���X�\OȤf�9޵kW{W����/b�x�ssS��R�d����O|�g���σ�8�@��x;��#��/+j1�cj���`&g��,8#���O?���Q��\|}UwYo||����������X�vh�G�=vرc� �K�/ 9<y�F�H��7~6<<������~����A2C��K	Mc+�x2lép����_��z���]~�����㸎4��$l�lm���%)M��]�;Z�q-����qj�9'�8N� �<�;؅��2��ҍ�L���/�b��:t�m�eRvFf�-%Y�	 pѶ]��j���m��}�͈-}EQ+�8���F�j��{;�~gָ�o33n�h"��S���7o<3�u��OF]�5�m�e��Q�CS�8�Ta�1Uf���#�ϸ����!��gwHS��3�M�Ac���Q�ks�a$�
���KF�E"���M�ù�f�����B�(�W�����N$˗����]�(�/-�G��irp$ҦX!��N�8R��x~�k����|���/���-�:���������>r�9喫��J�>�ē�9�%�������\�|%K��|O�����/��/
���5�/��.Id��k��'�Hp�paq��C�LW�����w�u�1�]��b����6�%G����k?��M|v�M��j6��v�jh1Xxx>l6�e>��(���I��YHHn��R�y5��R/��*�zL�WY_e�~�%T�Y4�B	�o�)��r2�<���"���n�=w�#-� Kc+ 1Q�V���� 2&��E�z��N	.�:�r$�of̏�9N�-@��&R�<|-u��%�P�(VVD� ���Z\3��$k^�n�f���n�ZU�Z�����%+�(bO˪2cE�a�N&��%KJ���M��l�R��hW��0�:��\�)%D�i����jHc�ׯgrY� ;v#Zidz�/� �j������K�[��u,��:�R�X��AG���2�+��*�0=v�],�n�\�G���V�Q'��%��i�Y�\��V�"��#Ru��nH!+b��%md��6�HZr�`|���8��s��6-�"]���'���r��s
l;���1�񳫻g�֭�-Kp�k����&���ޅEB�PL��#vLʎ�����Ĵ�-EO`��-���i-�����>�y ��H����*��1=�TP���Ai��K�(�=]�o{k�[�}���Źٵ�֨�/z��CS�@q�=��tw����/���~�Ɓ��pB1���\�>�,d5�����!�Ϟ;#=jh�ONtttt�W���r�4Y���:ׯ_�S���X����7a�QN?�p���.,,�4��v�X;��V,�>}ghoi=v�H"�6�h����]�֮~�������J�_ezU���>�����Ua���2<<��pQ�����ܯ��z����W~�W!����={���'۸q�ة����>lbQsbxt�b�P�T��7/���#���Jezv�ڵя~�������?������krr�ֹ!`Z��
���>FN��L�gl�0%�49�긅r��F��d��4j;����!���
@�=ы�-M���5Tz��͂|��L-�T�hE� �b�NC
l@E�
K�S7��[�gw���"�!J�}Y"xR��n[��-B-�g��e�i`w�_Ϥ�]*�1D���"ˌ�4a����Tsè�� ���(�-��Q��6����a���C:�mI�C�����51>~��A�L���Z�@�1���#�0i�m۶��z�ԩSCCCX �*v��?������w���/H\�dI~�ӟ~����g��Ç���ݸi�L���7&�:\"�8�r�U��
N�"\�ï������(0�6�f<,�������&���ͮ+�N����k_��9t���d�N{;;09��� ����5PJ�Q͠z�v{Aj&��¿�A�2$T����a��`�e>xP�EY�A���;!4�B�^:�zޭ����}��ȸU�A�B�Q�RtB�e�|�z�6���'U54��<A f�Z����a��Y�v�5J���E���?-���P|�3�<�"�ϗ��$˘\��(�
���jD��%.��&��yjaj�Ät��`�J#�sC�5�����!4��8����`4�UMF{�%��1��5���B`?���Z.�6^�k�,� .#vr�+QL�����;���6T8N®LF@͠��R�	A��T��T�a:/�A&��r8�ؘ�fƐ��St���Wx57r�me<�?h�}c�M�059E����l�D�`-Eܚ��ˤ��`---E�3
�WZ������G��0��
퍺nͨ�/z�\?�-�ؼ4�h�u�#0���t��ݻ���ǯ���{##ý����ZX��5�X'<��wO��@�a;JZ-�����}�vW��?���9v��/��߿Ǭ[�^��������؏��sh"��}A���-V���&P�N/>Yݻ�bQ~Mቕ��2�l�/_9q������Ğ3\J�Ґ�ɠz�xG����zW���{�QWO�̉�����ua⾸/=���������_��W}�Q���ѣR*jy_�����[�S:�dN_߀��k
�9	m�ۇ�������h"1���a���"6����u�ʸBcر��C�Y�RE��@T�V�T&5�O�^�L?$A���Ìc��n-�Ί$d�Z�W��,7t�	�dg����!���gc�����Y����l��Puw�1w���25�+�ʔ�f]�Q�`	�3�˱�t�C]�f�9�!��Oeaax�9
����a��>��h���8/��:�h�R�T�'�Q/�nnjjihL'!{�jo���ެ^��^XUB���A�Ʋ��V��===�e�f����
9lsKK�������L����ׯO���kժ���)�dx��ƍ�Aa�@[�mh�o����g����?�����˯����x������a��G���+P��=|���W\��y�3��p����-H�5t6�����������iX�O�_�x�#��r��	�7�=x��#�?�9�˗/�㒍�#��;jNҁ�,���Y:�*�<E|�όU�q�L�P���WO��D�v��!WNEi�џ��l��2K���
4��8�5l#����al�E������I��Y2k�x�W��ċxB㽰e#�d��ZF��Mf��XTj>��<v������T4�'�Fww��lffzZ��m����I�T��5�ZթZ5Eif����\��/��&���L#S��U��3��S"��ut�����%�X����p��P�!1�`W�`��J�c�x4��._�Zbu	e56����p�����n��j�,��íI�ƲE��hߊo��V ��01�jn".�PAt�f�\��A����e��6�B�Zbu��1��5�!݀³�0�'�����J�N�����3m��%ڻ:K�G`�m�8l����Cl�f��Ş�:)��h��hXQ�]̟7|���{S>�{ٸukgwOvxXЙet�!3eJ��nl^\�,�qS/0N,��&�e��8s^��6{,p�j��n�D*�`������5c'�f����P�ҔPY�+�T"��yˆ�=�a;o���W^y�]�k�JvA��T2���<='h��vl�ᇜ��������t76]���]���{�
�)��Fl
�nqq���W��?���{���<w����M�O�>��r_��dJ� �::�t(��w��דN�"�5l1L�͛7�[�W�����Y��2�����Ç�;V�寏O�<q��!�vuo>�T.J�j>��p�\[�xbc������;~�����_�z��+ij��~�>8�X\�~�]w����f���%R�|n��-׮�����?��?��3O�+b����ؾ������̼��I���$��й�B"���ܚH5�����3=GRޞ���5�]�\��ANڟA���X�v3�Y�nl�.�b��!�NH,���|eS[+l-bjvtt�>}�'�v�jb�SEFT�{�'o����N��{nf%�O�Z��d�P^�JhE�qc��
�,�ռ�:��ݒ����롧US`��jl@�ޭ��2��	���P��8X�S��򱲌 ~�,�U���O�M%^�cX,`�12�β��@��I=M,%���6v�A*�O"qd��-�g�)8���__��_�����o�t�v���˸��	�w��M6{���X� Khc�z�8�����!�mtlgزe�ځ�g�}��๳g����冇�A[f0s�l�1����vy$��b�t988855�{ܹs'��	��-��a`�������s�NO��U�ݵk'�N�ǵ}�Vl.$�t�OͲ�B��E@~/[��!�/Fn��֘Qg�����+5+�w�t�}Ǎ0��(;Z��Q���#�W;`r��;�>�Ϫ��9�6kL��k�q�_R
î���a�	[�m����[���{|�c 
�׳Ӌ����.Yμ�5���"�c�F�	����0w/qׇ'аY#A��0$�h�%�Xq�6�0��7[-U�4����甄AR��1g��Ve�m3�'���D7Q���"^��b|{b����2=?L��[3�9�3���!!4+B�)&��ٌ����3��M]U�Z��Y�À�*8?�Ф�}&�Ѿ(v��)�ްf��Ͳ3�m�D�R#F��r��׊p��hԻc����[ s�\�ƍ�j�5�k��hjJ1X�419f(?���${Alm߃x����$Y�yʮy�kH ���o�����_�T�;�y�s�9?7�7��k��>��S����9�k�N�U*��N&�9�A�￯���ԇgO�:�́�'� !e�V���>��8����?=2z<��o�w�w���������b� 9�kc
�"Ŀo�>O����1�s�X���T�� �o�@U�~s���K��@'[�nUd��2��t����M�uJ��m�n��ѱ	����k������QF=R�G	b���e���~�����|�+p��agg��v����-��%"}Eg2�A���ի���$RW�\�����>>
j�hΜ� ��թ�VY]̊@���  ��IDAT��?_nAC�u��`��Ã�m�p�8��r����٬�N��2=(�ن2�^;��҇7Fg�3[��u����pX��Fu#n�l��O�>|ݺ?�f�ȼU�ڍ�2ͺ2m�t]��R��JWys��b�[��c=~���[Z��!�jL��Z&��*���)�s�����,wbG�3N��j,D~�8�����7INP��jI�G��F^Z�������"Ѹ���^�ti����������:>��{`�m�׮]�@�'O��[�s��F�^�V}����F��^�<�q�T����A��d]��۴	�_���d�{:f�0Ox<]]��N+�Ⱥ`!v�`1�.���v!	9��B|ppu>#�:��)y�n�rMqLs�7gcnn歷��0пc׮��{�һ��6.�X.Uq6&#�lE�V�"�x���� ^�(�^]�t���Ѭ����o�t�0� 5���)u�\���j��?��@Ó3�Es$�ޑD��w��;�VX��i*"�;v"��Y��ʭ��d��I�|iP
C��:�Q�������?.�5O�����'S�Ϛ9�i2+���c;�'	<�J7��҉�z����E��bĶ3D��?����}nŷڣ�]�銚�HD���d4C,�jtŜ���ęS��	�~��v`����U���' �*��e�pFXNN���HDcQˮfH $�n�6��V�*?���5�U	+lpL�XjH�P4!`f�s� �xB�\��1S��]Sk��0�ţ�t���_KF5�<_�q�ޔʅJ�Ԑ�:�dBʥ���V���J�:�>G�j�x����Ar�B��*���$5Yl�O�4����YELv��0VE�T���s���0�P���ڒ���uYn����!�hǐ0XH��,1۟�$�E����xmZy�έ7�>q����e�m�PbKs;���ڦ����;�C�^�|�S�)YѶ��k##��-[��y�:����ֿ�����nX�ti���������c��O�$c�#Y(Ɔ>���iAzC\s��-d�`Ӭ�)4���0��M���R�p�����~p�9�4x�d��-� ���b^�����V�
p���`���|d3������Cڜv�Qg-���L/X�~�����=��C��`���W~g��ݹ��q}A�|��3�L�b�"6,�LgW�m���=,H�j~n� C�m�x\�Gl� 6
�[d��jy��u�_��҆�:8 �k�1�� Sq���X-ݦ|�I�,�*�����y��l(�g�Va�zh���U�X��݁5�,&�:n��?���$�JU�o[��<=bc޶?����*
��G�i�bp�l�ӱ6a�iy��^a�ݬ���<��^ן�C����D}�#,�6�>$�Bx�[��;������V�<��b��.�'k֬u=������O~r��͗.^ ��Ⅾ�wq0�Cgpp�u�4L�@�T:s���ȕ��|��6��g�y���_7�f�+������"�����x��Z�e�A�D�EVt�[���S�(nY�S�v��m�<|G\Q�n�=�s97o����R��_��'�DX	3�R�H�l��p*��y��8Hw72�t?����~0�t5��,�v�旋�c��f DbTT|4�e��Ɛ����
��xak��l�D��-��Yu����B˓�8?�vS��/�'T��N|�1å̒����zE+l���nh��< 3�hlq�����3g��ȥ�`��u��ݱ#���s�j�ЌCCCJ��j���/���{�t[cf0PE��!O�ƮZ�b�0��HL�xL�m��Z���)�~v���Nj�A��,�iX����HJ�=w�Yڎ"�0���F��������tF�Y��:�̉>Hq����}ݺ�&���Aj���%���1�	ы,�L(�Agh�y�|�H�s?��:�f����)�xZY�e0M�A5��S��Tm�����:��ms w�X3�H�2��I0�걫�ݔ�TPɷ�B�>�GX�"�C�sTЙd��w��0QCC�0�6�H�I%���Af�6Ln@sA���f:��m�dOD嵫WϞ=;22��҄�4��4-5/��ۻZ�m�|������hL���g�KŔt���L����P;u�����߮Z�C��z~��~��_<r�N��UFǖ�̙�B�7n�I��m``��
г��wv�9\�m����ً.A�qǛ���/��'/�(�j�2bZ(@��E"��ܚVN[&��B=��I������җ��i����=�c�����)�?�e������c[�V._��{|��Gpι�Ű��)ݪ�l�*q���Ң4��4m��5İz���^x��|}rT��|�?��/���e�oZ�2x>�G�
�KG��(d)'�HvO��c\����N͋y=/u��x\y�2)=����N@|�_��=[�[�E渢�~`�+�t������dg�.�?���3)QU��e��2fH�J!?bv��T`㺞�d�
�Q(��j�67?��fm-�_�.�uH�<�5�J,.��bغǕJ	'�A Z6���K��M���_��J.��d"�_)uu��f%�*GZ�D�(;�d:��P+V̚���j-���E�rz{%�^��k�X2Vu���-��v�FRcצc��H�Z%�Z������ޮ�驩�'ONL�}�Omܲ�݃o]�z��pMXc���R��)�}�ݹ\���䳹�b�)٘��vl�<�~m?���W^���ڵ������+)�y�1��?�Գ�����+�|����W�^��ĩf�Ҝ��co޺���Ψ�7n��$<+b�3����6;.y����H,���ON]HJ�C$zu�j�W�v�vau�|�0��� >2y�Ż�gVV/����&�A�p����� :}��k��^)����3�p��Q9�H�XP�Ț�x�[*J!�e�TB0����i�T �k�V��J�2��٨r�כ*�T��=�pQ,jj�Ӈ)6��+r��p[E�ML�*e�V��"�u�F�H"�X���H���2ѐ��m�¥vĔ��|N3�֌�����|CU��{^�v�=[
Q<���A��W��[�'b�s�����.fw�T(��Kk�<�J��J�#��:e[p0$\��ƇY�$��e+T����p�R���GaB��[[�m��P�4Ҙne�ɩ�,��L���\MT��������8]��T�Am8A[�P�����)6��ꠥ��Nܯ�fN"٘��Q��Ӕ�'�#�ꢰ�H�q��Y-VK�I���Y���b$�J&���R1�ℜ��y���#�(�WK$a�ȰZ�E��՜j�+��,.&��5��7�$�W� �����"`״��$d��h� ن��l.�bLkvv���cծFD�.ŷ�Eg�Tu��3+U{�Gԡ�l�A/f>�-�jw6
��Ș̘���ӡ���2�쉴�Km��FD��t��'LU;���%=ݛ,9��8gˑ�v@;2E �j�}&���|oϚ�u���MMσ���cJ'��rپի̈X���5��p�|�b��VD��nՙ_�%��R�╫xDm�=��@���
^GR9Z�^��9��U)�Z���ݷ���G��i�N/B��`CD��=;v�f���kxbM�t�h���+�v$;��NFa���s����O^z5����J�aŶ`g/_<{�]w��J�v�ҟ�?�g[W��1��ͯ^�eE�3�N�����@?���N��G�G��'�b�}���ؼ��p���-�w�؉���K�=t钩h22��4'����R��M����O��/�[C<�8?;5y�yCҚ�X,��\X�F�R�\��in��X�$L� �ӠI|k���tt�ڝ��au���#¤�9[(��TI7�R6G���o��fߺu������`>A�㯾����}k�%�1+c0:[:R����RSC¶����v4�f��%��TӨgԲ��o�xr|buo��B0�4��f��3�2�S*�56lJ:rI��`��d̲����g�Kp�bv$Z,�)|4�Z�e* �ێ��h��Gl���i���.p_��O�1�.'�=�N�x���[�S<Uxd8��9j���b�L&=/�T��V-&f��>?�n���U��:=?�$�A?��������j���!A��x",es��>��^{�OI@	�85a%��� ���>����ً�<�tS��˗�ֿ�����`��s-+�5��)�Q'�<�쳝����~���������'���-zqx����F\�7<<��݉?--̃�~�m�,����ʜ�NH���74��}y�W>��� ����y�	,$F�s���]u}fw�n���7��<�������)��L���W[�t��[�.���SO=��[�l�����Cf8p� ��瞃�����Sݿ�曏~������������n,lǎ������FOW@��NQ�?�)�pJ�z�İ�ˁ�e܈[:�*�M3�7t�\|�s���q/���m�%��b
�"��1�Bn��of�_�e��h���%7łɭ,�#�yX�����*Iu���cN�u���
L��uN�)II̦��d�A��-�<y��2��$����`$��^�+&�hG���u�ks#�ŸuLw;::��X�Io\je�%�OJ��m�jo���:>ol��gM1$=�%@��h�Ғ�VY�g�[Ϛ9<ϖt��OL���vutVt�;�Y*:��� �0�jG15�C�i߮T��$E�Pf�i�9̳'�8a�xf�w} p!�|`:`��g� Ĳ:�X�'�1z�h��� ����{xh���LJ}���
^ڂ��uuِ�SXcק,m�p� f6`WA�@���bA
�xY��j1��Z|b������ږ��2��	��=�ec/�!��c�:N�*f��p�-����e���РL/U��L7�/^�:��۾};�J�0�AS~1E� w@�K�m`��H�����>�ζv,�3g:9b۳g�{���?�ӯ�گ����ȳgϚ�����'&��+��ShC������ߦ�ƞ5k�	�����߀޹uG��L�ǯ=������ُke�@iT*�ϰ/�>��/����W�����蕖�wp���n�����'O�w/D�;��F�3?|����� �1��A���q\�����q��Jw�|��3��
7ɘ�o-����	�"�=��NEh}y�W��frtl�����_�tS#�K��_ق��u٪ O{?� v���A�����̐��  3<�a��m�KdX���e�IJ���c*�9嬡����hc�Ґ�d'|��#��6����3����
,ESzff�N�c���X0��P�@Լ�Ne����#�n��%;bVk��q�"|{v��O�D�d@O���_?q����Uk�'�*x�m��=0��>���G�^�"� k�v�{eZ�š�`]|�������'�mބ596�eLO]�f��������￯gͺ�����c�#Ґz�cO��L+e�	�0z"��9a�J����0��̩��"�e���0׀'�|䥗^:s�^�R���g��زu����k���m۶�߿l�g������\� ��YRB%��be��n��.B ��8^{a*&�X�Tu���_�(vsP{$5�@8��;�uh��me�!kp�g�*��a3kf~�m����M���X7d>�)�%Þ����6gB`0�Gmh�%Q̠Z�_���rUxV9�)[����A���;�C��$����L�)lkyU.HD8�͝�����`��
F5H�Q�Z6"��J[[�*�����M���l&; #��eQ/l��I�g8Ae^V�S�C��r�-(�c�
%dI��q�5��|�^P f��̩n߶���KJŝj"�����~��_���L���>cƄ6��gMx�NM_0�C�9|8T\��M��ǥ��~I�ƍ��.^�z�V�;���9�(��X�X:LZ
ϧ��M��4��a��VZ=��'-i,	T
�/T$�]��zZ���	Of2��:JHL�X\됴���r��Դ�W��i�t�(�#0=	��rp<)g �:�!%���	a&3���nn\����)5>5q���v�ĵ�c�{�P�c;�ۼ����h
���b1Hl��M�y�W�
`U�;w�V��5/sj�?}�?��W�z�����,��!� ��ΩW^�Ì�TI'bF[ҍ�S�Gl�Z��DTj"�17=�y�f��H*aT�?�����?����۶e2�\fUoowO'�C�8q>e[�$7\USf�����-�������ck��T���� 9�G#LP��p���}�d�l�4rm���߸a+TTڔfmG#d<I��b������z>�F�2��;=)��h��P�@��u�Mὄ���qR��	(i.[5|�r9%�#ޔ�Zj�
�`w4փ]��7VX�Z�`"I�2>�"�܈2�2�
�ˠZ�7�n]���7^ƻ}�	����@v�;�36��.�B������;4���^��&�_�D ";����;�L�5��Ul.�1z���6l�$�a�ʸ:g-��:����u�*�L�� A�Y9~���a˖�����i( NO���c�NX0����t���{���+:荦*L���k�{W��qkԭ��"H��ɋ��_��G4�5��--?��O�z�S{���I�4��u&e��8"l�"�:V���t��ڂ�^�xgH�|��y+yy�:twv�r�U8R	o��~X8�$�ر�G�!l/f�u�����}���q�,���U�,-k#`�@��I!ӎ��!����a3'lϓ�Kc-�?��co�����pS��Ǎ@�*x��POe� ���>���
�<(S"�e�V��K��I=�
���UGbʔ�!e��R�YJ1���dx��C)�`�|�}L4j%JDCnڇM8�ꆥ����d"x�*2�L�%ج����얭�}���z����c��Q�o�椌ϮI�4���"�3׉)�,Zu$6[��M�\.W+Z�W�X�0}6���%� 	���30�d��drL�I0�&�G1�����5'��X�ŇlP�����l��΍$Z �� c��
n�|א+����YRY(��="�)�Bs�S��[�1D�b$�p���d����U��W��������(�a��['��t�"sH�+� %i���\ɾ�������pBBl���	�^�f0$���)6��ei���k��;�o�f����?�l��·��������X��i׎��e����8��9�bG?N=|x���Sf׮]X�+����_���~�0���y�[G�r�,�r̶�� ��c�x�K������7��M�AOW'13�L]jaC�rT�<��=����G��ٳ+���g�Y��t1��~,~�cp0ˋ/�����8	e��Ç_{����W�1kfjJ�������+K�HÂ>������+9�
�43=�T)ef9���&���3m�u��Ay��kHT5�A+�RB��}R���P<E���h\)־���7K�ͺd�� ������8�З�&��} ��W���u���ڍQ�ܛ"jn]�M�]���o�Y���I�҃��~]޼)���d]�����|5�΅�K(��G�����ėk>*����Qҧ�'`$���x��1--m�����X��>���8�]:p���5�.\x�7��j�p���HL¤�/_�zd�`&���`Io��&̗�ٙ���]]�H��ܹ.QS����l��t�޻q0y5M�s��Ɩ���q��@��dｂ�6<:ko��� P`����vtu�^qu��������%X��aVc##�(�x�ţ�-M���?��ذ��ᇐ8�����;611��Z�z5n�#$��|��U�M-͛�n9��	<v!�?�qڴ��Ҩ���54��"v=�iz���Wf���UXc,?�G�����Kƺxp�S�u(8V�`2�����1�rV�cGl����Ebv�T�D�t���lZ��|��7/L�ʩ��*(���qfَ�L&ʎK;�wmj���q�!�YW�J-�X5�u��������ڰ_�kkG;l���Y��H�m���Z!{^�D�>b$�XH��Hƈ��j���4�U��H!̋�x��q�JK�D�g�J
�3/7�HA�V+��-��4�QK�b��
��;��$�h�p�(#�\��W���Uw;�;e٬�W@�����@3�A��SըU�u?�J�����0t�7��h��,��%r �7��b9��L8�X!�0�ސ����xu�I�AtϞ=�w��f��;�������Y�oijdg���N�P*���������䱨	���ם�����9ݨ&I{!q��et��eH��Ϝ&q+�C��ғ� GlT�T���7eT�q֫DtFp2����{�jKS3kI7� �K�)f�]�-,�)���k�r�/�׮�&����\ύF;j�]�<��'��ѡ��Ђ��Ld��r�*~n��3!�j����L�+v��崾��dj
ڸ��?x��;z����>�я���BN�_;��� �׮�>>��S�tk���&�q�;�j�brUoW5�4>>����!�=���۞S��T�ZY?пz�*P(�8�����hȐ��V�a�k��laxd�;��-;v���̹sW�\���af�/�9�ů��]8^~� H��'��9z|Ƕ�gϜ�[�vrl����x�M�w���Z�Az���2wҞ�i/47��Ca��4,3��;�"��Ψ����\6L�è2��Ε��K>�Z��)���~W"w�
Q�`
H-��H�
����������<b�ĕ���,�;W7]��3�F��z���J�p�(�ݰ��B�.쨧�
M���e�i����=�1>������%\iOДD�=�?��b�m�1�r$ve�p���Nv��u6JsC4;3�Q��ɳgϦR��{�g���ؿ���� D5��ᗀ�����N�]�F�'��׾���w��B#����B+�@p@7mؠ�9��)�!���'N������?�����l�Q���S�38?�<N���:�jPZEp��p�ؠ������{���X)�P�gx�3�ؑ0L��x����C�aa�S��0�𭾾�=:!����R�;�v�И@!�m&�۝�2��u�(���qZ(Y�q"𵚟�����{y��'!jaY�%�C�|��HW�
�z6?Ϟv�i�h�����_>}�M���t�"ݯ�|�� +�7�z2<[q�i�	6�Zc���>�!�&R�3�&�[�R�_����2PlϪ5��R6��6641$zK0a��G�bKe���D?�Ă�e���D���ɳ*��*��6�dUsH�իW�K`k׮U���m��J>�FV��`*�d׻�<5�?J[����� ă�B��-�IwO'�~��i؝O=�5ɧ�8�Nݦ��/.勔Tth1��>ߓaKe_�%��r�Gw�ojx���e���8�Bw�`$w��
/�	,K�b\�%�>g��F�D?��)���$�}����+�x�?�`��'SS�P�4�å�Aq@���P�X�Ց�`I�-]r"x�f0��Kk�4�@(A�⛁|���qL���I�����:t�PX�(�*5EMk�}�GV�����d��M�0�����kU.\V|�nm��}����^��-ż3��`�}}} ���Q���^y�XXhX�g>�(�o}�[/�����ɱ����I��G�Bg�
��d�$�r�С��9s�:BR�G��a4N7�.���x�T���@۱�	\��>�H���|�M<���v�V(YA#O(�S>u5�uq;U�"��ݢ��]ټy3n�6�A��fg�3�&bvl5�%� �[�����~|L�4�:~�b(��K�FU�DK�� X�I��p��bv�'��eIW� }�+�}�`C	����(���(��V(�ÿ�o8�IG�Y��9"B 
"���Ϥ���������`��g��A�֜dJ�{�
Kg� 8[����5�::d��7��Xt<�Ќ�mic��P^�F�B�Կ��~�V�q����q�Č7�¢�0��g���.�gu�m���̌[���m;wf>��4nj��-��η�7��eՑJ�������y&P4׳�O��O����蝻`9�r2ޘ+#�ٜn(泣��Z[���=�HV��S�;z�'/�ȌF?��SS,�����]�.m۱mm��_|FdKKs[[+l���\:,�����$80�#�j��@@���x����_�B3����t�x�=�XbC:͂0�����v?~"[�zG�<pO ��؅���*F|�����X������p5�����'��|ιF,��15�ޠL�v{��&`� z]���X_����wy~�\����v/.���Q�vkE�_��E�W�6�{)izW4��iQ��4����A�*�<M�Q<łɆT��e'�7����҉���ܵS]Z��3�E��񩅹Y�h�%!X+�l͘�J�ż�אhYhġ����ex��u���e�~t4&]�ܻ
�[&�g�o|t����^��V�E�ۭJ7V<.�"b�X�%]>���f|��,#^T;����q�B���j�M[�㱤�M��5x�Jgg��Ց�C`Ϛ��5fE���8�V�� 2�vG�Q�%ئ��|�X��1�ǒ�2)Zc��f����M-�}��K�2q�2�ʄ'��8��i6T�2�An_(�T��n�!]�K��@�K��t�D>V8�ޭ�.�|YJ�^���/S�K��&gV9�FB��R4b�5|r#�!���ZW"i=a��t3�j� �^g�X�6�Ma؜٥Ր�f$M���3�\)_�O"J�c��O�G+\��h$�8?59�ZZ�\.����:��L�y�#�?��}U�
[K:r�d��Us󊟒� O���������~�����o�ݻwllD�HI�t�8�p��p1_H�����d.����m[�GF��o��7~�7�u���7�3�O���8y��O~��'�������À9y�$�
��Х���F(>�]we3KgϜ޽{��H��c˹L2@��G��zf��r�\VFb���]���G�ߺ��;�8:�7��7�[�Z5H�'-�]�7�pe�mK�<��|��=��v�ڦM��o=�����O862ܿy3��X"��A�`x
�H��*S�� m�d����i<�&�x�F�b�z��2aB	F�m��q2�!2N�P=�@r����U��B�6�T#�aaYޗ?4�� �u�����o��֔]?��&ȳQG*Cܛ�se�ٲ�wS���c���z�R5��a��1�-h�\�5�P��˭�ރ�Gm7��$Ih�3���\�.NSfՈW�/B��*>Ss{�x��m�S����S�W�W������Z����U/��3�D`T܅ �n�75I�>,�e��@0	w�څ_�'�^�R��;*%IJ���D,�Z`�8"8 _,I��ȸ`֤�����̢@�����Ė�w2����m�=�n,�ld
V;4t�ܹs�Y���Js��"D���(l���=J�s` ObF$����O���w:$0��s��U����n}�'Μ9�L?U&�����X`��|H)�(��)$�q�j�2 '�*KW�:S�Sc��!��of ��0e1� A����s�=��f �ŀ�R�OW���l)M��G��J��
��n8�۪�@2w���A�癑gi�=Lh�?А"�0�����\A
�8�kfVP1��'�2��vaLG�0I����K�p�۷��F�.^�'��XR�K���짛TU�,ξ�>�:�$hittt%P�VT��%|�T�R��i�ð�;�;�q��T�JHl"+��=��;h�q��*h�?��8�{�=s+Y�*u����$T��J`�������,WK��L���(IN�Q� f�Q^�$S��a�PX8�����\r��ET��;t�C1Ȑ ���=�-�snPyS/E��җW�Љ���A�׋o�Z��J��;����:�铄������LG�P4��H�ox�B9���&x,�8����^S��NaI�k�f��pP������T.�*yq�tDJKo�ğ�Ŧts.��HSɖA�R����#|��'�ğ����?��sP���1����8������1����~w��O�{F�q�炕:��3�A� ��E1(�
w�kɖve�s�?��{����>������=�ݵt���d%R$E�	"9f L��ӹ�j��}�j ���mS�LOw�W����6%�)E���!i�:���7��[/��
v ����z�#X�̤$�!��,�J?`����N%J)��Y�'1�Q���_������>|�رk7���hA�A���_X���%��XF�����07��Ae�[�v;s�d��$���!�م�8�7o���;:;��/�:&p�	R���Gӳyv${�M�N���0��3u}Q���;�\�4�5�'���lY�Do�������-�E�}r�D�g��d��mD}r�9d�r._Acg뿌Z���;8�~�R8F��=�0��7GFF풐vBu>h��p)݈*B<<���i)��mM�teҡo9v���\��
�6�}����8w3\���n#0���cY��c:�,�w]����w�blJhji��Ob��P���<X-U~��uwtJr!�a�*8�_
	�����cU����C��@�<���{l����H�ި�3�S#�Ovww1����Z^ڴyC:�<y�N>ӫ�����w���>8�R�Ŝ��kC��xF"X�3}z]���3��6�J$*�R�f؎$m���}=ݛv>y��q�_8�]�v�f^�u��ڦ���������s��1���\�~^Y����n0m���o�q�֭�~�#���g~����p�ɉ'��a��YO� �o5A{��K�)�s�&��U85�7�C���;;�����š�2���MP��@-Q?�ϲ�Z<{�<G�}����o���I��F]bΎY��˵jw�{`����9�֑�o0���&Ӓ�[��ke���߃�}���P#�@E�$�pG�8�������ya�XFÏI殻��- 2�6��UM�L^�h��0:r��Z�ܼy������ql�ͱ��
�gV+f��?[�=�Z��,�@��.@K�����8ǥ����²���F6��?��Zf��R� �����G_���Ç�=yF�~Wj����Hǳ�\iU��ҞLJ}��+�$��y5�K
Z��7-	3:1i0��Tq��i�T�wh#*�P�4�׭��U���A|0��7m�!����5Tizu�l�7��!x� i�TUꪈ�J�
����B8����l5�%R�J$��T6����71ی	�ē�]�S	�F�(�vF�Ԭ�BJ_E���K���V6c�ë�WpG����뱺MCDTH��L�2�N����a% �f���ކ��o�]5o#t1m#�T����YC)�`^0NWpF���cA(
�ĩS�ac�⬜��x�d��f����E�X�9E񥕼�4O����:Q��M������ϷY4Z՚}L-;�`�+�A��c��Ʒbyi���+�t���������g?~��E���l�����;%�^.�>���ipж;�/���ųgGF��ڵcaN6��p�м�TVpxՓ�3�K+E�C��O��@mݸ	�J�{�a�f�:d�Ֆ�8оޮC���������cˋs�-��x�1?���C#�R�>ƤnoU�����R�5==��\�43��?����{഍\�>4�~qy�]q�Miɒ�u�K�i"Ќa�� X0��@�T�ƍ�M=q8���2׼V������|�	��VL�f4��i��������Q����ճ��@OëK�A6�P�E���%�`�l(d��hyE�dcK%���<{F�;���O��IA��ҩ5�D|�Q�f�x�Q��	�2��5±��6V��Q�P�bEIB?�ˊ��Ȃ��5/D;��6�sf� N8���׾�+���0nPgA3��n���x�.�iM&��! 7���,7�M�'g�_~�+Z$բ�}�vf�gsm=-G��_�(8�'ɖ�hU�p(��	�@+�k׮�?�qPͥK�$ȴ~#L���Y�4��%��!�����ZY�+�����a�3|��w�������7�5ْβf�	%�}�eA긧���ONO��_�u�� �eۮ]0������	�ܖ-[z�ݻw��=ʉ�+��C��V��x��;�����{5"�!��_<~���x`��ʥR�] � &�#�؂�j?���|߾}Яآ�>��n�J8����������As�y�R���&��4�8��S�gKÆ~�%J�J
��a�cT"Ø~fBvnzĆ�jY"�r� =|�3tIs�գw�8�+��w���tv,��'_'[�|F�IT`e3I̬j��K�l�4��� �7�|��$���'I��TR���Q��������ڦ�9��g����5�K���M���fܝq Xz�6(�[��ֻﾋ�0ێqS\m�$�;�ED@ X+s���h��Z�8�S_u���'�3�A=�����̳ɉ[���z�*0�4��h�����4���u���G�F!D�=_�MW��9V0FL�ό�#h��3{".�N����c���.$�w4¼jIq4$���,�k�M ��&�\��~������f�W��^_wx�w�U� q�Ko!�~�AV�sY��a_���|�I�)��Z_W<tرB�V02�D�S�啲��ͤ�9��˔FFˬ@�� q��&u�����a�!<�WX WС��r	Gi�4C/�IH���!��p��V��D뵢.����O��� ��V�C�8�������)��*%t��;v@�cI�|�5P,�c/�øZ^��� ���.fI0u�`-�~ur���?��~� �Ϝ9�����d��h��ŋ���sO��UI�PF��0B����|E�9��Z�������w�J��J$���'X��������+l��=�3�t?`O�%����@n)����k���~ذ�Oz�0� ����'�l�������?����~o�g��=Y�i2(�iU�A���j��i�X��J6HG3t��3�Ϯ:nz�n5?}ŏ��pMpV��d���BL�uKl�5��Ac�����]M�k(ST�͔�Nbz
�J%Dِ�-/̟<y��>�(��ׯH���\�D?:�����Uv샡v��><v�X_O7��~���rY�|X��D ��'U,ڡ����4F��2&%/��s^�r������O�'p������%L��=9>�Mʼ��_��ܲy+�Ν;ǉU4M�򹅹ف�Xiyi��co�) �Xk�D!�`���Ц��{/V;15{���8Aɟ�ӹBa�捃�C�ׯ�����?��������6���xL٥D�v0� M���𙷛�V�l5B��(}C�uCXZ�� ��>�r�\��R�"mZ���2Vu�V�r�w�� �DC�@nHԪQְ��VdM{ξ�}?�K��yvL�:.W8���X�J�'*�m(�5����I
6��q8b�:�elB�ua�3�#%)��\[� }��^���8�Y���===ݝ���د,-����.���)���HX^GG��֦���J�ׇ���޵Og�@�7�y�c�:�j�������~����2R�- �q9�	z��5s��ݦcZN<-��Z����D�o��h�=�x_���lߺ�s��)\���O<��ŋ���+�lj��Y)C:��$T�6%��˭Y����5gW_����ʕTG2_�r�'3qZR��f�#�n�8���R�.D�5���/���4?qǊ��fdY��K�ٲ�ZM\���r��_��5!#��j�}���xj�և:A�7��0��G�e>�)�O��t淘���J�5��S�)d�So��$S2{L�2����"L�\67;5����R�W�gRiA̒Q+��'&����a��H�Db�`Z�J#�J6�D>��z]ߺ��-��pZ2��v:�.I��*P,���;a�l߱�z��wΜ:��&����R"���IvG���.o�&3*[�6u����g�ڹs�sg����|��ѫ�/b7FFF���7�L��=%��t�Fŵ��������l˘����]�AV����[�VK�_�����R{W7�``����p������L<s$�U�״<��ruW� " 8��ٹ��������훙��J�]�pq��=��L��ؕo�Ͷ|:�L�ҷ�z�#X"	��>�Ʈo������R�7L���\>E��1���+��H���k*�����Ɵ��w�K����a@(Q���)�g��Z��C�H�k��;�4ԲZ���6�
�5#�����{���]s�Z���o�/��wB�Qw���r2������9����o�����@��Pn�zf��.�,��֍��U��$/N%�sQ-�����Ѡ��L<T{�=�1,|���C^����mnzO�u�V���l���eYehF�Ei������~�ڵko��v�LҐH��˗�ȫ�]R���؈�J"�*l����C��<��*��c�=���?�~�&�F��/���[)5�<\�����
��{��.�0��pGX�ؐ}��㇟��'��`��:��|v�f�����?|�=��3�b�D*��l��=s�4��ɏ�ۏ~�#�d��z��W�3�oذO-�C��.<����7hcLƱ}D���)Kcu:�o�~F7�c}1��Ut��K��T�r���gt�{�ق@i8nPUpG��{�C�/���]��&�A�F�V��XWt.F��W�h�D _�B��:V81����>99937'\#-���FFX�V���tk��,���[:4`Ю���|A���Ukb[�^5�nG\��&0�HL�����$��`T*<�)���(�n��Nq�]%	֔�u��:^����z�*�T`h��X�-[�&xAE��`�ؾe�\,�>�vn�-(b�&@ o��P���*�51>����g�Ⱦ3Ѐ����m`i�8�%9�9�s~��z6�Q������D�����oB�w��_`���A�"R�J�VؔQ�mi?�˶Ar�<�0��7m�ʁ� z啗}�f����C--0)[Yt:�gP�E,�̀���Ȁ��+�1ШI�T��:$d����Ԭy����0EERĿ �u�֭3g�P��,@f�r0��X�F*���]>���kG��ʕJ�D�hx�B!�*���g*��C�B����<1|s���F$�D��.�_!����G���k$��q/��eF� ���3�,P��zX�G����P�{������>�̿t��b�_�.(������
]�K&�d�%�8�����!:"���R�\����;N�r���b��|��D�ܐ M�2�E�c������<A��	A}�_)�8^�Qe���j��ZL�c��Q��m������ݦ{ﯵ�|͏Ft�²cR�E�٥,W�;�&��WV����F�ƿ��q\�Zc2B ���TZ˸�M$c�f��	JR]�=�;Lưr�ѯ���u���r0�X��ܦ�ť���C��c]�-p��݇����+P3��st-�^�TZ���ڵkjb��?�9��с>��'�=~��%�ӥfg�	��eܔ��qCP�����}�v�V�h�Q���D,������0�����}�;��N_����Ͽ�گp����T"9;5[����O:p���
^�}��������~H"���]�� <��W=��cF,�裏�����9�ŧ�և�{���aPx������w��/~����3�N/,H��*���O"��T�y�.Q�$�S�ԣ`21�#��+�;m)*$�'�]����B�*��`h�&� ���J�/K�B_�~x�[�M)#s�R�`LE�Z�q0u�ڝ��ޡ�L�����RS�����kjR���"t��ʃV�eC������T_��4d��X��p48�c'N���ˁ�� EN^XI͂_A��X�2��JvE[[���ٽsk�"�-�O���L���!�F6ۡB�T�+�TX�ba=�d�$Q�x�=�F��\�Z)1�Ѭ���qA��ƫ\*�XN� ��X�f�N�n[�ڤ����'#��ux�3���Ʈ^�r����,��th���Aa�V��q\�e�8�s�c������m@�m۶M��������㒉B6���h��ř����Y���y�cF63�@k���OшY�N^�d��m` X�����b�I���ֱ�=th��7E��,R�E��� /̻ܩ�����;�M��'2�@�ѡNa�I=��g��b|.�oe���2$qv�߬L���%�i��|I2&��R���$���K��6q�j���1�}İ���X���ɤ2Fg+R"[��ܹW���aaBÕ���F#'fI۲cKc���K�����up'՜���%�ӄ)>��Xo�?��v���Sg��bx�Gz{�� "[F"�e��l����8�	�}KO#[0_j��l� i
d����ظD��ݞ>(�=��3[v��-��'?b92::��@�]�|	*��X�@o��\�XZU���Ԧ����PUsӨ�\j.ť�hǲ�{��g�у�?�x2ӖL�˕j�\�}F�&���ٍ���^��-�й�Q�ߪ�M<�>p�"c4���� ��|��?�|mq�u��̸�3A��XĹÒ�-B��wpGd��w-�0k�p����&��^����<���W�R"s2J�0�S�V��(K:�'���(��
t�U����g��b��>��
�`�L;���2F���s���谖;31e@S�0N��_�N8
��@�A"W 4�gϞ���K�.��YGJC.Kd�P���U00��!��[��?���A&���k�~��<���_�����j�W���
�nhx�� ;&
!�K��i��v`T��?�3���g���;w{Ϟ�4�``?v��)�կ~ux�z�
W����o�A�=u��S�����&��NKG[�� !n�g�z�ʖ��<x�W^yN'�i]����w����cG��Q�ف�?��?�ۿ��k׮AF� a�m��m�VK粸]q��nA��	j¡�P�KO�)�>��kǨ��'����g"%Ѕ�kh�3�|MysL$3D��в�����C��|�?�~����5W@�b<����B��Lly��Z�����&D>���:o�8�W0M6z6��#�cRB��U�T�x]�x��w��:���c�	Q�X *�5�qáO�6�c�9G�tK��@f��	uwt�]�ݽf���T�:X��0�H�Kӥ���CqBG��4,t�������./.��e�5�_'����g�������M�_������|�eHN��cU6!�e� ���ØVG��|�S�X���������ἠ��"c��\���]����ئ����2�ȴ�w���2����C���F�q������n޼���H4f�N�
��d,M�/���	l#��
_�?ȆE���D0�	�v�T46�N*ߌ��ti�2u[ahbz����7n��97w\]�Нo�k`1@��څ��V�@�jj�S��n��)F���1ÎW_�.Ϝ9s��!*�.���cǎ��XI:�!�S ����ԞQbN=:�mX�%��{��{�|9{��ح��۶�޽�ǿ;v�8q�]��AS�D�R��7�V�fC��]�#`i�q��R�g�re���8"��UmtuvX��SA�E��l���Yq�p;*�d��?da�,:qN�s���) #�Zp!"A��5N[�X4D�D)3�������A+S|@R��"4���З��I�ﶀ�gw��ն����"���pS��k:�����$'i�]������BM�;A���D}ee�hV�����4��6�Ѥ5��ZJ� "�Z��D�Du[��E�
���e0̾}�z��O�>�A�3�S�s�d�Accc���^��J���쇰�5sct��{�p�y���3g�x�	\<	�!Px^s���W=�=sg�|�O7oބ&��ЁK$�^����矟��������[7!bF��@53ۻ}�o|��K� ĥ._�{�e��_����H�
�F��|�W��s=�xAL@�I��N�ѯ��ʤ��Z�Z�Ա93ssK++۶l��9q��pp��'�|�}��������Z�t$��<�1�B���$^̬ �e��"UDb�Hb������p��f3��SՍ0�-�1x�9�J�� �BD��&�Ek�B���?�(����ʪ��
i�D���`(.L������<2$/H�&�ux�p����j�XYYeZ��&��my��>??w�ԉt*��Ӌ+$�vO/�eEFzf-'fT+�R���*}4�h���dS�m4�(�#�V������BwO!_H:���MeAo�)�-�.�KF6�K���t����μT|V���uvu(ز���J��m�~suqn�w����&$�r����������67�'��3�&��N<іͤ�b֗k��陸��5�`4SdHN�\vÆa��XF&�ޱ}{&���y��(��8���oNMM��hC�܇m���V�qg�2hHYd&��r�5�Q�� �l� G���Yk���07��I����b�.+-p��m`vB!2m�e*�7q: �,���ƹڐ�Ţ�;�� ?�0EWWGS�c0��l`.#)��re�Y|b�>��Xi����[,��]x�{��7��[o�337�o�~���-A�N�s��e�m333���'��ٍ�����Z����&��n31ޡ�m˱b	3A���4<8-�K)�DfA����`%!�>Ч�&��D����T�`���~3���`ԙ@����G�Z��}�z&Fo�={����a����У�����?���~��׮K��9����[��"2q�̚��iH���'�|$��	��,!-�k�!d���$A%I�#����4��b�4[�\$p蹜��\�$�Z)�-B�$1]�S�1�Զ�yW�02Q�Q'�Y���᪽Ȏ�}�wD��
7��9�I3�{{������x�(B�Whjq�}���_�l:8��d+��*<���~���ԢE��Y�fR�P<nN�i&6��h��cZ�]��EL�?�����B4U��tH�p2����xBE����IN
��k�ٲy��ڍ<ڃ>�/�짿���e��@���^�@SB�|�s���W��7�7�U����6�(�0N��bV�E?�&XK���� ���L�n�r��s��-�-�����p?��O~���Ȉ�:�ܹ�G��7l���§�_��7-�~������~���L�Iȳ�Mj�Ν����3�l��8_�����I�GJ�]������a�
����{��=�g��o�^�%S�(���!l[i�r���,�/z���lF�ʕ�\�� u�~��f۰�oM񈉣Y �D20�Nr�6����BI���*��`��o��_Q1��ע.$�4}�\c���d��� vI�u�cq�+�z����i~T�!@sO33s4y�����x�&'���K��'�,;w���~�m�rӒ��rI�)gfՓ!����B[��--�0fI 3���4�^��4��8�������Xl���#���֎�T2���)�u��];�6��]����4��@�Ke�u��Y���ߜ��&���w�s��&>[،��hgtuu��)�q0>��_~���w�{�#�qM<#�����eW;�`���V�rt�"�zĭ9����+�%��§M7��q���-��ۛ�/����]q�;^�5�V����x
>7+U���!�9;"WCI��#I����̀蒾�v��n��{�)6ś����o���:�$wX�E�KM�����(��;v�K��	���A�1[��u�������n�`���1,u˖-����u1���"��,�b2���l�e�I�}Jj*d50la��K˻v�Z�1'�Z�!Q���֏�6���Q���Ӛ܀[��Ca[��g��ϯ����3�{����u��-..`�`��:`F��w���T��k�S�Y*�[�"�fkrƮ�3M:��#��m��g�?%c������bT�.��ݚ�j�ZrS�nN&�k���<�xD'.�tC���n������&&�+Hf!>hD���e�ފ;3|���XC�
���,���|O �?��+���0�#u	�Z�R��:Ĳ.���D��/�d�����7덮��tBV�~��J���"1Aӂƅ4m�q�)��p��(�Y�$>e^�zT;<Է��$S���8"�ȉ�:	gqf)ᘱ��ĥJ)]�B��w���uvu�3y����XRsҨ��h��ȱw�|����*��;ڻ�Z;۵wϏ~�#�		���-��*d����-ϯ,�.�=uf��� ��-k��M�����w�\}�}��׏~]0���L<�8�h6d�W�����s[v"���������W9N�<��w����-�65wr�f!S8pρ����7GF������q�U�����d��~�k��^��4L���������%�Y�]m`]���Bi��v��]�����؝J�z:�{z���<�J����.Ke��<�_ʟ�s��ޕb��N;���$��V3�-�/%���z��j���c�T.[:ɱ
��ѷ�J������,/m8��h+����qG�j3�l -�O��5*Uߊ��	p��W�D������v*f&L߭j�Q�Ա�Nj�T�u������zn��ս�7\�s��b������?��f�0�8���Xl�T��ġ0�܉Xʴ�t�mxͺ���[�hH��;�:�fj�;�����q<M���F���{{�	�`,,��ʒ6PCJ_K�2H�o�W�\����maŜjcη���Ex��׻;{ddg<�Z���L�3c�<Ⱦ~����[�][�n����ڵcl���+��{gggO�0�LFFJ��dXM��:ڻ���f
r7fZ���sP�2�
�V{^r����x��X�4��Ay�X\ʄ�2X�QWhK&PA��;������t�+W����(h'�J[ݐ����WZ6l��({~}xxH�X�]���Ky�G6wn݂E>|x���6]��V�5O�z5p���7����k�6mضm��`/t~��Cط�������r��*�a����r���)x�UÃCOŤ�qaa�Ѱ��@�ݫ���К�jX!#W�K��sK��;W�X"�+�S:�Z�,3���3����6�P$��<Mӗ�PW�m��0�����V>R�4n��������Z�HTˌy W�ЗI1��Hv���\8��Z�l�l�}���:
WF���]����z�f[[��]�������g���J�c�GG�5����ĉ���g�Vd�J2�L�N"���nTk�_���2�lP�
B��Y��U�N'��7ƽ��O��
ȜX�#�c=��PR��/��ד�ޘ���j/k���m���������|f]�����?���?v�XG�:�{�_\X*dҬ���+��3���힝���E!�,�ē�,	(&�Y���T띜��|�.eyb�$�x*��ى/�z�l1�`�3�V�L�s�	��X*�m]�<�|*i��釠��}�O�.�ѱ�?��!X�����m��Vp��z��Hϵ�j���WK+N6+m�9���2ĭ�k��^`|����̶�;�NÌ--��{｛7oɀ����I|+&�8#�[�TK��@e,ʌ �J�N"^��:>D��Jҽ]�|����l+tB�ի6��4A�ؼ�U�~�w�ɹ�R���s�+��hϵ7���sdZ�fg���4ܲ449�+Q6�p�r�%^�4���76Iܦxg���Q0!?�Z`l�V.,U���H��|S��
�iʴ(�4�P�`͵f������~����X�y�;�35Cle�:���k,�ƾ���f�3��B�`�P"	|�ւ�a��5+�L���!�D�/gia�F���W2�1H�)0a���7m�
}��-��Y��ܹ������~�|��O<�y�F<淾��.�Z�cQ��<5�JH�g�}�;���Zu���7�(6���T������#sX�Ew^�߶m�(_�q�(��ׯ���3���4�o���x2�gϞ�~�{[½�ff�GK ��d)V�#y��`��Cu�s�=�;�7VV a�a2�q����b`�+.;	3>ζ�S�N8p�?�i�Ո\=nH�)y�j7"��:�f%���T����Q1N��3sC�	7�A�=$r5�"�;CP���8����0;#na�m��)x�/n��?�;�����SSS�:bZ�^s��&��	�����v�|�>��}qy�t�Q�ϸ8����%�F��NX6R�w;.U(丙2��k�;w�;������}�ن��A�c1OVB~P���.(]�:�PP�{�e\-���~�4$d{J!�:�2���i�B���B�C<�����K\Y�E�l��bJ�zju)���&@�j�T�x��N�:}����M�0���l5)�N�)n]Ja��rs���l����<����o����C	��d� ���Fw$$.����c�O<����x|�kx�ё1�_֫E�|��4�(�P�K�.u��E��E����o$��G�
*ut����$�N�Pa��==2�����cc7�A	SSO=�Ժu��v>��C������"�O�V�T�Q�B6�����0�,J���^<#V�a�!����/�X��_\�Աc��!_z�%F�<��!
�Ҙ�U@B�����a�0����?���k�^}���G�
�%6aEҵ���M%r�~i��,N��V���|���Yl�8E�lH,�^	�����k�.xS�XC� �(+��l6������aa۷o�N�b����'��1;7�;
��`�|��R�O{�v{\D�]#�a�H�L)��x0��[�nf �kj�*e�q���;bD��?�VJG!*)�͠Dt���9�^C-Q+�߲�x맺gJA)pm�3co�>#;�.�j��Z�C㧕/������ފ�՟�����e�e�����}�7��h]4[�T�TT1Ct �;t��$��H���
7�b��TCT�]nկxpB�Ae�eZ0�Jt���-������.רU�d�	nޔJ�+�:��A!qד��a\�*�x ����3��;�N��!��C����Z(����cG�^��Z)�u�
I���%�����W��<��g��{�͛7%�%��O`qi)���'*i���l!X�V�����<jyi�>�_*۴y���",��90��_�_?�<ߙ3g�qx��g@���T__/sF�I���4q�QWW�x����N<E{G�ŋ=�-����|K���;�\1����>���OCꭖ˙l�Y9��q��Њ�l͘��)#Ϯ��j����u+��bȅ5�>\7p��/�7�le����ꢏ� ���#k��ՀK'��ۭ72~������y�;���s�!e��H�����2{y����Ծt�:�d�E�̬��񚮂6�A��$ш���fP����p=�U�/\(kz���BE6���t:)���$_{�5��4�hp�8�ՒL�0��y�e�񥍾�M�v2���BZ��H��O~o�Q[)�2ɔYo�U�e��Si�)]�ybb�\Y��U��=�2��e��e�#�yoo��)��w'ii�r����K���C�Yv�����Iq+��m���.�߿��G�8����,�]�(\�V���+T�rGw�޽���d���݋���_���������M�0|�VVK��!�h�$��]�k�b<Qoz�������b���ླྀ���[Z e��ڱ�kz�tg %Z��K! *���b�E�񣜑lJ����O�)6���qǭW�}g�ָ,MA�q4z����ʦMI�]^^�O;>>	�G&��֏ã�8{�4�E`�É��f�^-W8���]��-�޻q�0�$m"��m�7�/HS6����L*���zd�����Xv®p|>� �bC�`��M�h���'`^�|	�M{��c����[,Zs���!q�Rx)��e�,�YA��BC�3�F��dؕrEܪZ��Zu�Ғ	DO�� �4^Yň���%א�����_y�QK/���=��^x��'���o��;w� +:;���PG��՗6!Y����"j7u|YQ�l�2�eHYo �����(��$/�Dr	�̵�' ri��}����]�P]['n+������L����TpT�4W[�����HʹcG�|��n�z?�*�ߓGZ�o��L��3�C���G��]쳵K���#�/CI���a��J�˓y�^��*Z�,��wMj'�h�"	�j�Υ���N,`슕4�o��ްd�**��M+x��A���ÒfѠ1��� .Qª����Ly��wA�`]|r�֭��1;�%��*�nhh��ˎ����+_��Wop�'���.��5�GO�<�v���a��������ٳg�:��W�4	�*��ĨRɏ}�c��Clō��!K
��0�M��F١u{B��������~�����>b����=��L�D6��L��>��嵫W�rs~�СC���7�9�Y��`����D`���$k���D���V�ވf�4�mSE�~�W���]3�RS������a��(rM������̨�������sa,gQΥ�ީM�Ry�!��`�P?����8}��E�-Y�����-�h&�H���х?]�vu3^[�ȼT�R�����z�+.�Y�����$�%�@�.^�����j��6O�ݳ����[��rض�` ����{�n6,7B�{V�\�|Y}|zf�p~n�eXQ�*�c\���
6�N�9������UGy�5,��h��l���ڵk��!�o�&%��'��#�y[�6�c+3�۷oǥ��o���|184,�\Y��W�c6����F�P:1)���J�ڨHi��?�y�o�B��3%�0��+l�"d� ���h)�%T�W�p���>���+����(`�-�V�%���9�"�d۔�6h���ӐQ�C�R٢Xe++��l�6���8 ��dT?4�'�q�bRڼy��nB��q�L�@��iVdr���1���',�E{��J�5>��
�L��� P�E�-�崘�4[I�,E��`�v׮]3S�������/~�~GG}y1�镢�`RB�ct`��"N�N�-�K?L�-ظ�"R�R�C�!^7[��)����%S���6�F2E���̹���^x����˿���n�"(H���Ӌk�A�E��Y�̩�k-�%�R6��\ H�s3�N�E"�0׬+��n�)�l�o����<	�0�1��_3�Ak��#h���Pf/ 3{׶bw���j���eqA��_�{-��
��]Ɨ��T�/���u �����ߒO\�R�2B�� �*��&�Z�x~8iA�uP�ߩ5��j�j�=�mM���=���T� @>�>K&���r��lNz|f��¡����������AR�
���2y����a��ЙJ{a!�e�=Q�����z;��4O�<y���m۶�����1*�FKK��g���fٽ�g�C4�m��jd�E2� �9�CC�H0H@�W�\9y��SO>��3�|�����
�U�pk�}`{A�gt���AN�8�
�;��֧�a���J	>��{����R��j4ݟ��߱�Օ�B��6�۩�����K����(�LM�V�K�8��>�	l�͉q1��b=$�Ҹ��	�E�R�HGgF�B��
�7lx衇 4����ͺ��)R1�0��]�r����i��AH7��~`lq��X�3�a=����+ �.���,kҭl[�5.�XB`{��lȈ���Sԙj<�C�5ރ�-�i�� 猒�=��Xu���X��ػw����G��u���+p��q�DB����ɇe��r�a�W`1�y���>��7����7�)�f�ƍ�Őh�-8�������Y�.0eLC&��/�����?p���@�Ps��F-/�F�(<Q2s�l/dA�]��-k�Ɓ�[7�)����0����c�b�����F *��];6�LK%�++3�եz�Zo�̦U�	꡹�8��×����)&��,��(vUzY���鉸 ��A\i.�cq��>-��ٙ=�w���Bh�
qǙ���&�R��X���Ȥs=��u��g��q{��Y�x�=��[㓂���S�D9�m��3Q�A����k*�s�<>��4��}�nH��s��Cԙ�zAa�Z��P-��ry;���Pg4�ha~�
�����˿=�F�A��o�|��qΘ7�0��L�O-,���N:1�ǙJ���~���C&�@�d��\�����::�fg��4UJ�
%.����C�Fe$�c*����8�8���^���UYX��=$�wO���X��旖���`���VQ��F����3e��%�%�:���ɰo>��W.��h��8�<��I�HYN��ҥj���?�ϤGGG%��D0���ѐ��aV.i�����_\\����T��S1��FL��d3��m��ذe׎0��Zm���;o��o�!H���_~��Y��ȕd:1�a�Z���~����pZ�'4nZ#�QĄ8>��p>�籤�7n5ju�,4��)b�XDZ���:? ��}��=g��uZ�YSJ�L����F���TV�R)]w�F0r��#�C�*��"���#�K-?;�[�B��;�3ߌ���V���8c�iM�����Y�~����g`9�B3�z�m�c�$�|�WٵKpsFw%Z`9�geg��]�&�h����3��rNEl���/�z!O�K���Ȱx]�6Ö�tC�פ%���L���I\
?ë��C���I`l��Ǐ�&�0=���ׯ_#���������5A�Ԋ_2� ��<��S��Ʒ��!Mw�P����v���zA��6XT�[h����c�샃��9Z���H�ق��	�T�9w�q)*u�A1�)]�f>5�"�C��ݲu;��{?xQFu���E<Z{���B�?w�b s��x��'>|��qhz��s�ySq�ɰ��'��߅��2ٷ�XYb���̦�Ђ�O9#]���x_;�ʤ��O6yq&i��%U�L����D��?�:#�Nd_Sf6���Q�۷�����e� "b�wu1�Ǳt̞0�-�7bC%��`1�?� ޙ���1A���解�'իS�@`�L%���{`%õ`�� �
��]Y��8M�6ٜ�6��Lb�6l�"�}�CC�*�5 �u��M��e� p�����D��ܴ"�RY����J%����,��C���|<`�m�>�1��<��#�3M�#b�����e1�]W�ɲK䐈G��}�m ��0��Ӂ�ږo�-]-��N��C&s;����Zpc�u���<Q�<8��ٳG�y��xR8b<�M����^X��B���nIƥR������0+�vG���;���>�U��k3��)��ޤ���*�a��tp���݆̲��
ҝ�h����Z����.]]m�f3��R�N����7��Ҥ
-��;����޾'�xbrj��4,u�8V�8�<9�W`�X�Mޗ��Łg�\����j-@���!r�U+1�j���+s�?��^|�E0��#byv���!��;�"�#րl"�m�����vJ�1�Ex�t�eʅ��ҪA�Ű��>� ~�p��a�dgG'.�uu��T��x@
�}������ukÆ�x��I+3[�e�|��4g��h�n`{�1G�L�{���ub�[o��s�!�� �R"ܖ�cK�C�uT�r��L�&��}бa��e��D�M�ǧ��C�Vg��A�Ti�y��"�;὚a���^)����X�-���3�4��*�e�w>$�y7�F�X{_��fh�>��k~XuޚVč&?�;�0�!�&m��6���?�-���t)�u҉;�FM�� $@+���`�lnni��Z�B�Wˬz��M�M���N%�1���1l�&P�j*{�V�{�D.�½�\�!��Bb�A�hig;r��k�.�s����_�{>�O���G�!��5ؿ���O5?��L��+��S�7=�أ�.]����J�{ߋ�MZ~*�$�~���	9¼�������������z{�W�7*�s���jWg;����y��R�fR,���`Q�b��V=�wJ�J��L�N�Ȇ7o�|�g�;v��<N�����
���K/5�n�n�2��?�qt���}WF.NNO���w�AF�����9�f\3��a�+x+R��8�vP��J��$�Y@�Wm�S�M�ڎ͡lZWb:� a����)��u�zO�4��M���]���hыD-¬���nMh���3D*�m����
ԸEa��&���)�^hi��i���� >���W!�a�]�~}rB�ILp��3߸q��|����x��WW˰��9��.<ȥKW~��`��L��8����l#�MgS���.���l2��5�wvu\�t��+Օ�%���v	��v�1��oVJ��U��+��1�f.+��M=[,�d{e8�k ���c��Y���֧; �ryu�`M_�$�@����b0�RG���H��������ĒZ�V�ɀV���_���ٲmG�����ٱ�'�<�Lg�9ɜ�s������il�a{�Nn��@��vI�=(x���~��O>�6M�M&����ʈ`��L6\3���ȩ3�^�0�~sJ6[�:d>lO�Q�i�D;��qM�AJ�,��~����lo� <^O��}����S�1MO�g�G�S�]i�U�CZ��Wo�Ԧ��*I8���Ip+�҆���<��W/�X�D�R���Ic
��ꎎΞ�����!�^�S�J�A������+�w�ƙ������u�/|�P��N	n$l�\.�8?bh��-�g�Z*�й��a��L�gF�\U󴫻��*R�3œ d|��U�)�[F֯~������h���.�W���'&z<�<?O���Y��*$�Ԕ393�����\���Ĥ�j��7����{ה�皦l�E�Gˉ��
��~*��*�r�0���z!�	�YF^�^��fs�̞7��"���|Ʋ!�L.��m�*��1�Z�v5bgHޟ��:�D<���9�+�+�$ZゑC���m�!�A��Y����F��g�4�-���̡���7�W���RDm^8��U�L���sǲ ƴ�(�b�+����4By��1�ڶ��ق������tFZ��8E�VR�B��G�s�d���n��:3Sф�@�CC.�MHm|2�]�`�w��q^~�e(����Νccc��qID����y�fb%�̀�~��_����\\(�1*դ�Qq/��! xd�	`aY���X�	u���ޞ����X���T+3�A4]�<]V��E$�2�C���p�:/MP��7L������L|�ɏ<	���y�V\��G�������!~��'�b�
�|��p͂����N�r�c�h�0	Nf�@��l���E�� �ֈ���a��͖�zU2�
�$��~���R��!��~��"��uߖΆK$ŭ_��g��PW�0�@3j+�_�NwA�����~�[�!�������N17�����x�ntI��r�
̠M�6�R�eVsq}0�o�1 �-���x�'ٍq��}�"	"Xi��س{'H4���!xJmj�g�F�LG[(���iH	���`<2��3A�;bxq�_)�pefTY�îj'����g�/.�O�2۫�eZ6�B=�����Q��4�a�+��5j�`�rȶ��"�~��_|���������Ӫ��W\\�8� 31��i	�+.�� �����f��K2�)�_g�NC�����c���	�f��x2(2��{��F���/�]++:��W�E�5��H� ���XUɵuR� �	��GJ�uf0�3QL�Ah]N��ژ�&�����  јN��~a7VKů���>�^G��!b�&�c�8#�c�P���b򅵁�����S��ŋF8��!&�{b����/�����������_{�U��,5�
9Gall�%bx���^�G�(�2�ވ�﨣������R��$%၀5Ɩ��A�۶m�V�}l�tF��j++ ������]�u�u��;r�V�u��uh��~���B�ƍ���~#��Ӊ̋���;>6V��P��E�~<���Ss��~� I���Y
&L���V	�Aa.CicV?��!��}��,�J#B��FmB�+�L����p�G3����[`ϣ�Ydx���)����~  ��t�s�E[�ћ7���Q� ,�j��D=N�_�QR���fH���n(uO*��_Գ��Y�^�U#ϔ�Ǝ{���"q���l�i9����2������5�4��hqn�t������,��w�F�����e��m&���<_R'%�Y--��㕥eǴJ+�z�:zmD,{�������rt�q������S�ϟ9���	�=s��v,M���ĠⰜd"��s�=��C�~�U8j�i�&�����4��ʒV��vuc��+�27�\��vp��FO�0}����8ޤ/7�I�8�$��)ʼ�ۻ�L%�O���
h���Dc�XF_w�Xu!���җ�%��#�����G���q��X2����g�`��]�2�$���0�!t��փaSN�O$�4���-��B��r}��aH/(�	��a���.Eϳ���2�_o����(k5)&�'���-B'�12�
.'D�d+����H�ܕ�yS�{M�}"���2���;>%[͖�l�f�:б	D��i������� g�"3�52r������@�2��YhL��L�X\^���~����x������m�²8��ݐ��ssXb2�U*�L���<-�"�$����la���v� U,,,o�{��7�yu���s�WV����\-�I��������к~��8:?7�ކ�n��6<����`O�U)��zuaaQ���p�!��azkȤs�5I^T�a���p$s2�n�ä҉�Cݥn��-��qe�4`m8q�XA�i��,�K��и��D��S��/.3��������Q����l��}������_�}���޽g`h=vubf:���8��:��w��V�/H��5�U�;:ڴ\U@k��w��P�m��٩)�?`����rq5��VJ%�CJ X��<Ec��O&I�,����6nwq#⼛z?T!	�����蒋�K���T���F*a���׉�iӆG}tff�W^I�Rs�
t���X���Fhz�\�*{�L��De�i�����9` ����e�a)f� �tZ\����[��=���#�w�z6�w©Y��L���mh1>��СC�F�&�ɕ�J&'ސ�|5�&��J��&���E'K�S�?���'�����}�s7l���W�M��
y�lvw�(��NȽb��ѐj�B�=O�E������!(�;|������}��&�-cl�,,��.���Q�%��l!�Ƙ��w��'N��>�N�''Ʊ�L6W�V��m�����~O&�=!��al�e�X63�xp���M6��"%�7=VW����/]��H�[�33¨Jӓ���(I,�T�[���9=;�Z��EO�$.�p���o޸�'�
��8���Io@�$�!}#7+U6aC��[�Z��X�8���hҨhGLg���C#h�!4f"{��Z�\����Ys�!ku`���5�Sͨ�c���R�!Ȧ���gf��� 3�����w��� �{�Ma?��>��Zt�(�h�.V8���+�L0�^z9��=S��d�έ[��A�,��\XE ���ۤ$��?�՚,P���|�MK�������`^0-�)v� �
�f|g?22�7���K������z�`NP-����:��߲T��i~�̂���9ƓJ@D�_�Rh�)����?�A(E����od�D����j�JlE�
PC��I�&طN0�pӾ����;w���>��g
��x��Ǐ��@{˰�j�
#�w�l�B���'?a�7[M��c�
%����[����c� ��ᱲ�T��Y"w'*L�<$&)���e���cҺv��u/�H2C/ͺ}���a��ܪ�pԈ'^)�A-����j��}���Z�ޭ�lq|Exo��ੱ8�Q�Z���$m�OV$��]�!�5\{嬺�-��q����s���pӭ[��>}���u{��ڔ2�L���b�09�m���L�����SF�I�`��0f;1�T�B�ܝt�o/��{S�ڧ�'����N���ظqcÕ �ey��,;DK�%U��	1�x?�Y�����?���r�g2����DRP ]����	A�ʦ����r����p�&Qk�ηZ�&�3g�D]��A�>��W�^_uU$���,8N���������������
D���`ϟ}�i+'��S�3B�FL�4u���DV_��X���iE�$d��f8��U�wXDVب�����CdDn�L�$Ah�*p'p܆f�ymN��AS;(ls������E�z��0�͂��A�tt͘8�nzct�ܹs���x������#o��t���9}�sR%����[�A�)�A��x���H��"����nϕ���i���^�u����d��n�կ~W��?�����C��<u���d����
R��i���4]q,��~�4�ò3+�u�j�p6���'oܠ�����y!6���ٷ���~f�&�T����!U��ӗf���aŜ8S�V>?�ȱ�� .�M�u�4�5��g�OA�'Tm�5D��M��4��� Ŧո��ɝ��V�͵;W��a�mw�"���j{ǚtƁ�Z�VK��TW{���Ն1���^�V�A������Zq��і�mR.W���ҹ5.a�U�}O�#y��7o��ۤ���g>�x��;gϞ����`�ٵ+'�R@�e��f����\�o�j�&1���y j��t�N�k~n���s۶��(i��}=]ݎ���t�Q,��wTjN�I�n�V�~C��
�:c�8���T�����`��X0���#hp�g&M\-6��t�6��£�E[Ȥ͆#��1�Ьj��*��I�n޸����oxp��{�bp�z���Ò ����>��\>2���%�k8�m۶��fU��,-�<_^u8�ɴ�j�eBj�j�2���HO�c�Z��p>� :65/����<˨5$ O
��:P���4��8�y�xM��S v`���cr"������>�o�o�-e�~	6Z���v��&�jŽ3X]��m��K�i�\\���\\^�oM$f�mœ	�\a=�����&30�3�}

�V�0�mq��Io�"6-�/i�2,$'�H$r�A��.,,9�v>/��٣��;�c`7�soHx��AC��뇤�Al����9�>VR/U��|�m�֤�:st�_��;U��N���Z�Ch�t���:_�^��K���JS)aaI*
�f�]���4��rm`]�����++K�����l��R1�O�%An;xht��|	d;8���;�(��R�Ph�ŕe�p&94�_^..��q�JǝL*XN`Uۄl���F��N��r��%�щKV�����sg��w,�R*[F��Ǹ,���h�� ��o�2=�R�ec�ҀD[G{wo�����l�2�S���f���^�:&�7hl)��ԓ�h3Q�>mNJ'��<�'N	�i}J�bttT칢 5�����J�J���
�����X��Ms�[��lJPgw'�MN���Y����҉:b?S8�#�./�W�V�T\%����e�~?�e�]Ξ�Pk��<��#����G���51?+-\�tjzz
O������5��C#���.�)ֶxe��79�̂<��$P��>�i#��0�V9v������G�c AcO<�u������K++2N�Rj2�\����@���EGI�ǭ�Y���nwuqϤE���uwv�\���%]�vT�1�-�����Gm�O���f����{���S�Z���_����zKn4�����������6ǬR��Hj<�56!�o���1���m/��?�Q
��y[����/w�)d��~��&��r�]� �q�ɨ��5���:4��S��j?�3,�_=}��5fSP+ǅ}�%��>!$�ք��n���)W�:)��/���D>3�7�IM��`���S)"y2/	+�ڵk����;v��#��ڰ�|-u�p��E7zHF�_ů����G,7�8���f�ǒ�� (T��ZŪ ��Ԙ4��c�<��47w/�i\�_㺬� v6��}��Z����ώ�ɹ�j��{��}��W>��lں\O�c2�}����(�ϝ�:��Ϟ<C&�Át��B)hބ�&;��=s7���oo�#�y��ݥ���}�陞�3C�p��P�"��#�� ۰� �� q�?��1�|� #1`C��Ē��q(�"ErDq���ҳwO��ݵ/���s�s�횅%)�buս�}߳/��f2e�l �'(Hj{�񜶢a��E-@�j1�'�P ?5��0jw��)G���������|����y �:�5=A�K5��`4S5��p���$=����G\�X,�=g�?Ɵ�,��1�
�oG��v���h�znn��h�HgV�gIY��qp�k׮��{��`[caE�b�f:,EP5�[��8�$Y�ui�/�!M���7eu9������^Э}�����u�|Cm��l����5�T�QRam�v�� F!(
ܷ�~�U�J��=;;�i�3�a�J��,Za���ٯ�,�D�ܺE�4泦vLphԼr�
��57R������uiNR�a� �^���3��N���U|��(�J�c��]�k3��g��]�]�A\=/x�{������^��>%~�S�-�7,t�U:�n-�+�(���E��t�JЈR)�֐Ui���6�bFp�(&��p��T����Ú=pZ��ꥬH�F���(61�`j��L}M&����-���
�v�4�e���C�LI2��r[��i�M�:�,Q�L�4�l*Y�}��33�����u�����B��6[��=E�+�`z���K7\��]���f���|G/�����+h��T��s/�8 �/���7�|��yS�l��2�-],Ȉ�<X�J�:h���SO�:�IZ��4��4�LE���0�h�h����L@-��$6v���M�N�h�lF
�VW[8���Q�=;M�Z�jC��� {�{�i�L��,�d'33ELmY6k��0mb�ރ��ϳ�� ��9�1ui�����1���//�C�����;�ϥ�E�9 U�L�q#�#���r�*�d�tR�<�]���m#���X9[�|y�p���!�5�U93S�G+u��U�&�zyC�Y��ݾuV�7�6Es��1��ڳg��R[�n:=��\6_�5�_�� \����]]=�jP-�,�m�6OʨW��^�z�p �|�n �=��"�E�G�b�iݺ!�~!��F�[`*���!IB�S�T�r���A���R!+sʧ�� wG������u�Њ2w	#�m%��7dn��X*%�ch�\H�S�)Ҙ-���y6#vQ�Ņ��ݻ��|�񉥅Ł��|<Q�����S@K|[Kk�޽��uޙ3g��������?00��p��������?��Y�R�2�3��'m�d�1tv��:[ͤ��.,-BB�
T����$I-�X��)1�WHF�	���fpa}Î�`��Ղ1l�.4&a��r���9��u�wxu�0|�!�1�H;�&���|p��5�0u&
�O�U��!�`�0�
zoe� )��Hv�qUǙ��*�̴�mO<��O�*N���nun}viqYB���
$~O�������_;�Jb�Y+1#�=���]�x�^�z�,�K=h&�*Kk�%	�G���!j�p�QGT�
?�J#�m��8̰���|E�d4��A]ҝ�'c��<B��76����ܟJ%�K�ELdB2��F[m9�R�V�l�y=��Վ��ܹE(1F��?��x�,�-���?�䓏��R:�>j�S��#xc���h���õ�v"���A�6���)�P��۷�~�8���k5�� 5�0І
�3�z���/C�A����_Z�D��ԛ��t�ڮħ�G���M�:y�Z.�MO�3-E�H�f��Aq:��*����>Z$�f"�o�^_+�� ��>}�^%tGf�n�EgPj&�]��5/�3�+��q5:��SӚ1#.�Ⴭ���s]�X\��6�P![H�,�cFa�w�����h6����؉�v��e[��G_���w~�ܿ��е��*��#q0٥�ĶdT@�TM&�1ģ�ex��LZa�a��qI�؍r)�#��Y��%��6�tYIܫU(��b��fg��S��A��V�ڕ�#��=�]m�P��"tϋ/��"�΅���G�)�B	���ě��ݐ�+�K�(�M�ے�,v�~�(�~�[�b8�HV�ힾ�z��LIH^}ay��(���hJ�U�8����Z-�ہ�N�NֻC0�b�j{�c���6�k�u~���[fvT�����H�I�1����8�13�Sz��z����7Z�c�ȇַ��'a/��b��E&I���=zV0��k���n���N~R\�������bq�Si&�Eg(T�o8�#�:F�������b�&��(H,p��QH�7ù����@:,,,aٸx�_�I��)K�R>I:>����Xw��1V�H�ʑ'�7� �w��P,�2.>��Ǚ�7�)�� B��&bR��N"�. Q�Z�ƌ����y)VjD��0_� ��V�������ĉX9�%������p������l���ų@��W'O�8r����{|X'!�a�AL��%MY,hτ��ɨڔ���&V7����c���o�����f�9; ����_yA�0K�x��#s�� �\,bth5/��^c3�o*����C?1;::	���}�� �JMѕ�I�P0ʱ{;w�%�w���aX��H&|�Yj��ML/� !�A��[k\��Gf?� J�쟊�M,z��3����>d�#�9b֪D�j+�;l% �v�"Q|�ֺ"��Φbj��Д���J����f%�.i���iN�_66��7�,�pM���ut& �% �pZ���/p���n)��c
P���n�ݸ�G�^d��رc�b��7�g�+�3H��>���o�y��%��J��@o�^	���5e��X�iPrX�@��bD��:��I�S2A�7��h�{��$2dE:�$���<�ߖ�%i�[S�B��g��#���ZO蝝;w�l�{2b�^�Q�**��\��/Q�*�%�K^S�C* �'�$NNN98�e��T.���o�.x.��_�AI��:-��PVT٘a{������X"-=���"~յ�u?�#���-���������d�.cۖ��ŋ�v��vw��fl�%�nЁDJ �Ǣ>�.��Xb��k`ځ�&��l&ր��`m��ҥK8�q��׼q�F�"Zrtl�!Ц���o������wdm<�o�q�ܹ�e��p��G��4������ߑvcjs3b�k�fMX�c�x�����X��V�BèV�,��jeD�eq���(���t[~�-�fD�(�aS`�@��㩦�7�uV'�4�i����7��e�C*`�j�J��"�#��力B��_Q��޼��fP6Dh�,2���\}��y�ã%�Von�v>%�F,nX6�"xA&J�am�����5!/�!����I$R͖S*��8�t��phh$K\�t����˗/C'��M����츸 �e2��6���T������I�����E��\���\�N��(��6�Mx�a�k�Z(�چ�$��}��-���W�{�*ڪƀ��u���C��8�0~���Z�D:�����5}���~p5,NH�F�	1�}z�J$N|�����=^�L���ٳx�04�F�c�xo6֏�C#BL�Oxv�6�rl��G��:�r�q{Gk۩��2�v�ORS7�V�SW�֪UNˍ�1lK���:�N�����l9ɤ<o���n1m7;�9.�1~'�����j�o_T<P��\>�T�Aũ�L�wo���T� B7���jjhLg9T���d`�F�M�Ģ�H��iM5�2Y���n�8��J]��҉�*'��_XX�9p�!�7�5ܝ��u�u[��9��t�������P��Ƈ�o�� ����h��sҹ�D��}�κJK�?P�j(.Φ��7�ڷ}M��P��fa�+2C܄������?�oݜ�C	�nπ����bA'�C���z��H/%6��z�R���[�է�v��O>�p��������������Ց����|���:u���h���t��W;j� a��3���)�j�����W���'8z���f�nٲ�0�IPq��Z�0�a��.Ǘ��/B��
Z(�Y�$}�����VO_/d����֭[ye�?y��H��K��y������L2M+�Wz�� =���Y�ʻ�F���m���d,[�?����l�#v% ܵ�!K+`C��R��[Ԓ�G�iB�Y	�D��q�w������ʩS��޽���੮,�H�lhw�w�������?����Zx�k���cAi�g��"n��@C"�� ޕ����f.ەI�N�<Y�(��J͉�K���!02�<3s�$6qa��l�c��ܹ7w�NG��<	�;�d����ލZ0]]ݭ�7�GNa%T�af�p�ܠ��.��Dŝ���Π���H��ȯ��"�Cr��J�p����E�)/W���Cv�Y�nkx%�OL�QFbvX�+�-�#f�#C�q��Ho������/�],�C塟<$�;��M��δ~����/X�c__���e�}�3`�&�CFc�o��15�d��d��K�h�IY���%�t���@���k�����h�Cww/�=�����[(���fZ��t$&|y��ܚHNt�p#�z\�� _� �^��2�5����L`I��^Z����	��g=~b"~��I�|+b��xv��J�O��"�>�8^�̎����S�:h��Z]��穃�8������Ra�>�t�2V5{~T�7�<������.�D�ȃ��w�wG�>���̓�n�ٱ��K�$DYj�*,��K.�߽}G�;���4:���A�*�XR 5"�<k5���&���H�
��i�,���r;��V�˸�J���I$@�5:��uj�N{�����w�do޼Irtt"򊒊�z��O<�B`l6��O?e�P�⅗*��̢�4�
jz�vP��3�y'��j���~�VV�ra��.����8\� ��=�H2��˞`��`ٮ�nn)�匣q�I�W,�
F)�q��cXCwN�gM�s˖2p���1퇶�� ~4:đo�~�չL��w����R)MLL�_�����~��o|ceYz���g{&O˴u�b� 㖎��#�����<��/?h�N���85�Qr�Q�S:���[��¨�A�D��ex��nJ� �еk�p#�2O�8�h"!k�(3ٖ�D�K�G����Y�/ �έ3~Ki��V�}F&³ڶ��'�W@�پ�uN��3�/`�''�H-Ja�0�"7�
T�L&⽠��\�j����|q��)��	���:x^�7E��x��	��u��.x<DV��	;�A��|F;D�ئ�v�l k޳g�����ׯi%.���q�F�w�����;(!s��O���v8J1h�d����Xf]e.��0���u|llT�f:!=�ɼ���nj�CFfi�3�������>�ɑ�ҩ�nk~\P{~��_B<���ؙRM\e�m|t|~~�}����K��۾��`��Ua،�%g"���@i����b��U'�O�|pHePG>ť������v'�i�]\pdldia���O��hjRD�il�ggq���Vp�-X^#d����=-]��gm��T"E.����δF�_��|IG����ԈX�t�������W2<�`�Ouy-���MN<��'�E"6��5�t�f�B��k6Ll3�wR�f��Zrކ���ޒ��C;���q7����ڹlzT�l��hg���S�ݨJMڝ,Q�r��p����RRe_,W3��s�fn]��W?}����Y7��_�����%��.��_�q%����.ܟ� ��������q8�)�yǎ{ꩃPw�݄���kZ���;������?�쳻�`J'e�u�
�ˆ�n��� ��9�Ё���>��/�s�����BU�55�mmmrP�$,ӕj����gөI�RSI$�9��%�ە��Y�����ᡱ����:O<��dv�{�������"Q���_~��OO���d=����ޅ�%�X|�xbbl|aaqll���;CSS[>��c,ojj*�k����L���fޖӈD����Źեy<��=c��їS�R8��rq�$a�zs��\���L~yq%��V��(���+M�@�,E�}�e������� �T@�Ր\^�T�>;J̤��-M�
k�r%��ЬC}��U6=�9|�Kd҃
0��4MS�$�dz岔Q�~�ͤ���2V�ҪU�����uӈ�uƱ.-����۸v�:������͛�j�k{2CFt��m�dG���ʁ]�&G�`[�
)M'�^��W�7��'&�M?�^�����y��[���k�с|O�ʕ+��bh6��\�x�U�pp�۷ݽ}�RZ����	q��l6�J�2��綋��d"���\)�e�q4"�g�:�|�D�h{1[�H0�G�o�&�M��$ӀZ��о}Ӱ5�u��7�qf2�����=�e��)G`ǫŪӂ��V����^~��\���[�n���c�����[��m���;3ӛ�2�m�ft�罄��������gϟ��9|�48�^�-����r!�K4����%�#i{��zITiqD���G*�J_�;���:s�z�Z��7����ҙ���0/�}j�$��LK��aT��m�JF-���8�R<��-;���TG���і�ajk�LY�M���z����Iۖg�qn3��������@��\��W�hĢYË�9��8	�!��"R��Y�(IM�i/��%1O�؟�ƚ�j&) %�ׂ��n�l���Z�`�VUQ�lW��Da[�S8�AV���>��m���Z�`�T43�wo�F_��gG*�w�aq)�Ij'4c�i;��!-؅�T~ۭ�[ؽ�I�#í�gN%�����[�V$�MᐬՍ��� $^�.�G2�u�w�;8wgΎ�wZo4��L��j��݅��]G_�:�`������hL��2iЏm�'���@*���*[ӎ���J���;PXY�yMs��(�O��	�_pn�܁��f
�%bPv�����/����}���?{wabb2�z��������IMa��f�-պ��9IDԫ�Xfnv��矿zE�l�'���n;��tF�%��T��z�f�N�Y{(�͚�&�@�)�8��c�1m�\���V�x����u�6h����Nz�۠
7�A}�r�ބ�Ib��x� ��}�J��1�]��M�Β�H�UZ)!qj��\�r�^K �Bl�m�a�;6�z�G���f���;�����yA\�rI���y��R5�0EҴ_&e�e������޿��Ӊ�͙���������~0��i�R�E4���=��I��dwr]��w���"[u� L��b584MG��V[dk�`�́nK�����Y|Et�+��p���s�N��F��kk8j7cU`�ӧOo۶�XP���� U|�	7}���w��D}�6�����"z�X�p� n��X�	A���!�k�1���HDvn(��\4͂�K������~��*��&4�ѣG9R��(�T6�87�T`DG��R��,r�� ){�ʕ�ݻ�y�y��p���i�����ai66d��ܐ�ܐ�8<��'�O�W�|��֭[�c�E�5)��?� ���c��He�[������E�)�.��������C�i����J�:�Bl�6���c�<UT�E<MrI(��t�i���b��`y�S}
;�$d�ed���Zbٖ���	�Ca�� ��so��������?��{��?��A�D�g�&�&St2���Ў��'��,���2�Á�ōu������ʆ�87&���g�0I#��
��3;���������1E��Z4M�t�
!����i`��Eu��)�Ι��b^x��I�Z#�� �a��x5���R�Цb:� ײ����~S��f�f ���vS+%L%oOq�>��?~|vv��ű0�jEq��f%���|>GNc�a�,,xl��M��_�e����D�����j:t��ŋ�eݎ;�߸Q��K7�k�	��nl&29���|V��f�>���l�֖���k��S�
��(ky���u���R4u��v����`�22\�Yo0�G�Hi����c[�y/x���ߧ|�ڵ����׾v��M�d��Gp�n�"�l&��[����{g5�p�f�2.�% �E飲�r�X�U������SXX�����a���0� ��z�W�>'N�����g0iY-+�	�ޕ�W����C���p±`d�,{��س�(��ܿ�ҋf"a��g.W�����ZەӍji"(�ݔ-��m���+���(�oH$[M�O>��#zO�8aGD��0eC�vGiᲹ9�3#����?�1K�ވ`�Z�k͇:O{Ny�� �SV�{�f� �m������		|�B3�c�&��yA�2�'�@��9�z��п��w@�?���t�r)��Q��F��2&.�-�R�g�nW.υ:�["���
�uE͘�-4$&�\�-�K
�,������w�ː�h�>99KƠ�X�L�wܚh��-�:[��J����9�k�J;s�><x�`�ZR<�
s�&5����w��Mvc����d�<,cffw��`�A_r���ZY�.�ߦ����2�좼�*7����!5�����Ǟ{��ե�ޑAW��`��������?�opt}��R(������;�x�$=쇐�֕U9��V*�@7t�\�Z�EE�DI��v���U1,6�/y�f����L�� �6�W�R�T�D�L��dUb�#�ڨ� ��ၘD��f�R��v�6�®c|������T�p
�Z��}s��֜�2ƞ�+�T2C��?80�G��m苗��f�o!�aG���ݸq�JBj�td�.	_�88�w�����R��6�\�~��a��ߐ׭qp����z����wq@���O�m�>M$t��WdR���D�]Y�'0�C�������Y�H�چ I��GlS�{kڔ�C_�m��*�
(!�K��\x�N3�5�R�E��##C x_��3��\*��לt2��כ�e3�T4jG!�၁��5���U��E�P�)2!
�)�Z��d"�[�
m�c��0���^{�щIP`*��Gb������0������v�^�����Aq��MRu��d����N_�8���߁a�Z��gLSJ,G��\����͵z����sss����Z�k�>L&#:P�.�|�vT)�w�W%��& /�N�F�L���Dm��T��jKEM�����`?�`�cL$㚁��R�Z��X7���j+K˭ ��I�_��V,BQ��j�����|N� �Հ����X�f�� *�<<M��"˅�8�?��?|��g��`g������3ݲ����n; 3!�}��=�V��5i���8�pBp`�~��G?z���0����~+����������W^~1��mK���۷�:��.�V�`K���27]�)���.��U��e�����_�jlbϾ��z��%p�AW_?�䅴�Y�{C������;oϞ=�<������u]}}N��j;�L��[t����."�}4&��TJ6�]3,���M�LY ��#�+(�V�b;�4�O��i����G�m^��r/�M�a8��}	�ɇ���訕6>��C�ɗ2��%0I���h���� O˽�B~��;�Yx}G���j� �XB�:u�`(*�4�km8D:+�4���o�a�$��m(�V0�W����ؽ{��k3��Vn)�S�e=���EvB�H�x�%�Q�. P�����'�'�;����4�(]okkrG��������҄e�B+C;����<	j���;wJK׈��L���T�ww�0�������0��,������'�pn�5Zj#��ư���<<<�˩4��҇��{0ء#Gf�_��将{���$�%mٲ��#t�s�F=���a*:������W����Y�Bڣ���^,3
~dȷ��q�$�i�20�Ԫv�������-��X3ĵ���Pu�c�g���U{�nhJ�T�X˃}�>�6Ĵ��k5X"��S��HolR��L.��!�DA?TZ�����@�8)-����`|���8�5X�^��.�&5�F8u�^����[O��T�o�Qg��e3a�U�H�m�a���v����v���待���t��Fr����2kݶn�
^�:/J{�x,xj��ں}�QE�u����-9���$Ĝ/+�L�l�rS��=��R^�j��.���Il��+���~��_��#('�Q�x$e[�	�O���x�V0�"�fCi�"��}xG��3�ځ�8����*3���e�J!��1�j�����&�!��*Z3,��_ju�">�b��۸)��T�j�D� A\"*�+aTz8�ID��0|~$�B[$�a��:Ή����Dq�sy�u'���P8�����ϟǙ�ڵ�u��I֐ʮ�n��֭۰�^����$�KX8H�DE"��Am��O�28���i'��ã��o�t�����c�A����-��b������_|�Q����t��[oIB�q�)�2.��%��J_�d��V��իP��&����ۿ�����VTKl�0��.�p@��p��F _\<,h��{����/�/���z���Ǐ�i���wr�.�*q�	�:)3d���ek�o���؊OK�?�`�J^��f<h�l.5pu�$$V�?�ŷ	l2�ͺa��hS
�{��~x+�O3Q�W�����v0�T�O�p�y+�	��Ria|�����I����+'bmK�����,q�D` ������n���\v�S|:5�eR�~+˸��˗�	�t6#���|�Ne�<�,��������� ~%S�xN�㉔����X��g�:Zh�$N�I	 E>�k�+�Ջ:����R��J���\m�g�c^�j��O���㆐���|�1\��?�#^�#M����j���̩��#G�Tk���ݽ��^*��� �lZ5���\�p�тi.���N�s��O�p*�U����Z��#a!�9M��U|`H
)�RTI/Ć��{��O�v��i��S&&���I�k�Tu�@�F;�O7��[�R�J�H�ٍ;���l+������!���K�*%����̀�Οfk$�6�oF{s���h��h�F��e��B���j�W*6VN�1G�b��X �[oT#Z��РK�@s�
 ����.(��
�֕�F�������!䣢_J�, ��d������L��T}�7`����iN*I�ԙSD%h5t�B�Ha"w����3��a�*AoӴ�]O���1E�f��x�G!m���r���R\p��X*��p�0�zz����{s���7�]E�V�a��Q�uw�n0Cո1s���[��u�Rn� ��p=��H��U�3$IB��D���痖W�7�����S�{ｍ�u"2(EN+��)E<�͠/�?7'St��e�ODd�������j!���(D?�4/�6<*1Rm�i��dQ�0�ä���d��z��&S�H� ��2i��+f܋�P�IhJ�s�G���X"�Q���4N���uf�ʂ������~z�ŗp��F�V�$��aH�K�I��!�.Cҭ�B!K�S�t�DGQ� $yݪ[��fgc
$m>/�������Ș�rޒ� ������m]�2(tҬ	"nwW�ٸ�� �J�p'l���бcǠ�>��Cٽd�Ѫ��j[�H�i%-�Uc����!��s���L����['ƛ����b�\l7M���}����k��{v�r�m�����'́0�	����R��_������s���Ci�]\^���X\��L�t6�C��)m��i��/��߿??7���K�.�(�-��2���;ҢT4�ݻw'�1�!؏+wn�ޱ%I"��@�� �v��ɠC�ʇ���h�T��_@���> ����_ �]*�\EG#�+3��+gpt�,5��3������<��R����R�7#���L7�b5g�?��Om@�t�o�V���51�ɀ�g3"�4h�lJf�5���������km�c�t�v�1FY@X0)z{��h�AdH��^�Gl�Klܐvw��khQٳA��������	w[�(�]׀{9�?nm5���h#x�孯���I�6[ť�����K&{��#���X?Ds��H=I�n�
����O��Y^Y�vA^��9R-��Q�N:����a�t�JO��9e-C�`��j0;;44 �魷)��q��:t�I�NA*a'ar�WTGbӋ�Yu��۷N��q�N��=�w�x��W�i�(
�`yu�����ݯl)haTǘ�=����"��`f�㱈Gb9��rXy�b����ي�mn�W���5��a����@�l/��;*zj�;�I��bM�A=Ҟ$}�H8�O{�����E��b'a����<�* N�'S����k� �:v��?���Le�6�Yߝ�F�r���8��1�ytZnP��;���*֫���'�>�㴍 -���}�������$tHN/�1�ކF���P�'O��V�X�Y��El�=ط-`guDG��}gu��O	B���B:���������$��/�����������JG��	�������9��"�qB��=`�>��x�޾*2��$�Ҁq��ɤ!�F�@�RO�:����)E%.˚��_� �Ǻ�A��L!*N�#���hC�����n~-�i��nԉ%�tm6���\����Rb-�n+X�ۖP�k��C���E��m�!�V
gԨJ�����,w������뿾���S���v횽=#���E��˖qB�;�����0���$��X0������P����~�i0�?/ �а��ȷ��),�Ū�����y�6L�yc�����w�^��˿������7�����������\� �v)��\y�yA�d����B�[��0_z�tV�)a��;ɴ�!C��&^ha�b���9A��y�AmX�劷m�t��	bŐ����f䦑$�3����r��i�)������8|��X���ҥl�/C�I(�3DhS����r�#&�����'�FH��w|a�~<b��K/L�����m9��E-�a���:��{�N����Y������hԚ7B���*ٛ�xR�%:�fе�+*4XN=l�\d�Vz������;����W�"����}P���Oȼ�;wh�M�H���{��8�r)b[�j�Ѭo�����%v�#�\2�`�?���ޑ 5�H"��p���ːt���q����Ͻt�=���p�,�	�������Hk�)��re�^�Eb®D�3,��<80�g�u�/^��c�v��������{��ض �K�.������d*�؂����������u�(<~�h}��j���<7Z��������j�.��Z�,�h$4 =���L��w�H�-�����Ŧ�m�~�Z"�裏Ğ0퉉1\;_�
�iDX;�O$z�[���Lk�{���2
YX���35 `�����
�W��R�AJ�hk���U��NY,d4�!9�҉����9�����hJ��%POqXG���b��]���RP�՞J��N�}J�֬��kk�X�C��-!��[/`xx߇$���Ϫ�����9��m@Æ�q�Ɓ�6�&|���n�vuC�Co�m�FJ��6���:�ƙg�Fu<I	*��T�%�����d(�M��6�m�J^	��V���	_�GE�� ��-�/���V�jG�Ӓ�풾�o��˷�*����#/0#�^�~���wNW��rq���2��X����b�8cې<v�W?��V,���2��X2�LF��O~�h���n2��i�FF۞��%Z��G�z�ɦ3�j��R)�#��� �d<��34%�)Z��7�:�%��6����T��u>��\? ~P��
�{���z���ӷ���O�P�����9��}�=ո�G�`�dr��1�B�<|�Pw�`���-)So���S����Q�C{�7��5���4	Y�`tR���ɕ�^���V$�j�,WIW�p���[m;��L:y��iZ�}]�0#`aL��ų�V�r}������+H���
����u<KNm8�|-���q��k�;����kk�ǖ�V��36��3ݟ���~�'�XKc�m�-��F��bBF�k�|6�'>�Tz�ُ��ҹs������Ƈ��~�9C���vw���#5�`�"$x����"N�Q.U �����@��4�]��q�6V>��l>�%��<}�ZOON�(wВ�td�/�g8L�פ�m���)�̊]"!�|��j��=�q�7Ɇ8-3R��~[��uK�9����C��|S,L��
Et�4�?|�~��������&$����j/��.�'	I#�}����՟=~A�3� {6�`��1'�aCu�`X�v�3Z�ɇ��d�����e>��$���X��>[u(�i�yAO��%�,�T�$���qcc�2����A�p�;v�;wNnі���~v'1\/턵���k(*X?�6pA�Q���-�
�|tH^飌�8�#�`��`dB������)�!�����M�p�bI5�)TnK���Q��`K�&E�c��lY���������h���ￏ��ݳÊ��^���-R'w}F�q�5��^�HJ�346��s���?��� ���'�E�1LR��a�+�7iOs�,	����8U�Ϟ=pc���]Y+��59�r6��8�µtF
�!�!�0�0�dti,���c=
	X�]�˂�Ϫ)�{+a��+Mp>�b"��j���Ӟ)(�dBڗ�V�΃�K�hNNNj!v�]�0X���9�,�Ȇ8�8k*�g�y&�lش� s"69.��w�؁��O�F����?�c����������t����ҖPt&���e�(��lF�+�c`��H$a�"G��,���U����<���\"�(�`q�T8Nod���H�֭[�v�����,E�q�i�bc�^�v����o}�[P�� eP?�j*55��%�`R!VKO�HQbp
l��j�����̙3/��"�&q�l����{��,;y�����oѷ�h"ּ�T��/�~ݤ�gy��?@ϡ�z�a �\�h"���O�gQh�{
�3	괴玄Ǣl���3Y�08����/y�^Pi�G7|@����x��\]�*�6KDD����b�g!��
��
���CYm�9F��#mm2,��#Ш��\,_��b�E����p���ė��D�p��[7�<�쳠@��?��?e!)���W��?a��|^,�0���޾>( ���2����S�T���V]��%�2x�!�e^E����㯯��
�
����~��_>����{�dJ�}O�K��K��Mq��v��[�Dm@Dc�,�<r��+�xU2B%�X�?k�r��ѧ/�P�4a�I�t�v�܉��b����}:->��Xh�7GO|]q
�����L��Ti^���*( ����>���V���-����XK���?@+�dM������r-��0b��Cy�DY�YG�M\M�m�լ,Hg��u�4�8��|(�m���$C��n[��m+j�hN%��@o_*���e�*e�KA���f�mwTlC��jj@��Kɘ��FQ�n�rB{�9�sG�VMe��f���3��	g�(���9�FV�L��I�z:�g�n0�|��nޜy�ݷ=������ F�9u�4��T��m~[�,�a���H����Np�Z����͛7��]�=�m�{��]yB��!qwVtr&R�ު�*�D�O�eV�+.�z�d_{�%h��������\�6�}��ɩHT���D�Gc�v�	V�<O�0����Z�g?�����mzǶ�[�JmY�x���詧������?!�x�WV
׮��,�)ތ$��Q�ų�
�C��+k��/]��{���^�x����6�J� ������DfO/�g�B���&��z�Z]
Z�-1e�)�h4%��Vz�w������N�+�x�����?`
9�o>2s�w}���f�C`S���9�z+��i�466ƊF|�-�<�Ν۵F��
}2����T)4horRz*Aۻw��i>:6�=�쳓�C�(v	�k!(g�,~�,���ￏ��ԃt&jn"�u�(���[�a18462�Z�5>2L�O���Jr*W:�=ҋ�TTh�����W�O���_��x��-1�"M��Ӫ�D\hLJÜ�T�Q4	�B�ob�u�E2���Y��JU
�_������c#C7�_�w����>I%b�O?���
����a���*�$a%��P�1mG��tD�&ض+fK<۴d�������|�������o�
}y��E�7���Ă�G¶a����`7ꕑѡz��I��6��X��/�8�ei���be�yTN��_V�|J�vLz�����<�8�ym�:�����䖅�kD䑊xMɔ6�]�ۦ�8G^��������[��AWd~�_�&,K-��DO�$��"x���}�����^S�67�ǐ�gO��Wk����JE,3���g�"���y`����I�u�uH���С�{w����\�<7'ؓ؁���\Wr����N��kǴז�l����cR�%-����]j����p�րG��������z��0���%�2bK�\�u1��������k0�>��ӈiml:LO_�����z��[�k����x�\ɥ3ׯ\u[N�(>���� �_��[��q��x�L�6�F2K����{{[г0����$�O����������#պ���J�و�;�?�&-�!�{|l� ���CC��eK?~v����5*d��J����y00k�R�H��uE�[����]'��m'���UP@����H&әd�Vc�2�VN��@�!G<�Ml">WYF�F���hGNX�d���S�ك�N���P=hJ�!⭱�
MK�q�Fi�x�($|"݇a!���n���|����AF�F�$�6�$�iߔ���1/C�?��3�M��x<N0��np�������A'��aa���ؘ�i���L�!`������=��!(H���Çi~�{�;�������*�ݸ��(L�~�s3�e��3��|��b��:�u��`	P3���"8���v{mU�腵iM�XT.����cǎ�ɟ�	ȹ�PO`]������g����SةT���g�|*���6������V���8������ ��m۶�֜*�X t<���Y"�pC���|�� ,[Ѣ-�3E�Ebqį�Y��y��H"�r+�&�klг��4� �d+����9��U�}I}�۾:S�N0���I����cǰ���-"Œ�����	�w*�K4�"!��.8���w�ٶmzϞ=��H�T�jE��B=��Oº��2x�x}0ڸf"q��7��	�;2�֧�aW�IS����Yq�i5%`�M��nM��C��3"��4-�i��f��_a�_¹gs��V�5�~�*d|#��o��Qk ����,�U��g�$)<���k�^��7����X�EiW��'v����v�H����*{a��q�����ƍ�196���2	�'b���U�'P���أ>ҚF��1G�xYI
����� ���r����Ԣq�v�U#L#�'K��W.�b#ŵ��)�!kE86T��P_���F���#��#/07"�`���(�����P�G�2�X��gk��r���b�+9�r��{:���jUʔ-iE��mh w�n�0�
���$���y�d�!X�2V�Efˋk ����Z�ņF�3�R1��kH���!�L}tw!��x\TPn�n��DtHN����Ͽ������w(d��͗a��^��b�[�̳ٶ}4]&�饗���.�g��:��p(��Y��Td������Ex�,��b�wwW�E<c4������D�G%�O��
�[L���V&�����i7�U��	ZT�M<u��B�!tQBk��D�{n�V��J��#	,0��ƴ��tȺ������^�{�,Y��~��P�<4t3�*�h����`��T�>EpH4T�3�?��4b��.�e��}�@���ٲ�A�J��O�S�����ڕZ��3iMn���1��n5!ᡊ9ED�LN�HN������mS�X��'���9��(������R��u�2bL'�?����WN�:��𿾞^!,�=}��=qn���+��HG��=+(��4H�Rs�O���;wb5�r���%��㽀�K�s�~ey�w���z����]�W�����p���~:
AK�����Nܛ��^eW�d��kj<5��x$��4A�G�X)��Pk �2Y ��$b��΁m����-!�*԰��.[.�Q��DM���ښg[p���e��O�X�"���8uriQ>�_����Q��KѸ�����;*Z�]U׷ϔ�#�NqK�9ЬW�.4�R��ii��4d�N��q�r���b�w����B���P/8�:[��CC�%�=�F�TV�[� �,��T'�kź[�A�7H9�1p\� ���Bt�8�K�.�p��-�ZMB�2����9�CZw��j�e�Ȩ@���@	
�<�QX�y}f�����i
�1���'�Q�䏈i`xn5�ti��t�(��o�)�I�I����&(�M#���F�VF�r&�����|��^<sm7��"1FL���~��� ?}��%��իWEN�m.u!m�z_�-������~��r�+=�ѽ�������ǟ�H6�&�����P>(T�����J��f���8�Z+s����$�*��`5:��M�C?��2�οjNdLI��!cvMe��@�	Dz�+{��#��HH"-�`s��T����򹜧~5��z�Rkxǎl%��奥�2oR�cH�y�t��f^��<��ш�4#Z�RoT��C����#`�t �����|�͕�uSg���Q�Y�3툖��A,�<���=f�X���R��m�lZ�׶�5��J��#��^*u�������w��V���T"�NB�W���&���lܻ/xr�� �T&i���r�ej��}�㛰�lD��Z'
�" i�0s�Ft���>�$� ����S�����wu5���o�}��ȇd,
�.��IXu�#C���ҥE���kDc+��!@<;2���Ҍ\,�#'��[.���y�K�c��&$�??w_��=���O�?|"Ŕ�x͖��nȞ������Xh��}�ɓ��5>N�ͨi�ЪP����护ڬ��i	��7�z>�)���v�0����2���/�6�ov��6� �=���_f�/F�`~*�߰��ۄ!q̠�*�;K���5�vn��b��y�l2��Z�08����9n6�p���3�����/��g���w��yI��<p �d����$�u�ޟ��XYY��s?p�J	�����?���K������С'ACgN�>w�\ae	ǥ`*FiC�ӧ +�FH^���3�)2v��ДKЄޮn�i�����Le\D�$�U,�\��-pm�iq]C����>ͱ��*�C&v�֙a�"����g�+߶m���p�޾k�l̸$���"�
���Xˀ-<���ܵkׁ�}�k_��`W��	lF��h֘��q�(rJ���&��$�i���hh�4Hי��R���bNt�� z�f���T���Dq�_�p~Ǎ���|����	�Q<ç��xR%Q��)�e�p`yA�%�e�+�����&_tJU9� ���)�˰0�ݛ;|���'K�� ��=���ŋ�m�xo߾�a���0,$�Ղ��$6�l\�}�DH����n��Nz�*�v�L�
n�nC��v=�d�$���Hi��g�m ��(��)��l���+P����K8:݄r�f%h������žI-`*J{�W.\��*���^���X&���z���������2D�O'j��7�x�ڕ���	���Ĭ	Cb�8�XF�8e�@���Qv�SBv*�+��QH���_`�K���<?n.ƇD�"x��  �����CnS[,�f�6�3�����k�����?�j6M�'l�e:�5Id�56�����\�N�La���x.��������X��XJ��ZC���@�o;$z�x���%�h��N��2�D�#�K~^ZX���g�]�Om���ٙR�/�8t�]�. 6Qi��r��d�D�u2lh�~��gs7gf�����w?x�ן}��� ���q S�Q�Z�3�4b��O��?��??�̳2=E�1-���I
9�G��O0x����72}Lv�	�C�P�G(\M�\Bf{n�=��"6KB���]Ʒĥ,W��i#��W�b��_���ܛ�ϰ��š�bAg��U>���hD�\K�[�N`4d+0<�t�	Ù+F�%���J�&��9��suJ�������=T���6
��ٳ� ��s��AtM�3�X�_�f�Q�S�nӀ$�X�^����NP?Uj�$�!A6'�p�p����J$�R14�A;O�o�t�����
k; �4Y�]]!d %#V~�յmz��ɓ �C�A�I8�޽{���]h��~����΀�M�U��ضu��g��G#������'|�AiV���؈���p����"ЦΤ��'
����Va(� rC�aw��D �%�pay	��y�W�cĖ~�b����Y�YS:k���d:�v���,~%z�V�˦�6��0�lՈ/]H��>�dhSK����F4�O2��s��G��o�x����'��'X����z��ZpIL�3���F��;��W_����qm���8qB*�O�JH��u��Xb�J��錔��[.k�I����������:��� ��ki��+6}�\�k�6OC�h��4��wyu0�f^Km�-T 8־�H�fc^&�)��7��۷G���ɦb��jaן�/�|&���(&'-T�'�kvV��A�̴�תE�� �rx9�	���:`nn�9Q�k�����pF�Յ>8�f1'
\
V�� ]�1�g��F�m�T��_v��I|��i��~h���� ,'9S�+�?�ԌOC�=�QT;>�
�d�=��2�U��S�4<��/=�������~���|����f�Ie%肓���&֥�b���vT|���S��ҩnI�6�:;6���/a���j~Y�N5�/c?)��@�D�]R=�q�4�|�.'l��/A�tk~�svSS�Y��Ng�Z���ɾ��0,��R�ԙs  ə�b��ؕX��۳��3�.#te�y�Z��	�J�Y����K]`2%���N�yq��D_I���p�tpxQ}����ܭ7����n�y����-�%��Cp��J��0Dm�@Y;P(X���44h �}6��q��癙k=�]c�R���h�`��_��$�Z����0��q���ky҂f����Ү!i0 8R�笅�SSV�n�-�l{m�ڐ�EQ�z���fD1 !��ܹS�Uq蹮<�4���ҥr����ޞ�ވ!��8� ;��_�?;{~��3�?�쓵�Up.n$u����5O�O�W*���zY�:��sZ'-8���aG�޽�����)�š�=Pk�m���>�x�O�̴ޮ�i��G�M�=?.��V䆌�3Y� :X[\�d�F�؇�u�����-#��jvt�e������{/@V��ף�g�ä�T�|mZl���z��9��|]�?�=/B�ڊ��?m#C#qE�Y��m���2���&���LS�Y��.b���֦i��t���XE���aw�I]*܈��~{px�d�+x���HO���R2��!VSZB05fg�*l����紲�Յ�g`���9;��� <c��Pa�a;@\�,@��
��-�w|d��?�w���}�ߴ̈ �޽	{Ѵ�XX.�s��ծ�AȠd:�fWu(�N���V��j��	�hH�*�k��7�8p�T�\B9�O?�1��Mc�|�e�,��U�x�;�ϟ��d.�6N2���cb�V(+��~"�N�4!3S�����ŭ�JSbz���6�<Z�D�Q	���E��K]^|Fƚظ���bF��B�>/X�,J��i}�������A�$m'��|����?� 'K¿�=ly��0"RdX�^4����0��3���}�{cccۦwbC8)kddL�Nn߆��jɱ�(�q�_,�'d�gђ�gff@o��5�U�C�-�MS��A�VZ|�vG5�WR��h�}Mim����Iܴ6:�Ѓ���9;e���(��b0Y-`�~����|�0���`�{w�1K�۰�� �'hƠ1K� 	HQ��� (�Q)<��vF��P����m����BbhcD�Jf0Ը[ ۺقG8�f�F�<c��_��`o+�����4�-f���U����R��_��ȡ8h�
ߩ��v�4�́q��_���ѣ,�pߑ�c,*?����j���m� �D7@��_b{�'!0�W����X���{��m^�P��P�7�j�&�_.i��2X��}�f��l����������ݵs\|�tM�(��,�>�:{����P�zZ���d�2t�eU-�	r�f���	Ew7.r�ĉw�},�KK��`�K�M�f�(1n���ԙ"�-;mY�-� v"�H��U|m���s�X���]�+x�eHͫ���G?�v���wg���@�cK��J��ۦ`�6�x#���\���PX� �Set����}�C
T�4���L*Ԋd��6�Z�Z^;�j��VSW�
oݜ�s$�l�x�EZ�$��j��|�3N�7:�s����'89ʌ�a��Nݑ�+r#Y�	�΅2sO��'��$��B\r���m��28FKe4?���S���� Vj��}��ͱk��3��)��E�pa�����d[�B�?�7�x�-��]�l8���I�[�D��}cFj*�^x���O=0� Ǘ��6����{���}�c㸲�as�s��<u��z��Y�0�14U�	mA����������<��T���(h ;����={��I��J����|���g��sdg�ؘ��=�ƍ?m	��>�?2��V�r����p�Y�$������R�����D8�D��xu���U&� h�y�ĉ˗/��j����cs��#G�`��$9:���aQ�1��D�
Wt���������^F���O�r
[�MC�SӋԆ�O'��r")r$����5��ݝ��q������mō����@qM,;�rG�?�I�PۍMKsm�+y���Tڢ!�O��=B<)T�ܬ�e�e��`������3�v7��3�L�A|��pҺ���C�����q5	g2�<�E洨�'S�`����'(Q��~a;G��|93{ۥ�x��r��c�Y7F��(�m�Uwҟ�/��;cf�D��G͎8��?�#��[��+���<����1O�Hb��˨�%z��U�&0�.	����>;�� zm��KV릚ǲeP:�%�E9s�l6ZimTj֛^ԫV*���F`��=�(!m/
�3�j���DH:�VP��t~�w��L&����D<ڒ�8{�����|U2��uع/��3�h�ŉ��[;>6��"��	�:�M��7�M]uy��N�T�7�X+ 7pMV�Od�lh�Y��a6£��p�����^,����e����o~��'����^{���C�ϫT*�hӳ�R�W�'�b?r��'�IMNm���wu��0����@_?���GF�am���TL�\�-�b���'�D$oU굖?K*.�{;*�0M�f-�G����6��ݻ�0"�/^�$r��M�ZT��,���|���W8Z�Bamxljt|2�U��ݩܵ�W���뇸�C���F{�U*o�%3s�� �~뭟��g��N<��SP%��ʪ�c�	k*�md��A��R��4V�
��"�����	����$үx��(i1�N��y��5H'P,Y6
yA`��BY� ��!Hx�&l��P�&��ڪi[FG6�fG������}���G������Ojj��~��]�F�i�u 1s��^fP�i9�vc�X䡝���`�� وc�t�
܀���_3�3�����2�H̶ˑg~}P.�D���{a_$c�ʺM�w�X����@,���'@������Ǉw�܃���~�m��b� �q׮],���l9M�+�1\�3�r�W�����z�
���7�i��$�B;���q>�K(IjL#���Z�
oq~�:L�Q��^(@�.-s�"�.��La*�l9x��;Ｓk�N��,V8Fiyv�l���Vx�5���u�~�~CL�\��ل��.]݃"��V�n�.�ø�~2�K%`�`�;3��h*3L/]Ɩ�Q�����eܝ�Eqǩh]3��c�p�[ã�,�Te; o�{��>��M|��B��Om��G�ch�y��-®��"���t"��=s�iSj]OE}�9�yQ�5��\�б��l�NDy���9,����y�p���?��Wc�+�8,��U�ßpL���ӧ,����k��ַ`����?��������Z�-�cc"��/\��ٳdF�7"�1����95�E�����j$Z�v )F�Y��e���b��Z��+sh����$�G���:C�F8�S�xQ[��QK답\�����H�D�AdX�҇��j�ac���s�6T�,)r�Фd��V0z�6h�n��q���N�iX}�p�'����P�:�HZbw�8|�04���lNb��G���WE3:�3�wdɦ�H�����S�JX^*?~|�il#���c����?��:��:��w4��$�Iq)�Z(ɲ-ɲ�$�_�J�y�䌝�3�O29g�s�29N��d�|�$�$z����6��(.")n����@���U5߽��� )Gr�IG��Fw�_���Yrs�x�,���A\��)ZR]*���T�Ma+n��r�D�ɑJ���
�7��_��֯?��4<��d��J����T���9��/��2f�.��,���'l��D����������HNxj��]�����G>G�@��K��T��r�u
��� ßpGK���"R=, !�O�8q��A��2m.�.xnf0D�$d.�q`�l�>-�����q)*2���r�;��N �+��S�8�0���pq|D�D���/�}�eT�Θt���DO]�p�h����TL��R�����p���Z2	���,�'6����2� /��*O�Si��Xw�%��R9��J���2�V��c��Q$�l�l��ⲿ1v`y���'Ԭ2�X�����U.�`�dK��37���έB�∢����,n�V4��%F��[g�p���`����8�`( ������08�O U�\��Ly#�:W��AC�$4�)QY��Ϭhm����1PRe����,8���KTP,ħ�_��_�@F�i�ZCb�"��˽��}�ȡm�7nZ�15������z4H�:�����;s�Lɰ>��c�;�")wu��|��ܹs�<�PQK���z�(���b��(	�D����@�D06KV���X�|:J���q�f쟑5._�v���i�i���E���������H[�B�J(�U5�֭]���|}}�.tE�U��W�b@�Ϝ~3��imnhn�[�n����/�N�G#��x�U"3z�]��x�Ε�4����G@�'N���'�w��Y���P�2�禦�*���OJ�Rclp0�B�c���BUs̮�UyS�X���Lra������33S�[		�Ds�"�ĉ�@��f3�����U؊\2	����ݟ欫D�=��X,FM}M.E�)X*>�MR��˦����V�kA�Ԫ/�5�5��i��k	~�R%cE�'���
�Ca�}4-�L���C>75�������q���Z9���c�8e����f�``����V��
XU���w�����dcG��_����o�~{dr�eŊXepb���̥�\���Ҁz~.S�S�r:ō��?�8���!ߦ�6%;R��k(a����VTP��T(��>S��	�Eu:4�@��;a3=�H,����Qc���'�Z�^���^��|b���N)�#����n������)�%h%է4�&1,7-�%Eׂ��VTd��߇��M_�@D���Pȇr�h^��?���ɔPd��ԬL1����8n]�J���aE������o�i<��r���	6�΄�����H����}x/�0�PW����E��� ��E:��^Eu�/����e���������t��,ZvP�+��mj�`��JM,p��q��u+�S�����'��U]YY*�o\X�O����a!C�Bmkl�īkdT�L�ZU]���A���⍫}}�F80?� �0(���$°$� 7WQ�l��D�qa��.0}e*B�3XE����L/D!�������CS��d&VC�>-h�P�>�P�9�C�� ��!!�8,�޴qme$88p�cu�#�2M�߾����\8�k��#�O����D�Z��b������b[�m��K�3sQ�`-Õd��z&[LP�F���v�b*��۴y��z\�韝��3��vjv�#����UQ��OF#���g0�EXD�U��t�nM�ς��"L͡���~���X������݋�޽������dj����)�V2���]�v�"����}���u�|F��Lz~EGK�*a�������E�+��B�ڣqB�m
+��߸q������[�s�,�66p���پRQ�_"VC���˄���%M��J�P/�Ё�����WM����N�r��6�ߋΒ����BV�!��jV>��X��(~ŀ�QT�R����*�N���.⑹���7�1��������,�*dx��n����\�=@�݄5Ŝ�w磻 �����3^h�<@�(�(���=�Y���T��v/Q�,�a��L�@��U@+�v�F�(����RA'�n���S�z�R��'n����Ǜ��@�p&�\�"��6��=���������9iH��<���Ç�S|�\[�<w�D=��8^�2��;C��_��{�g�֭0Sμ����0�u\�#R���9����?�W�����^c��D" �wk�X�q���o����"����f�r����,	Vr���ק�KX|�~Ӧݻw߸qW�viG�Z��^��kג(��!�${H}4|�x��|�#���k��:���L�Ka�����(h>A�ό�w�[�6۸%�М�.�D��[�$�	�r"��BBpFO�>���(uTX���*�[�2�W~ӗ��җ8��CdM�d|�0O�'�88���VI/�!�8	�H8�F�9��E���95�J˺�P��*%n-Y�!��\�@x��،LjW\5/cv�RD�a�I��:k_������
�@9	�9���c�S���/ϋ��xI6���.B�yC�E��$�o*N۵�2�Kr�=
�i!Ǧa%�g�3�,�M�\<'�u��  ��IDAT�T�A��(�o�4?�W�\����)�rñ��.(�����I{��y����Oh(����&d�90�)N�k��ՂzH���?W��H\J# �4�*���Uk�	�X��τxL[�k�|+��XO�!�E���9u�ԃ>�M��"�3'�*A(�?އ�,��)v�x������)�8�ǭ\����###�{��k�����=�W��u`��S�$�j"F�i�>'�]�$�X�1D��q��h#��Iw$.�@:U%����g�y�ڰ~����}W.	,<hueg�Vp��?@yp(,�.�+v��_�"�}l��9rdhh{�Vpy�"�Ĺ�ۦ�n�x�G?�]|�J�mh�e�"4L�UȑNd�K�w��T�Id�+|~�a���ď)�`Y-Ei�h	k� ��r�ZR���徹Z=*aT<Hu�^���g���Hz��R��B���L^J��LV�$4����D�K3�7G�m��ٳ�<��}����J������^�R$kh��J�8���n��+�~�ܝApܬb%	K�_Q����T��_�
��ѹ�СC�a#(�W^�g��Gl�k+��N��Q��穧�����]i��ę��?|��'�M��:�j��/��P���j�"B����_)����O�իW�\��i�ʟ��t�)��	S��4\@F֐�T�",L�G�|MU.c�˩�y�h6%#��HJb{9��%5*�҈�/_z���Z�H�+Wb��djrrrbz�n�ac(���O����G�x���($�p�F����{����B�&���<<F8����>���)��8�Jg�9X���*�B����<Kó�s�9��8��{KE��	�2���]W�¥��s�œଐWg8C�	�^03In��%*�y��C-� �I)�>���?M��ul�ѣGW��'��e� ��8�R	���S�ې/��$-��a+��3���9'2t"uN��4`��7P����p�B��0[�̶WT�f$�@��JAq��p3J�?ǈ��y������3��C!�b[����F��e�0�l�hOF���� �ɭ�T�TIݒ����J��;m�0�U�GeL3�c��,*긝�uF�B�R.�چ{H���fA�yh�pnڴI�C&�vU$����� �����.��,ح���QR|:�S�S��kr����h����Ď���|���J� O�|`&`�����Ib̒��Q�Be�|,M���Є��F#�*�d�=�h��M�FR
/ u�P���N����Z]2M��F��02Ff`����2F4y� �Q��]#�	�� K�$,������VR�%�ɧ~��o;�JNM�oظ.�M��߄�O�ۊ����}�{�	���TV,�����0�Ϯ]�V�ZU][s����7��Cn"�I�ZV�Ya��ё���W��>�t�����a���hPr��1V��:G�d�A��S4<
�`�}�Pd�����m۶|>�z��9�}�����IzZ��`�pp�P[�n���Z����%�$�R����P��iS��6�0T$�+��D������g"$�E��I	w��-�T\��Rʢ�*ch�Շ~�r�%�>�����.����P]�[�r�����*n����'T.ӭ�f�[6��d�SkѼ�x�W�����ͺ$����t��ۈޥ�r�qQ.�"Oe|v_��1�X�H��hq���T����!���m�ϸ2F,9���N�<`"�����޾n�:i�Qx0�Gz�A�o��L��۷K�ġ1��
�*�~{�~����g��ayLiׂ��wߝ�o��*��(Q � ~��Up&������Mʼ?���D���9e0��iL���B�474
�S ij�� ���q�3+��T����0�����`��?���/����c�>u��E%U#0��5�W�D�ukΞ=���~�Z��؍M۶]�x��^�U�:nJLBaSL����y�0����V��4k	aJs����y�F�'C�ͣ���%S�j�}���hI� uJю\N(�g�T�0���V�Z�%�ǰ��Ұ�V���Xa6Mù��N��3sIj%��l'uK(L�'�c:	Z§��޴)��u�v^X�&n���g2i��au��je<�&ꭈ��q�ᨐ�zV;��(k^͙ ����}B����{���n���7���=<�r;:͒S�/����A2~!��T!���2�����4~v�m��8�߲)�>�/��ق�-�E�5�BD�E�����HR
���3�ob���P�Ei|����n`�L�� ���N�G���RF�Bf���k�"�83�R%-+
[J]�!�U�?!<�
��o: j�w���D��+%�X�˲�g�n�Y��7�Ca��-[����U�
Up�u����bÂ��_��4�#�l���dU,G������7nW������zdd�������XXH��0�D�lc�;w�狐�u��]{�n��'O����?�L�'��NML���?��:ک�g۞=؋�Zꔇ~��7�ۿ�f�
� 2�Bqc�Xl/лw��򗿌����'�xf�W��^xbߢ:'�@�mإ���o|�k�<���M�:�ty f[[���7��L��UI5��~�HNN!�x�D���
��JL ��LE���������"1JIq����n~�.K�Y�� i��$ل$L����j�)g��[���U~M۫l���د�Z���EΖ��@�-���ʪۈd�%�L:HD��e�T˷�[��*Q�BN��-UϊN��N���a�b�Ub�r��!HF"�bA�2�?�P�WW�\�x��#�>z�w���
���̾}��zZ���9s����k&Ek��w����"���F!��`���*W�?��X����4?G��[Zw޶}���@���taI��'�a�CT�w����X���h29����f�؞��9�_Jf���~��O� <�Lo������/x���|���[��+p0$��YQA�C~����?���{��MM-21���#���!���9�����?�jw
D��x�U(@L�"]]]�l�ġ���Ec�am3bgL���!��gg� ���qU�<��I��ΡA�A.]��I��R��`]��l���\�U/�G"Kyg��9Q�b�R�k����(W����^���y�C�{f��5㬱᭭m�W�����B:������{~v��Qt�d��YƘA1@���N0��A�G׳�,��:zqO%ȕ�yIL����1��Y�F$n��e|�OwZ+x�d���7|p��H�*��9%גX��"y���D��Q*7�*\,+�R��d��J|?1��fg��h�C�T��q�����V&�3�f8��������`���έ-����,
��'qp?��u�6���4oۺ�ak����|��P�g7/�Ʒ���~7V���H!��1b�ͪX���\�Uu����.�C���P�ia��eE]���.�
�������$I��Ք�+�g�\���)�!H�䉑�S%Q�ؘ*��K��f	���Z
2?��d��,�$*�g��wlr* %ҳiC1��Ħ��L.���x��෦�zlu�]}�xU���;����'�Ν;�D7�i�S$Dy������)��z���(�Ӕ.Z	��h�x�#����o.��>�����a���_��pVWGg'6FLMMEMEӱ�o�|��+Vl޸	�~�֞�vB+u��vtt�NZVP�6M��fx�U���-$o�@���_�uEEe�Hm��>�,�6��s�.�w�'����,��d{G[mS��/�����\&���=6zC�,���klnri�i�����N��c��&���,��93�O�j�$o����d(v*8C!����ӄ(�a��.Ƈ��\���#�Fr�V�Y�
ɂ̱'��\G�x�e,)�b"\����JF�o�*.�ԛr�}�]5����pO-[����މ�ե��v�Kqu��TQIdK>�fܒ�z���5Q?�R,Ro?���(�"7��c1p�Y4eآ�dO={IX����D�ar�4�]����{��v�ڵu��cǎ�}�П�(��C����g� �R�f����7���j�]��E�t�?��� ~�oV{^f֤ʥ���&��px	,��P/�x_ sJ�%���j�`���*u�X'��-����V9�~���{���k��	���w�����$���k�O�8��o޼YJS={O[
2h������]\lj&��6�_��������Po�!UD$*�}�G��Av���T�,�5�t�f<�X*�ľ'�R���M�ӧ������-�?���<�G ��`<�O��,cϞ^&�I�r0�^��D�V����"R�b�=��;�r媵k���y�?�iؙg.��=W��$���0�O������k��F
.���$!)��,��],1g�!{�2�A�9|��l7<!�;�'E��z���u^�}�PȲpHRM9��� |zq,�hE-�l&PK��ON��tB9b�&SƓ{r���6(^�K��(X��`����� y�\����2���&&o?%je�Uh7=�- ���k�jX�/��-ݣ0���[���:��*+W�Z�"Z�M2Z���u��_�y*%�Z['�'`��/u4�$�DW7-�t�����J!�m���$bA�H#ѭO��^916|������ѩY������	�o��l�W�����Z���n�����3���k���{��Whnj��}ض�Y�HzCB���T�)b:00@m�9�k�B���>��ϟ:q�o�_2B��T"�Hr���e-ޑ��sCÐ�?�0�j�===7n���s.�`?A<2��R���M�?�8�fܢ���z�ѣG%et��!�����[���7^:{�o��oab
�.vX�<l��ui�߯1�5�n+,.T*j��3&٨�x��')��&�Tas���Gi�+P4X������+ÈG#<����Z�<�<-Fb�RahCKqc�r�Bf(����o��\�Ž� �����)c�}�R �ו���'ܮ:`j�Mu	��⟼�PmY���r��DySj�_^Gq�Fn����%�I��ܲ�µK���-p���e#��������D P!�U��!,��^=���=���r��j|'�++�M���CQ�iJ���?�۟���j����w�d��O�#����o�ɩ��/�1A!��J$�1��|�@�PI�K�d	k*������^S����8�.�Sڅ�=�Ul��eyT�MhR�iX4:�N>v����?3̯���~�4D]kjmͥ�tll��'@��X��5:2�I�l�c�;�-=�����|:�cpuGGH������@[k+� �?u�v#V��H�{��7�[��k��c�5����<�6	e�Y���2h�ۙ
��Uu���9�ԕ�v�Xů4?��,�g=9�+��4��RP���n��]�O�.�p��-�z��/�a��H�K�B�t�ʰ��ʷ����s0	*S���U�h�Y6��#
�Q mf�H0T
�*bÃ7|*%�̢��d��-�Q�m�� +�"(��'%d�!?�Jl�t_U,��܁$��T�gq�C8���z��yUU�#g�US倫\�-���GLs���-D$~�%;֍ob�in����p�y�]�Le%�O沥�%�e����՜]PYg�J$\A�7Y�[�U%���Я�{7�Q�W{%Z*)?OW�=����{�b��:?�s�0��؋����	���66M���ڱkg���Ԟ��ޛ������Z��/KH:$�=���T�%5$+h�orvzRH(����T}�yWta�id3�Z��TWh�����O���*�&��2�ꚚT6�/��/k7o�m��U���ht|z�,�K|#I��Q
�,�{}vf��/C�;���T���gsݧ���K8&)	pD�����y
�0t�J����{���?1�/�kj�|���6}�/��"�~c�ҕ�0����9�?H�xUB �Z�!�aWՐ����GN��4K��^VtuWī`������߼evv����C���?�裛z6��X�*=7��s�A�ٳ��o��U�ھC����-�����'O��P__��KU@.�����+�ϜK!O��da���6�y�%�p���s����42l*�4y��]�1:���Ӥ>�\.��Y��w�R)����}�T��o���S�b�^C�`�Ȗ7q�^�Z_nϸ?���2f�o�a�wE{'���}f��ыQ�x��@}�5
�w��f��Z2R�.+�QO�*�E"�$��i51�k�hhf:J�{}R�%�K��8^l�{!4Q�4@������~"���N	H�)�14r�ƍ��Q��=x�ҥ3'Onپ�����yw蕗�B+@Yv�F����E6�L�$22���t���;�я~���\�xI����]@�X��;v:��>	o9g��T�d�M9ٹ�$g*��E�����ދ�<�Q�v�ڵ~��hM�i�R�����,Fp&���+���@�֚�ԅ�:d��[��	K�_x�<ށ���~뷰�4Ḣ��v�2b���2T�t}n~�r"�Pػ�ҧ��Be��|�Ot?Ә���V�Љ�g�ǭqe������h	�AR�>Asw0��W�q�4��.�9h���2>��I��Xs;��� �E*0�)�9�x�C�� R�腊qA�GXu1�$�#���=���˴��I�ز�;u��DJ.�3�#��s��J�L��|]V�T�К�-'k�����2��{�.�gAtR,��r��*����-����n�
�Xºx��gz�rjfɑ`��u���=���I��x-�II�oB�4�ܹSPL%(.2D/	���e��=���*5�^���nȁ����S�MC�x�����e����ȇ>�����
�O�z�D�mIJQ�T�4=#,��xF"!j"��l�")iq�#�.����e`��2���A>��72���f��8}^�ސ��GOE((E2T����6��X�l&�R��?A�45�VlB�ǣ<���#5<s��������:���'O�)���/4���}�$��a�f�;�r��Z?ooo�sA&�S�z�7�������R�M�Ά��uMMu�������� �BJd|���a��B�.���nذᮻ��>���Ky̽w�պr�Ǡ5�f�ĖY��%TBE�Τh;P��2�OMBY�C��E�;K�l(�^�L�q)~a���p�&Y/^�[eq���B��+T���05�I�]�gf��T��7����.�UV[%U�~�y'�Zn�I�D���7��ޥI�f\.�I����+����@ZT��{�=�ϕG�&��@O�r�bީS&�=���Lg�DT��3o/�v��Ͱ��v���
ε��A��
E+�P:ˣX�4���~�eB�RT2�	��������p�p�+�._�|i���{�cd��#,u|�&�R}8Lݑ�/p�С��+��D]m��u�z뭉�i�q.O��Z�`%dP�"�#k�`�u�,��&��+ۇ�FCы�.�2Y�m0Q��@�L�~�#��^�o_�:t D�~.3����
t�H4"b�)RS����x@����|�'�f"=�&0X�N���55?_�s�����@{����OȆ�ţ=��X����N��.��Ç��7����At��������&@�AG�����?�ꫯ�_8G��Q]��P������b1O�5>�{��I�_2�����I.�4�`(� �,�R��
Ǩ�8YQ��N��L�ぱ1'�'��$�%0	����^il���`���]r˴Ի�R,�d�]+�_*m%�	Ч��fxzL �3�F��DSC��ӧyH�O|G�X�Qt�\L];�J��Y_�H�]����)ɾI[�d�%?�3�U5&�)d,EFl(�ۜ9��x!I�;,jّN/C?Ջ�e��?�j4KM%�D��ΆYIw��@՛��|0����Ӂ���r.���Ϧf�*X(�Q\Ɗ'*��A�����[��eg������������Fcd.��!��EH��>���]�H ���G�A]�tR>��JQ���ٓ=�6� ����wk:�?�>Y����;ͧe�
�1�I���oж�3�A+q\rLcuȰ#ٔ�)>p�޽�<Ƈ���ݶsWs[{C}�L��.�m�m�Jx���(��T�\5j��qc|$���4�rՑ��\̐W]�hn�i�P׈�*����ƕϾ}��sg�l7S�0��e�D����������︭&Q�K/�PZ��@�cc٠�c�!uan>"�k�Q����B!�\�q�@_SK+<XT�z6c�s�Ӑ�x�8��:�$Q]F�ϓ���w_�&���er����z�G�u���a�����?K���7nljj���k׮��]�n-D%d{[G;�������Fq�]� �0�nSO��up�/�^޷oߧ?�)������%���8P�d��1��645}�(������������b���?�����f�/�����d���c3LRK�l>��"��6��~�?�����j[&$�x����7��S8Ń@�pֹZ?��|NwW�X��
7�Pʶ�_��J�W�A��
�_�%��e�E���(��1֞%���4K���j�^s��;�oy�\�8f�;��W'2崛8����o�����Z��y����7�ʃpl:���o��F(bl ��$���ae=R#% d��(���d�2MF�,(p��3���gEK�m�#7��q�	z���	f�7��ͯ���$Ή�'�@�Î� �~����]��<w�8jEw�`�Ш�D��A�	󳥱�[hN&��b8�)̸���:41�#s]�枭�ckk;3�́ja2B��]�*S�����$d851�pu�g3f���2WX�8+� �2�� ���Պ߯��{$_x��ǎ����rb�bm�w��Z��ѣ��?<3�|~~�����'��ƞ}��m۶A���ߚ���3��Tco������������8���V��(�Wy�hn:S%l)"�NOE�nH�U�P�&j�u���v�Ӝ%��l�� KY�@�7������~��`���!uT���`4�n��b �)� �8L"��������m����Q\@�8B
&8�#�jr�[�!�%HLi�:��_�r]�O�6R\��,����^
�@�%K�iB��PJm��u����%�V"5:Oج��s��r�����?��ݿl����T��UH{+s����	.�H�$]0l�O�K�fFd[��5L��e�IW8篹�/R����Ɣ\��{�b{�S@��;�N*�N9��������m���K���m/(����#�i�s�=`mJ����_�/	z��7:6)�\�����r�a_h�EET6(�����`���$!x	�b.��,���`��"��u(�裎�X,���E��˓�cl��\��Qj��Y�E4q���v�����!�p�k�ml6�)O���2P�r�k͚lz���Cr/^�+��I��Y�q�6	gЂ���>*]�R]#�Y���g��?��O�~�i���n�M*t��18�\�+#��,x����?���4V��H[��g�ܩ ���^�x^d�bffjxx���.Z]}���<�W�35p���J�!��8�_8�;BI{��rFd�Hf�	���fA�`n��ؼY"o9ĳ�럂�� �?6Bq�ʣ���&���FQ�t'�
�y��e�-��.�oG�I@I��,1j��a�*�~'������|9��=�3ū��n�y�1h8����F���3x��RnT2���}�,��2ܗ��.�]�Sf�n١/��x}�?7B���QJ�d�9�͜�J��VU�%�{^1�<�X����`�]�v����i�5U����o�������=��0�u5�VvA"Hd��9;t��;���{��������w��ݟx
&<�p4�/٪_���Z(�6�P���nn~6XY�l���zvݾ����{��R.�c��`(�uۊ��1������s������ON�~��k�w�y'd"�c�F�
�hE�`�r�p#<M��" ��m���|&[US�Z�0l�%Pqplt�ȑ#��֦֮��Du���������(����T6��ю��W_}[�����nÆ��z��bf�ɃJ<9���̥��~ؗ|�)��@�x��	\���a%/�m�5�8tpNmdt�(9�=e�}��!�%Q�|.%KuE�ټ���?�����u�hsJ���b������Nۻ��)N!&=��ex@Q��B6�e�M��p7n�p���\���)za�K��qt�>���
Z��5��d���<�O��rd��E�i3����h�ˊ�tő֧�X$)������2C3�XVqp��De**�gԃg�#��^"Pn��/C}l�_�R���tw"���%��2]�%�:��Ň#�
�-�OAn���&�U�5�ɉ�l����%�#�*b�luq]g��Z�J��[I��bI�E�v�J(ªD�Ass�Ν;ҙ���deK)��q��oa��ѯ��|�et��)�K�l�q2Zѹ��o3��Ϡ��occ���WϞ>K�Rm�z�Js����)����UUq�V� �t���k�kԑZ��+���3VN�A��c2�/�@�8��GB�R6��(�!'!P������e������/��h��������~�G>��C�_,Yj,
ӑ
gg�S>����4����/�����]���lhjĕaܬZ���������;��l���Vu_����TvFQ�H��T"U%�C�6�����7m�m�������wܹ��c�l������B�Bl�X�����[�l�������Ӎ����
&F&ĜD"���=�g�g0�^?�Zww75�JEU|x��b0��k���`'�+�B�n�7n���Q��O=y�z����K<WƶJ>]�Kf(����M��oH'h�h&�1�2��$�*�(�_RU���������j��(��r���e�V�-ʈ�b�R1�u�w7өqɡ��#b�<L�P,��Ђ�ZŖK��'��Y�D�%�o��_o��;;�1�,'��yե�}�����x_�9'w��K��*k)� �J̈́��E.�����xP&�pfJz�q����5
ж@���z�;뤢$�A�WXE��޽{!j_y��T���سg�Zh��\�v��>wM���LOO�ck׮�>8 �j�{�z���c��?���KW`�g��p�(/��Q�#��e��?�p}SS6��ք�R$�li[A�
ц^UWg���X̱�o��ih����?��3Ͼ��K[7o�!%F��N��$��tX��Cr��p��܍7��J)��P:���i1�e�)6^����O���J����2����2ة4��n§<��k.\��l6��GG��gHڗ�I�G��R;w���٢�dJ�L��q��)��A�EW}�"�!",�C��jeBYN_��P�d�)Δ!�S��ʈ���yS��<��c�^n�-��_W�~�����x��3x憍���w��I�#���{����vt�-2 (�ȵ#R� �M��T��
�LNNʞdi��c���iz�rB�������'!1��^�(!���HU�͍�r9�Iȑl��;�Ѽ������$K����`ss�I����zQ
	�~�WP�`p�H:[��,FL]W���1�D ��GSEjt�j�wn�Nc
;$R'�in��(��k��U�9�[b�KZ�INA�1�
o���0H������!��9�q��Z L-O.�QR�a2�=DDV���fp���e�!�5���A���^aj���b	�0EC�禅5��Szy�BzG�zf3�sۣG�~�s���?��ݻw?~���˰<�-�gh��av���ccc����a����+�����6n�o�o~�/���M�� �@�s�'~����V`����������78��[�q�`I?�4��i���;�{z�H�p�}�A�wt�T�h���b.G`�`:�5����nݺDU4u�q�F�������?�����ڑ7Ξ=[[Kү"D���
��W�{F!T���f8���/ƙ���>��"� U	�~6�%���0
R����d���QU^�_��P�w��ۇ�i�P���/�k��U��˗4���=�M�(������������e}���!]	Z��&���N�;o����+,M��W�z=/N.����J�S$��*���n�����zD��E�Q]�ԭ0��F��:n�2X�I��*�Q644HW�mj�����O�����ݸ����Ü���Y��eM��	9�K�ơp���������n�x<@ç�򕯜8�fp/�}���B���M=���B5��5�F6}���a��56�lݦ�>E@F�R�X�2^=91���z��૒���Cm���ַ�7l\OØJ(�,[�l����A@�`"Q)C���mQS�Ku�Y�'FF<88x���{'}dx���Y�om�~�O~�_ ��g��;w�r��)������Z�{յrź��7^?����J�<$u��4��S�N�3!8�1G:�; 8��J��	X������onn���UJ��R��%�%��dIJ~S��5K���K^�X2�&�`��d�Iܐ4�������#�ʭ|,Ov(K��∹)Y!�������`0q�
���ܱn{��0Yi� ���p��D�[��!�0a༺:W�k v)���Vn�4�~]u`+NO7��d��>��<��#��ƨ���G�����D���$���@�,@��{����N[��|�/Ӓ�>��;F���e�!��<�`��O�|�l�@r����_���g>��ԩ30�E[K�����O�3��,�	@NM��+�ƹO+��s�|���z�����I@�H1�<F¾U���z�Ԇ��5�O��=7/�k��PE���U�|�\abjvrz�M�����uuuBƦ����8�L��"a��K���"��&�$�%�����H�4&?ī��o�D\��뭭�Iy��obrr����յjpx��
q������IM����b݆#�t&ս�����Ç@��?�g�VgΜ�-���i�I0��_��"	�B1{{/�P;{�")�E��6�Ln߹c!�<�����$��"RI�ǯ`P�UWM�k>���m_����2�������-[�lMmh L8=��":<39Y��;;;��^�vm۶�L6zKK������@�U��w�رc���\���S?4H���\(<����o���\��(n�Z"Ģ�q#X�0��z�)lTSCM��7��Y2ě�?H�K%�W��(���%��F�Q�R�P2�B>b�F���R�HH�4.U�(��ڪL4H:��S�6h��tZx���te��̌)�v��(1�spnAJ���U<��,��>�I</�ꅇl�~�p�#�����X�,��%� ��_ڭ��LK-�^-����x�"���܉�w�<,�g�l���KtBu�	�A�".e�� {�qV,P?#��A_�p�a��$��f1�񁮮.�0�f��O�����O|��?��������z�+V�+z/]V�'n����l�̙3�@肹�����Z�6|��_��~ .�����ׇ��Z���.�x���p�C��/��ܲ�d��Щ	yzb���n��M�CC�,u������ؒ����������7�,���p� {�=HW��kѰ ����?.rcx\���E�r�:<��I���[p��Ԑ�ȠpE�ŕ�V@89r�ȟ��v�bUa�M��*�boo/w$�qMz��Ӄo��`p��4����UR#B��Ţ��[�e�V.�$��_�Q�J9���å�/���
#��&N�� T2�G�'K��	AI���,�<���×}��g��񋢸u�FP���ۼ~�o�A�R ��HhG_���8����r哱%KJ�%���հ��
��g�;����\�m��p����[*�2X�ʃ� C3�h�$������q,&l�Eн���Z���/���I\��!�ATQB:�&��8a�/�� 
`����Iq'�Dz�����p��S|%^�����@ ���*�>P�R)=q
kS�a��pEY.�oݞ�^�G6G����K�-�3�羐��ܱcd�/��|��E��V��N��E�%*�mI�K�h�j�C�H� 8j���
��%R[���&��S-�����/�422�w��]wݵoߝ�8�'%m�h�T+:�]�d��+8�Gy�ĉO<�Ğ={`��(/_�N�j�	�92���8�-���>��5ݠ�o���=~�ӟ��B�Ї?��������}���s�uu�2{�V^Y��O�yLj�p��?�����/@S�����4D����~��c����Ԗ����"�p�S���Ɉ?� �S�Y�^|	��s�N���̌�sc!x��۷�Pv���?��p�M�C\��5�.]��Y�u���c��E���a|��b��*8�w���d�������)R��/L/2T������M�3��U���fl�;P�(�>
�e���t����D=v��\A�*�Qa:��et���Z^e)�׻��kG�3ݻ���R�pF�d�Pe�%��e-U6n0�Qj;υ�Pݜ����*��V��Q��|��u���?�J�侢t�l| ��
<�fBD3I��E���d���\0k�k��I�1ʢ4i��_�������mmmW�����������Iq��诎ֶ���Φ3�d,�u�h�:H��c���")�{��P�ʮ�����:	1q�=����5)�@=Xz*5�+\��{���/��D+W�\�M�p�r$�'�+bV�����چ�����l�Җ�Ǐ776H�	L+OԳi��p%��ͩNT�'�u��L�k��*W.]^�n��͛D�vuv�RF�7�:u��������AXx�Ø�Ɉ�;�F+�k��,�y��_]��R}O=V���s�ׯUũ� ���_�~�3Y�Ñ�@��{�c�A����+ѝ����9nZ�Q�"Ŗx��b�e-��T�y�grqe��M�@DiE��^-�lQ��Q8%E��Z��s�W9?�)tĊ9 	�T6��3�!`��Il#e<����jJ8�R�]*����n�
h��Ҡ�%�0�T� 	�\%�c2$�T�IW�cێ	�H.����E�',�.��@�9�8���8'��@Q�5uw�
OVHO MO]f��Ҕ���-=�{թ��=I��G8�#�N<��>��RX�T�3|�Ç���D�X�N�3	;�]�#���o,\X�4��Y�+��l$�8�h��MP<$��n| y�ŵ�>��Ӫ4J�-U�T@��\�SW��%^x���W���6/,��������V�W]@��c%����G�^��ZI�`nS��X2Gb�Y�w29O�A�B6:|����8hԇ��56T&�#c�Xw,��_��L"�,YPCYט%����h�����L��W^y%��wUد�8�=�х����;w����3�u��p@�=���}�����޸q�[o�5<:�gIT�P\�燹�����9��w���ӧg��`�B�G���T�����~Ϛ��T ��i������X$��ʣ��t�|-x��`��*˨���R��6\��y�f�[�@���j8������<���ph^�̨���@��=��K��fV �q�`
��ż 0	�����͹Q$j�1.�ԫ�^$��V�"�yg��ӆ�T2#�$��.��,�S<�OJX��by U�®)�ר%S����,�K_�R�~ŭ�Y��f��Z�C_���ջ�e�Gv�S�
;^N�@YC���Z(ƬϷ�ͦ�Ft�l'��ĸ[�"���(|��*�nT��Ѝ,��gH!��I�VR��$�|
GT'uݺub�|�_���� F"���==��S����g
�7�:��m����{��^h��.M���=>���j~�H �u�+`<� ����BΙY,o˖-2��"å�~�$�"-�Y��5�"���o,$~��!"��P�ŋ�!�tx̹�y6;J�Q��#P�oj���J%���� ؟ɉi�4/��"��p��z� ���+p��R#C���D�����������#--͐ �V�Z�f,Q���ޮ_�Nܘ��߿?��Φ��d?�gH|�b6q<*�ǍdH<���)���m/'E.2����h�����Fa�U٬�"0'6����9/K1oI�73�gW����zb�a۱�4�JbFG�A��4M��a��� E�⹿O��]�y6|����  �	���c(%}8J;���dU5��)�/��"=ZY�W�'aHɲ)���o��q��'����_�.ȮrW��P�6�2/���2g��-��'�dRF���詭�V(뤀���0Yr�+��yey����v�/}��8�{xA��ϖ0�t֖�h��rqV"�%V� �w���AM�5ȊlŔx3އ����T�"B�-�p�+V���a&2�묪�À 4�L���B�Ѵb��?69��'�d��ٙi\, ����T ���#i��ɸb�
m璐���R�8�����n�28�=�ψ�%��a�� %�v�*��5��b=����}�O~��`��E���{�@L�ٱ¿��/�r�������-����(�;WQ�O+��Fu#���ӧ!0������ƚϝ;�ERc�ؘP�瞫�W�鍐 ����h�� �@9��x\x8y� L.x��7�x��Sy.�
y�c�Y�ݻ��Z\,�+���F\�}'~2� CE�#��d86����ؤ�p����a�G��33�D��iC�U��|�Ii�bv0�l��o�R�T"�K�9ͥ��[��b��FO|K��/��j�eV^q{+��������$���JP}��A����p�ܶ�H��<��I;�b�ō�5ݠ�N����q9�ͽ��/��!��N	^)�ږ�/���C٩��:�t:�,s�]�t��U����lٽc+t|,B�09>Q���9�b�J.n���<�(�Ld�[a,�A��͵���>�/)`�����QUu��54�4���{��Nf�_�/���#�̒r��ɕ]=�<�������[���wv�^�^�e�3�H�$�0B]�U��� }��^����N��F>O K��g`q47PA=l�G}tn>�w}���-*����bVq�+���9��Q�_���O�����l۶���??}T��RÞw��a��=�
Ҡ�"�(�E:�-����Л���sO�������mm-}}��,�G9�������͛6�4��p�̹���у>�HDo��}��5s��n��1
�o������E[k;����L�"�w�]U��o|��/���5�;�9{���c'���&3���1�5(���������xU���� ��<�X�P�tU�A|SkK�m�p�4�n�
#��^)F�A�d�T_0�a9U������Fִ n�s�x�K�T������>e�gf��[��E�X�w�+Q�,�ɉ1� ��L2USE�	zhfb2��h�}O��?�ފ
T)��d�p(`�*����'��e��D������X�"���Д�eF4+�� �T�Xx>_�K��Ժ���FK*Ĺ!zbz�ڨu5��$5�i�������P,1�Kj|r�����,��t�4��2F���UA��ݭ��es��3��}}��d,MWq��t��E#��#F�� ����G�E˜��k��3�b��f�i��t��"F!@م �ղ��h���`�BaFT7����TUͥҫ�w��v�A�S���V,ZN��`��Me�'��j����#
h�ʒ=U�籵��76�޶���)d�q;W��!:��3�bp_����TW�YFpb4ٹ�����B����S�ͥ�R�,��_H����#,��_���U/8�X���8�8R�����t���ح��L�pE8��w@e9H]
��۶l��S��?h�
��a�$��~�/��' �M�n2u���׮9�ڛ/��uk�Ê�@Q�XJD#�h$<t}h�v���r]�w���/��LM|���>���}��+:;q�;�S��f����r~���g���%AHfҍ��o9��s�]���]>O�/�v�zz���|r!_�C>8����g{���>Ȋ�_:�������"���\�t����y��Tuwo|�ȑ���������O�OB~����<4iUe�T,q�G����ЕԨ|�{�c���`(�����B2�)� 3��~b&پ�ce�E�$PH�[�"��2�H8h|:k��5v�
L&5	�*�#��TaT�2�Du&����gda�V�Ra���!�aANMM@��c1YA��4�C�)A�]dH�.�R��R����E@kQ�t0�xhڼN������ZF��ӒHt���M2�|�-���^8΋c�n%�"(��&�-T�A��%�-c�R��-E�35^��7��=��M� �U��E��v {��C�>Jq�9 G��3R�!-`�����.�\�f�@4D�ԍ�Ľ�I�S8�@P�xj8ݖ��%�h�6��Ϛχ+&������/^��
7�رcpA>��`�����|4�ٷo���8�F�����T>�1===�����S�'�<��k��5���|�I| ��`�ᬰ�O~��Z�����F������i��͛6m���,�;=M�.p��Pz���������+_�ti�m[9���ڨ�g>�pq����@`���I�[0°u�CC0���I�Ʌa��^�!Ǉ[��@����Ν;���'')����P������x�/��"�P������� �._����&l�M�6N����ɓ'U�N*�8vx���8�9�_
G�1�8j��C<LόI�	���Y�vF��t�W�w�G�RR#�,�����?�W�_(Q=l��ާha�t����Y{�aiUU��RE%�oɶ��9�m���40}|��; �i�(�xr�L�:rJC��hS��T�l����t���Fɭ�G�3$1-A ��Z^h��e@��5˛৊l��	�_:�l�(�n���P�X:�BZ�C�955<Ρ@,��3�h@Ё2!�l��#����Pq[:���u+��_����$�����WΛ��,��&B-Oi�L:> �����M,9z)R�,�����Z�^Ni���9�H�"�=�ɘ�c.����l?���ҸH ��V���-Ȩ��{�߹-D4�Ģ����'�����/}�K�6���J&鉸L��?��ַ>�ɏ�ɟ����\l|�&\����|�;����+V��g��`|�c��׎;j[����� q���ͮ�n¶����Ç�}w�57?'cα?�>#8d�o��VC}�ʕ+qS�P�5*������*��$T#�y|�{1��u��y��~�����a��f�V5����w��Q�Y�pE����"����$v	Z�{�E�F��X��M�Ar9�0�$��+�8�jI{>�����)ya1:�]-��8��J����2���x񣥸*˾�����!��J����%��sͲ�����y����7����+ed������3%$'U؜�,Hs���0�ޕ���ÂǙ�LAOJ���vCr� 3 H��	�A�%�pR�dZҸB���K�Duu4Fl��JW�P�
L�f��_��P�������w�q���u�eM+;�mX{��VTF�\������ar�#EY�Y*���w�`����[`�g�}���(�u��BLpXy{g�g?�Y�h0�"�����&!g.���5C��y�:����oo߾}��{"�/vsk��
h9���B��6��KT�B�5�S��a9uu�&$�px�޽����*"��!VTtvuYFax���˗��������	�FB`r��
JHlk��Є��v�Z���NT�O����?�����R�W�:�Ô-[6cI�1�i��6lظ~htt�C)����yf$t��f	ɝI���0��.�4��F%�Z2�Kֹ�ha ?\H4�sd�Md������qn�#�z�fp�(מیwJ�Ƒ�ջfM�3�<S��45�Ud%=�_Sݒ�1��p�a\��s~n�ˑ�4(�!7��d:��1,6��x�_ug�X��_%�*�Q�ް�k8����I��.�t�H�'iV�W.+]��?&�y��[��R�3J����C�NN�B��͎@q�ܨ�| ��6��W�ş�xU$Kl���Mŧ9c��eP�� �P�Ճ� wg!�č�_g�,��-�.�����-Wf�n���XLs	����� p�*�yy,��'[*h/T@�/��*�> ���ň�!(��k׮q7@��e��م��ڊk�).�!GMA��42�1e�XJU�HER��Яk��?by���P$��gN��y�C��GO��_��;����㏯[�
ndr!d��F��?{�IP>�GV��C�?�ih`W.���O��Gyd�굩dt�n�H8���`�;v�"��iׯˌ;Hxi��e������}�s���h�r�
�V��i�P�D�64<xcpXtv������{�������G>򑚺ھ���oi�a����A�W&��Q�-fSj������d�)�tfh�]�e��� 7.]���}������Y���|洙=�gAz��@��P8��/Q�k����:���&���D�Rږ%� 9Ͳ��Į؟|��>yK���a�r�L�k�b�4[���I]re�������J@<&����;<��=����8���;�dc3<w��҅f��p���uh��-Kz^xjTr��&��
"@K�5��i!K� a���	�����1T����/A*m�	+��A-Ȍ�U�5lغ��@�M����zj��������>�x�ܺu�r�B���S�N	 {,��Vt��3g�`�'O�y��w�ڳ'@(�T��O~��ѣ�N`-��߂!�u*���i�͡����ӧ�}򓟀Ut�����5��C��q��I�؊D<!.'���+�GM|�u��$�ݾg��ӧ����X�5���lV4���A�I_E[�Y�Qh���c/=�<D�T��MlH8����ۋ��\ٱi�&�hX����a����"<H�P8�^oi2���>,H߃����8�o��I�'���g������:��Lc)�bWD����X����4+|І�Z6�	?S$8�U��ō����~��� ۅσ\q�T ˖���1�ٜ�!��wۈ���R����֤*Q?)���U?�e������K���5�"Le�t��_��C��h�O����=��h��엫.N��&�f�cH�2g{����=�N@e�s�.���e��(5�����	J�%��/�<ؐ*���z@��2R)�g^ϻeݢ2r��}{�,Ҡ�!�%"]%�kE&� ��\+�@�}q*��B��R�(UG�ԩ0h��l�gK��gD�^��&w�zX�Vɐ�'|Rƍ4�S���׶J������%D�H��>���#x�����l�FbH�>�$!8q�֭��;�$0u��ŋ!�6o�,qkA�$j�#V�+H)A��Ҏ�������Q��u�׹�̜^p������-�r�vd��E��87�q����9Y�׍Wnb'V�\[�}�؉lYrQ'%Q")����^@� �A9�ͼo�o���e�q�,-<�3��?����۷��C0�����_x�+Vҭ����g0-x�ӧ��O�No%��E����իW<��<|���+�H�~2����;{�l�ٞU�V�v�m������M�6E
i���V�fD��ʬ��p��kr��bl�|Pe�w�ܪ�'1�݊eΊ:,d�4ԱU_bF;.�1�I-��X�?�υ�&��L��j�ڽ�"c��w��p��o�̻�`�<QG9���2�5���P̓���R�f���z�,-�r������b����=�3��<�Qy6�H
h�sȆ�Y�euq�$�<���IGlv3+���P�X�/P�+X�v�o`P,����氱�Ie0	c�X�
�Eu�ª�W~��_���?�h���ʎ�o�u��9 1S�L�M���3K�H$�F�|&���)�ϱ���֮]�tx-�H�W�XT�����+֭��v����� hҪ��Ϝ9���֔��o���W�ڶmۉS'+#1a��F	q
G��L[��rӗ��Dbmm��t浽�G㱍�7��M�*���H�' "��ի���*��-Xp��I�<��\���[o������@&�+ =C�|���5sfwOWc ���-^ �}{=TD��W^a>��(ž�>�>�S���#�����M1���5��������k��,�6�f��z�L�t$��H>�)��k��e��6b�>Dvq]XfY=�ס��r�Į6�ax�a\,Z��-577B��ٱ<6n�x��Q|.]r�����g��g�#�	�3�?���gϚ�NI�VTSS��(�*f��d��K2X%�&�A2�LJ��G���_b�`N��Ϩ��e��5�vl�X��X�B:ߋv�߄��z��r�ԩ��i3fa?HJ��&5�B��V�e�K>G�:(樈Z�B�pH�I$z����T�r����� ���R��G����KBg�E�=L��m_P�z�S8n`u#��I?{E_pY}���Ӗ�_��ֈ�s+�����_��+
K4Vc���knj�;��/����Ԓ�ד�B*�Z%e%7<�hh�lp�ɦ^��x hْ/&.q�'��B���_����Il��l�N�	�q,=
��E`�e��m�Hi�iT�ҕG�P	��m�Mcc飇ߘ7��w>�ۻ^���c�ҩ��޳��Λ�	�%ۚ���$�HYK��]]����E��Q��G?z���74��G�����_�}i���7�molo��Yx ��*�j^�ȫ��������ɭ�m�^+T��{zz*J��[`���[�Ξ���!>�t�4>\�|y�`���^طo�Ti47��aL�t�K��[�<'�*`˼��w����׾���>c�Ҽ�͵]�S��vH�.Z���"Q��GE���A��cw�W�!_!�-Z)�C1�'���m��L~,�1%M��1��-�M���%a�C}d�&��@�!�]���3&2$j�P8�Ϯ��|�qy���5k��țT LxG���Io���R�} �JJ�v�u�n5u2<UN�J������mm��2����}���G?]�Z�k�Ӄ�ü�H����0�	������ш�0�@&��u��T��\$�����E��˔�� �{�󞇿�- �;v,^�����ظq����-�<,��S�;��;O744������*i���	X�R�O�~�if���|�
������u�O^~�e\ׁq+��_���������$��G|��lܸ���}�/����N���$̓�U��5.�a`�JFZ&��W�Z	ؗH4L�5K��Msx@P#����&jjm�/�&�c�e0:B��K%�"W�c3���Ç=�̶�Iw�u�Ak������Ǹ�wމg�#��_�"��O�gɹ���1Q�,�S��'Z�\?X�Hkɷ��9�=1�4�α�<Z�4�|�&EŢ�Y�5�0+���+�v�F�e���T�r$�Y
*SUr�8�~X����ǅ^+VG�"�P�Di[�u��1� =c��僇�C+���)�B��[�p*&,R�j(��@��~
��O�2���]�E��h���M g��t<�g�'��y��tv���\K��M�BbR���\tq�/`��Bj*1C3�3�dWW��ׯ_��6��OC�o��GT���W���t/��]���C��E�"�[�GoHs��Gbu�?<Zi-�lp���ߛX��U���EMň<6l������$I�-�a4�QF6��.���$ R��d��Qbg�"~��W���}Мd���� ���c������.\���ࡇ��1eɒ%w�q�0SJ����y�7�]�T���ak� �@��1��_q��'�@��f`��3�MRSz{�O�����}﮻>$��,T1D��������
_�����BOnݺuΜ9��e˖J=���b0�&�cT�������o��������Гe��h���)AFi``�oƖ��(�^�X��u�--��~��n��l�E�Q��YЍ�?׭}n����������b��+F�9�</�8 r&L��`�WЪ�ӥv�]C�X��v��Ψ�y.��8��x�\����R�y.���^t�?�/=���	I98,��S�,�(���a�|�(*t
!����k���>
�a�P$�v�ɤ�xA2�z�9~�(�8B~8�N��C�gaZ+��䥳��?�c�H����7���v��/��4����g���g�L�F������z�7u.��s��;���
Y�VO�Fs `x�m۶��u���|��{�����p�%��$�^y%L|������^�͜;'@��|�I��큥駺���H$���u~�s�K}�+_��u�GGg`G�<[5�A!�ǥ��������z���X�����c�$�_�k���rϹ�G��ZO�YL����s=�[�=�Tl��_pp�����<kk[RS��V�Yy�5�B�k `�g���q_����O�E�_�.]�s��8��'O���X���Pm�ꦖf��)�Z�Z��[8�Q�q3��b�&�e{S�2� ޾T(�GbQP��X*��5}�p4º
����cʵjd�tW���/��:7�Ay��N�a�` �� �m�[./�h�͛{�|����MH�w��'�����K	Js542
Mo.�Z"^���p�?��R%�3-�	?)Vb�r=.��9�܊ϣ��*�����6O�������nw���c�`�6�\�
�x�����S�:�q-g��2���X;l�Rڵk��}2�D���"���d����
���$�.Ŝ�%q��q��qA�Z����>�M�����w� "9�T����BPF(��̧�p�SѓeV_�F9xww�ں��\3�mE�D墨MJ��hrxd���^���&R@�`P�C��Rj���ѩ��1�$&A$�S|?�N�9�%n�a���<�2i`�b��*Ѝ*�&!@a��!���\�XRk���L�lOo�$�)���A/�s�R�Ab��̳sYq�uLm�"�������C�']�eSjx���'~����>������*��J���\}}�ԩSO�>�8/���S��g��a���}���pV�8�v$��C#�����:}�x2�z�����z����x��V���@��%,s��03S�
��c�A�Z�mij���^�I�����xM�:�oڴ)�=��#�忭�E�[[4�#�nRHW*b�9��}sdtl�ڵw���+6lĖ�s�N+$�7�����#�.�^{��b��6�}R��'�av��Z���D}X��ڠ%�{�Y�_�'c��8<,���ƒ�Y/�dҥi0�ӵ�=XbT�u���Q:n��+ʓp�+��:��&[�ӻ��ִلf�E�%!J��N�Q퇞1Z����U�TC�fp�(jM>~jM�xX�Ot( �9��C\��GF�T�4"%��.��Xj0�����Pj�GG�K)YL��"��Q�����&q�+������h,$%�b��75�r�-_��W��a	�]{ş�ɟ|���L�
i�����l0'�[��l�����K/�mٲvtL��D0���O<��O�6�t��0N��񲴜 	��n/�(�r�4P��� b=T�P�cr0�搖�e��m꒥�/^�`*�����܀kЌ�=�HHnG����]0�믿�H+@%���p�u	���`�}��_T�>}*�$��w��;v��}'}�M7����}�o��kÆ˖-���w�(���T�N���*a_&%$#,������@-��bf`J�R�p�U�t��l�b���=�Kj�L�#�n��ږ%��p0�
=]�ze�z�.v��K=�<��L��24�c�jăk��T:����g'�@�J��xk����9ڰh$5Ɣ2�����TF|UZi%��uG��duE��Jz��|��e.�)f�2��+27��o�_�Q�hi��+w/��9� b�X��:κ�!��V-̒1�v�ګ}ņ�����K��EX_��z+՗x=���IB0q)y��a�D(̟r���ִ�d�� ���q�SuN��[>��r�i��w��u��	�}6+�3�!ϡB�u�E��.X� =�"��(U��5�#�����Um���a2Ψ՝���x���h3`��ͤ)���b��M^�g(����da�Ŝ0��۷oI��\I��P���=�����������܅��PD�֨ϏEP�̫�\A�B��~�߀9�s�� ��O���.X'�|f����;��߾v�Z��dX x��;�F9���m۶�·Bx��oϝ�aKS�o
z�|��e w�����׾Շgd�,X�HI�G
@���5�>�Ϭٴ9�ߏ���w��
�۷ÓͅӬ1��|�;��ꁁ5�'0�gΜ2�rQ�G��gX�nkgkS���4�=p�%�?�>���%)�~7��r���<0S[% k̙ N]`�z�.ux�hk���v;�ѹ03�R�������u���`��^D��c��_zL��K�d�3W0�]3�%�Η�m��F�!Q�c[&�E�,`mHg�H���E�
`��r�rH����&Itg}D���)��������T:�?aahh5䷂���lc �=����w��ګ��M�a������?�ac}#���mc�+@��� �4��*
h9w� �<G� �mmm�> +��χ.ۺu+[t��v��5�|�r�WC;@�p�F�Ǿ����ʕ+p)m��Cjμy��[$?<��g�#�)H�~���������Y���S,`�j~X��I�2�@�$�E�FC��z��x�ٳgC�B�Ϟ:�t�L,�~��W>��{���	甋R��� QG�M�]�u�}��V�\��O}�g��;�sybL�s�=�W^yÀ��Oj[�|��p�b�����ħtLË�:��C>C�Ų���R9W�kl����R�X*r�[�z�4��" �t_1;�����	�7�����/>�~�na2��9"'�f
���c��o��~�ȑ��)~a��BPi��fe�T��Z_ߠ5eS%��ݮ��`�k��3c2`�ri)�`�Rr^"*J	W���`X��¸�J�2��5&�ϛ5c�4�ޡ��h\��XGzP�'�#�&Ec1�̓t��֪0oJ]^4qAU��$��[l ���.�����ٌ�NIֳr�K�x���OIX�:���2��%�t��۔��Ĕ����������א�c������t�眣��
C
��劰�9�m=�*��)T��<����[��W�>ߔ�.L���c���z�g��Y�fA�!������_W�����U3D�`8�F�\�86���R��Dcc�,ۺ���	2D��yc�	j+S�4e*���VO��XBrl�M���������3�'|��ҵ�TSC���e+yr���h:�un�B��;�L�%��̛�su����>Dv�U�oڴ)	gҩ�hZ:%�����Ց��ٮ���C�c�Z��p�₸g�#ǎ1>�����0-@W��KA�c�a��d������]��������8c]A�B7Rwa�PV���d��D_o���
:JX<
�d����6��������կ~À���Ģ�/���-G!�]g��cٲ�����e8VSc�d
��~��5ke�t�(Ηdr�����E�-$s�XǄ��B0c�ojnTN��5h��E����ȫ��M}Y��jN��oK�3.�3�T�d�X8Ě�D����՛ �!)�`GG~I����	����3��6��Ĩ��kz��& ?F�t������z����լfT85��C]�u��횾:<��Y�Y��r�T�'��$*~�h&��aq!G�Y�C1��R����b箓S?
�\�c�L���{�����*�f�!�2�QK�~+����r|V�������|%��_��5��n��,_b�+	��Ǿ�ai2�
�]�h	rg͝�?���8�;c�t�d���3)�&�������5}ⴋ�o���D9z�n��Ud�aw�o�q���0����Jҋ���r��p	����d��勹��c�x(�6Te,$T��dX������kn['�:�^{-mV\�2> G�q��K_�Ҋ��z \<Ň>�!�	�43����GIeh���@�Ɯ`��~�uTaR��ar�5쓕0��7��z��y x�V�����P�, �w�šA=�hǷ�_l� 06L��*=�X�gX�tJ<(�[���XV��Dm�xC����N��B/�)&8�V,W"0����L��[�7cW[cI]gQ��ؽ-�4f>��g9�F紤��+-����Щ	_��~�Z�t�r~0o��ڟ?��u ��*k���UܯL���X
���0Ů�xW]u՜9s \R�����#Yh���z��7hd����k]�\ɞ������<��)��AnB�n����G�OrJ����"�	�i�<l���U��y���k
���0��"�U�ZpͲN>m3�I����.d���^�w+��rj0YV�P�~.��f��q௩�ƙP�xF�)��7f̐4�����w�s�`m9zT�5ᨗOEM~���!.'L3L�����,X��1{��@�����LPz=� &���[oN�b�CBa��
�ؼy3�'�\ƌY�[��	�ٹ���y�����b;�ӏ!�:�#-z�s244��w��^��u�bEp�%��'8�*�Dp��8ae�D(>G�e�J�����˙��q
iHP����<44z��I�_��鼼n�(�6��OXt.�3.h�#�J��Z/4�i�3��3#%����s�%�����q~ZO�K��ת
ȭ-`�W��a]�E�$�����]-�t�����X�ˍs��T�dR)V*��(�q����	�|�\�am�Wa�]a>̗���t��}����'ME�
�BٖV*�H������*�d���<i�MT����_w��aן�ٟm۶��=t���l޸���9�2m*9�8сǞT�`�D]��9e���g�|��{��{��q55��d����k��_4_�����v�ډ����0�t�7���w�ޝ�gpe+��?kᴎiXv6l���b�T&[;v�P��s�w���]{^�?��z���l��)Lf����]z ����ܑt���p��)k�׬Zy����|�;̽�_%��� Q߻w/�
�aӦ��G?z쮻���XG�y�{�,Y��#�<��·<_�u,ガ�'9K�OF�����d����&�a��VM�L$G��H�,dr.0z29��"�
y�b���F`w�I�ዡ�ϳ4��o����5L�Pd/\n�F�@�R!�T��vw�('�8��z�{�옴l&PH}�w�Y�F�EC�� <��� �+m��B���}~E���|��M'�!����&��5��e���N�N���+���O�b�� �]�,�O�{0G��/*��lVhH#��!�d�$�����|��҉�qR���Zx��IQ)��HBﹳ�U����þ��=��[^�=ljj�K���f�!�U�i�?ci��z�?7n�R큨�D����W�IHS�h<�|`T�7b)�O,Hh���� ��>�1y���Ų�·En|�HH?�	�z����\��B!�C\�;�h	��TS(���%7���1��e���)�G���
�$��(�;�M�����`*=<:&D��-�ሿ�I�wO���G�Jc���̟?���EMC���l���Ƶ%KGmx��'���cR�R(��$ ��X���O��R}�WpM ����C�w����t�
�-�y*%�K����.ҧ����ڵ��o��kV��V��t)&j�O�����=>_`��)��t6�j�Kʴ��Pqʆu���s�M��������M-Wĉi���ő\dY�
F�UۑH<����붴6	���c�.	�n!�b=���p�n��G�6����U�w5���%r�T�#�T�]K��v9j����j���6�
��a�&(՗]e�3�����)!�������@���R@�3!�w]��dv������8K�q�1�!يM�6�wF[0it�I
�f1��'c��p����0�ɇ<0��h����v�`��X�OS�<�W�ZxV[�j��4��T�7��}��������}�_\�D��w�qV'����X,�&4p�ָ/���1���$�$��W`�tuuaCŖF���x�G�.�S�$�⇋oٲj�FR���zJ�,�����Ո�k�������M�7��`gŻ(�1������9���>�9C3[_x�%�����ŋ�9sFuJ�~��`��	fr�ڵ��u�"|�'00�jW�iX#��x��E�0��;wb�_s������?�秿��/�x�+V<��s˗/����O�ǁi���N�L�d��Ᾱ��IƔ��N�&����3t��wUl2���x�I�o������o(Ȧ\��k2I	��� ����4����E]$z���M�[�2cd�hT�y׬"����j��dm&���aZ���e� ��^=��7�	�8.�	a��^ny��$������{�7Bn�>˒ڎ���On\���4 �2�s�2EA��o4,��\��<J�p�~ ٳ�S��z���m���:K&B� �$�a8q[�d�=��y�*u��%���h�  ���矻Ti��tzg������s[Vu�z跖��XB5�(R̒fs��H�[�b�-s��_�	�3��.���''/�k��k&�0)�Ts���Z���_|N�Qe�0jvAf|�U�������g
W&����V%k�'�g��_�iX���>�ͳl�J��|s�5�@�=�}�֮Ap��%���6JQfca}�㳤W�]����@-�s���F��0-Xx�`dV[�jգ�>
5���|R�c���5�b�3f���fAj���>+��ia)۸q#�����@f۞�
{~ɢ��+�$����A4I*������gϞu}�}���
RW%)�F��[K�ə��Cv�bQ�F��X�L��pa\�gJ�:n*]ޣ�{��ut(Ƀ#���U�g�k����W�
�*+�Cm�����Q�:����f��bNM���4_|�\`5E?oUR�b��0:�ڹ��y���nBi�}�K�d{NB��喉�8�IԟO��O�R�TmP7幐�����Y=�����ŝjV ފt;����$6*�?_G�%�F�̪�q���7�pQ[Kcs,��+�f��]@B����KZ��_Z� ��>��B���O�yeϡC�������w������̛7c���"I�`m���Z�(�p$X*�n��z��I�ֽt��{��ٸa������Pk֬�ĸBgf���9s c'����`.�o�~��e��/�x�-�-�rlo���I�N���s��)�X�nݺ�Ȁ�LH������7�z�Շ~xʔ�R���	���3�vL�GcO>���3gH>���_ݵc;x耎��XeM.(���-[2u�H�ƃL�<i���7�x����u�H� t
�*��/>���g�2[J.��*I�Xr�$;U�w�!h�|��1yJ@��4�ث��H4ZW�����.c����M�ƨ�u��2����K2��5Cڮ���F���A�ZG�A@�P�k/�إ�g��O���ꫯ}~+���m'O��/�%��W��4ބ)��(��֖v�1���]��;���YJD�5.ņ��3=J<׫�c���T�iсi�v���.f��������Үw�#_��;~ͮ5�58�����t�ٳ�b#I�2�B�X5�c[��{�S�.(��4j��J&�jHDM�t��alZ�~����{��d[K�m�$1GI�K�I��YL�w85��4xRo���B�m1p����Iv�j	7�ƨFB�O�J�����d�B��#�]�����W���Lf�����f3##�@����^���D��J�B_o}]��)��|�HH�N�{~m��;j	�젊�,��>�k�܊�!��`�*+�P��N0dd�g��lr$��e+-�bi�F�PH�3�B��I�X8�.����Db��hq����L������)�~��[�[`
�.�iik��+����Lk?:ǰ�9-���&+��W|l�,ێOJB �g�~
��(a�Z�|�I(�%K�@}A�'�[��ϟ���HK�x�q��Ű{Ɏ�e�pB�����=��S�۸��u�R�v���W �����V�x[0謙��B��_ �qY+�}~i�a[zR\�ɤ�Jҷ,@J,��&�[X,�K�Q�
%�(��\�������@ǈ�%$>�	'!:�5�4eJ�a����~����6�oP.A�_�I�t��*�g1t4'�
T�i�@V�[F&ia�"%I����'���j-�	�|��qg�SS}��eڭx6�78�.�{~:9|� ���1�B(2�k��<9�u/������]
iaRP����}�;��,Db~����FKe��p��0�.X�H��Ҥ\�j���Ř>|���,��t�>���K��3f|����?�cL@E��>�Q��]�vmذAs}r̎g�*��3z>Ȗ��Hy��H��(@
�(<X��X!�k8��}}�W_}u�ֶ�1 �444�w��+������ԩS���@���Fu�9��u��i��. ?��=|�eoH�Pb*��da��E,X�'&����ѱ�A<�Y���/��u�����/^��<���=��ԧ>�G�-��+�P�2�����#�&�T�d)�Okk�Xv�Ⱥ���-���%��0%��nq�$�{ķQ�+�:�#��N�|i�W��%Q�5LX��"��ɎJ���ĵz�6Ro�j������	������u�JR�7܀g߹���ȯ�  ������1 ߓ���aBH�U$0 G�U��i�pH��'�J�S\a�|hķ'���""��b�!~�V�"��YS%p��y���w�1Ù�syթXØ���sZ�&[c�)/��օ�'�p�FL�t,I?�s�}�mڴ���CYШT�	���9{�5j�	�ԞWl��Rc]z��&��wC��l���W��#�#B�?iR��[ۦ1a��Xn�U }�U�����	�R�91E��,��לQf��٢�ή�l����%E'J9]!a�L�b��ֻ����x����K����p�Whni� x��rQ�	�����w�;���������4#YB�s���G�Xb	9s6�)4h�3��5$�Ъ�[��Bq0��z���0{�嗹eH�QM'8q�����!��v�N��i�|��{Ψ�8��=R�~t��bh���ׯ_ņ�x)��佈 �e�P����qG��}�m9�����,	v�z��Yw(9��b&��Sg��)Jw�4���O��>H>L��>��UkU̚c�L~;��1��G����ш�
�K�����r��q)b�X<��g��⛞�օ�z�w���<�Ҩzф�gֆ��Y�q/��{(x���H-��������8,@���<�(^SM�L�ӂ���h4Aִ��d���D�d9�
������x�,��ha*�ԛb�_M�3�\y�ͷ<����ơ�����:gϼ��[W�X���ߏeD�ڈ6~9|���Ia%�c�?~댞m&�B��Ν;k֬7�x��	�0�d��pr���X��$�����;o/W��p�]S߰�0oWXH�g͔�W��|:�6��
i`�7�j��1�IcH������YH,�,��)SJ�0 W��M�ť3c��#|B���-mnide �9�2���`+�iǭ��������{�3�565� ��­�ۂ��؊���g�4���)�d�g����g5 p-ٿpA�:����cL�v�q*S�Քg	@4y/���I�L�D�V���e7�����j��F��oE�rv*�#=/���εkמ8~Js�q�P�� �^�/_96���]�l��-9����֮^��]L" �I((6+�A���tT[��,q+iw2�@^z�z��T�e������,��	�g�	�ׯ�����A��t������LY�0�{7�=���C�,8X#�C=XV��~�>��TjL2�[�.+�-�5��,sD|??gިfE�m5�L�K��/H�ԑ�	ܵH���-�ȩ2V�q`�e�r���X__t[[��@��m`3{z���M�Z�:]������{G�G0�����].f2)��P��4s���+U.6�9U�������8L��JX��'0'�ml��lG}���'�<�7�2����P)���s�T��)�e ��D�^׮]O4���?�9��/~q��-ܳ�U����E��j�TH�fTܶ�R1��"���SV)�����d�B��
ƌ��	������:� )��i�`Ci��P��@p�ꕑX��٧���w��{�.h����r^���C�lf����B���BEc��ϗ��4٢a�mhВmZA(S.�$�c&󯻼��5�`���Q���:�F��A͔��kQ�c�v�4���OXm��vk�����i�>}_'���=�=~�	�
.�}�<����w���75������2خ�'Cna��̉�Ϝ��j0&o��{�9�j/z�u�˔x��Qu�����[�:���J,G�nt���� �a�PA67K���bU���?\Y�*
{�c�I�'��֢͆C�!k*JT+����1�W�	� h���k@]�ui���t�M�^�&E���7�lق�,Z�h׮]��:��P����^O�=���7��x���͛��y�'�}�٣G�buJ���Z�4��P߀�t嚕�ѩS' ���p��G�̜9s�ƍ��ܹ�|�����)��������'�+iyX!�`cJ�sD���y��7e��\:��c���O���[\{�@~���������><W��6l�֟�R8ujСx��e(� \��[n������?���� 
��v^�={4�A��#^������?��\�R�ip�f��}	!KģP����g�����+�-f��ô"�F�F\
%}6������י3����Wө�W|x0�w� ��c�@�!�,�~_LO|�{�+,'{d�J_4N���vR��G_z�%G{3��� b3�� S���8���K�D��L��T<�T����X,LO	.���`�x<@��,Ҧ�M������ �/��P�g0�1@xHerDc�z@���K,f�aĢ҄+�k�����=���'�}�N��?���ːP�d���wꢉ��&s�Χ�-��}�^P۪��I�)�ք��X�6Mቺ��`f����Y�HCm��=�E4ab�]VE��
EVYI]g4�^X��x��Ų�:n&��.r"𰴉-��4ۄ:!hj�J�wYX�ؕAhՁ��>���\����E��p/n+��hB����r_�n���������56�b���gP7�$`	*�`�`-3Y-��1z켌�Nf ���x}�la�����ᯐ��l
�h/Ş���yc�����';^��0�0ϰ�I0���2�_߰a����5��ۺ�ڪC�hfl,V��X���?2ƣ�n��7��A�\<�$�iI����:\3H�,?Ǫ��LP�a~���ĳ�Q����b���O��BQ����̉X�.�+�+<0:)i�3��L�%| ����<���7��ˁ3�M��<����LO���Z��j(�	�1S���&�,lҥRA�?�BH(~W+/B�8蓼�bAB'��s�G�%X*����:VQ
C�9� �`��7�T �`�55���B&�'��腍�+ڦmp8�N/���I� �R�Z��20�"�De\�g�K�5:f���ڒAb�.���ߑD�f�5��G�~�q����s������U[֏��޽�v
����&^^��hLB����D,>wN'�2, �����7o�l�"�=i�����v�������Q�o}�!�!�D�Uvs:�jw��	1��9����H���ĴiӠ2�iI�,V��fL_�N�|C+.}�VI���T�444�<q�>���T�d�����v���y�;[�[����C��(ĐF��!�N���G���	z332���v�ꜷ�4��gO�k���}Sk���}:����3g^kk��sC�t)�_�@2�;��:��g������/�d&3%+*�P����� "�l:��[w��I[Z˥|:�%3J�li�V3Bt>2R�f� �BK��`�X:#Bh3��'.�������*���w5��ኺ��&���)�aUj)�bӒ�M猊Ole?V0�`&3V*�-�_,��ʞW��Y�p��O���=emh:�i�T�6�3��������<�!�"����L��%�e-���U�f�M��M��4շ�4�䳅`�x�J��g(���Oؽ����:�����Y���������/�f���W��ʎ�
V�r���u1!F�z5�[,{�	������B@�:�+�9
�������Œ�:V9[Hm�t�g��˖.:��gZ�\>^'U~m�����烖���y���$�֧�	�G�&�� Z��F5��p����G�O�f�ZO������Z�=#�Ɔ��V���EV ���$tY��+;v64K@`xx(����O"b�g�={��yl,�!c�e&��d��URBS�t,"<�@��^��&X͒6������l��������k��>�w˩�ۊ���&CeG�U*b�x8*1�Ԙy���A���6��`;�P[K������t��GR�Xm�Z�A6�M�3�Ξ�������%�y�G����-Z�T�w,��m��b�ii�!m��omjh~��a����m����aC #��B4��2�c`x,���P42:49����#m�:������^�s���}ׇ�������G�v��^႙2yjc�\��:6���p00|kޱ�nز��e;~L�������X}f��<IF�u䐸�Rc�����w���4�J8�"�ˌ�S�	4����o���x,�k�i�_D���ܤ�bI׳-�m9l)6�K
J�����1m?�cȺ��Td��2��$C�ɱGȇ�ԒR�9mUa 6ux�%٦U�\b)Up�6M4m
�{��6�"m� �JOH6�����g�a�ր���7׃���{��W���J�XCS�Y�D�Ib�����"|M�[�J�]{Y��?VrMOH>�p# R�0�T.4r�8�^��Ǭ�Fr K##�Z0��.i
:�&�.�t�to{Ų���a�_��{ <[�n������|�+�|�;����ш�hj�%��ǋ�;wn)_8x� �8k֬|N�V�^�0�N98�r�����<��7o��/ũS����q��X�w  ��v�'d�ȑ#�����SO=�3?ifAK8p��yd���N�e�g���͘1��zp�̙MM�Ui׮����K�2�s���)��a��� þ�ۀ�>����_{�5�]�IgϞ�s�N{��Ÿή���\+W��C��S��jnh���	|��p�T��^��5~W�y����ۨ�3�|���+�M�@���U[k�1?��a�+�
 ��n��y�+�o������)<~�^6����&Y��.�����;_z饊&C��:9(tw�'-&�e�l��zLN��C��R��VΨ�4�&M�':��^ Tw;sL�j);�q��}F�7���[���-���\�!�op���(ņ��JB4C�P� Q����W]u�'��.\��%΀�XL\�1�?��ݒ1��V��"d�c�a(�jM�� } -D��&GǘL�8<��>l:~*5�u2�\?�x�� ]�KKB�Y2c����B��X5$sfM��%�*MM����/��p;���[�3թH.T_��� R��Hcp>���΍I���(��j�2I�ݱ��}�{���t�]w]�~�)�kih��ڋ��5�c�	&M�SVX3M�F!i�Jm~\�#��I6��ߥs�:簹��-�Kku�O\�I]$��IL�`� �m R��5+V��ܰ:&�0��~���R_*�-g���\-���~<&�W�.t��c�<BWU���;�y�(U���J�Ys\zw�j{�ޝaM܄/ګ���-j����q���Dpk����j�Se��ǚRU�J�v9j�te�]��Ì1��O;ϫ@07�E�_��&�C�1}��Wv��6#ʈ�}`/�}?JF�\���B6rE&%�1����p̘�-�|��c{1\��w�����~J,i��/��+�^�я������^����˿���?��O|⁯}mtxdμyw��D)�b�X�7
kn=�JHB(p��)��A�r��6) �#4w;�zd4��I������K/nB �9��564��'?�fsK�.�.���;6n�������C�x���-����ys[k,ɧ�z����@xՏ;�͇�ɹh��s����=?FxAu��fp9�(t����n���[o����@i�7]I����2s��%&:�npx��SZ&@�L�>~���|��n�:v+ʤ��#B�4�c�mJ8�Y�FpU(��]݇�$��Pr��ɓ�(�B�`Z��$
l�NB
�JCPd��4��!�BWzw�+Y >�C�h֐��#�ݿu׾������b�zn&=6c�4&�-���v1TI'��B�ĆtJ�H2ayqaQ�E�%"����mU<Ќ��p���4bȬ6vS�e��J;��5e:��&r�8u\;VէR<P>W̦�n�J�
J�K�`��.��q���,�U+�����;���DhSF�Ң��	��D~ߥ=��*�tc���>$�V����P�ϴ^��w���@r�0�d{����Up�x I������PX���-BY��p�6 e�1J���K�lz1����1{L�L.�B�:�~�Ա�~٘�D����zE��m�K��5��`�HJ&��d��dz�zՉN�T�f����?���K��رc�<��}鋀J�V�ڼ���f� ��􈘎��z$��'Q`�dX��L��ϵj�&&�oU�N��%��+���.�$`���s���Τ1����moxu������i�~��9��82��ԙ��alذa����G��8�b	k���猈`�9\S���!ur( !���W�T����*J^��y�C��LNP%Y��ڒO�w>���lUs2+`��`�5RѼש�����i]��1̋O��b�n�hc���^֗yazY��̼L��(f/2��u�%��шW;88ĻP�Xţ��u�	!.��8���_[��u�0M��rQ,-�����e��3��5O����OM�����K�׋k��#	���Ùt������#�<�����}����ہH 	�5��!�HNF'9	���q���9�ݍ+Ce�'�����H��&�f6����P�o��l��'OΜ9x��i{f�����^�%s���%�w�^�{��CG�vW]wM�Ekϟ�S|�k�x������ͣ��Z�t[�?����aآ%՗��ݱc.8g���P��T*K�,�Ev��ihwQV��/��59yX0?�v��8���Æ�eD[Y�Ir�iJB��ܒM���<#�EO��j!?�^ \�Q�m������>��8^�Ðn /�^�R1	���W,_���|��\��?�e��Fo\9Dđ����ji'V9�YC��HO�k�F/6R���-�КS�q:-���X �za>ǯ��t�zF�S�8Ɍ(f@JT8�!Āv}��T()|j��������G?z�5��u(k�2�%��F��/�Fm�y�8ٳhUɘh�
c�Ve�sh!Rؔ�6����\)k�>;^PcH"�:ϼG�z�zVD
�)����L�bv`�>!�U��2���U�M�⸔W�5gՍo��۰�5DϷ\o�]햭.VE���s�, ��JǢ�N�U�8@]����X
�bϞ=�<������~������_���m24�ѣG��q_�ܚA�����B�~N��&��Ǳ�:;;.�����\�9s��<�W؝I{*�r��v�w��Z1d�����<Y��[N���r���_��'�o{9N�Ne��--"꤄?�J��XE�;�<2�� �l�2K�cڵ���s��/�]�~E�z�2�(W�[4jjA�����5�X��7.a���˺���H�D�X����	�
��f����	���!�x�X^.�gWyw��X�C����������/15
R0���aTI��/ڥ2sH�P���T)�
�XU��ƣ[��A�8���qb�F������~�\�C�p�ӟ�����?y�Q��x�駿���@3/��2��`�\�ވ��&F��-��S�/��cp�k�ƍ�l����ͦ�WE/���L��>���@Z,M���8z���S������::�64�dPx��x$���|����2a:�vǎ>�{�fjlx,9��Η�c�|������D��-�ٔ2�ysa	���6�r�9ue
�yh
��%����>���v�v�m��ݿ��v.[ضmi��E����G���ب���c	��ڭm�p�� �����_|)�X*��a�c:��\K*��)��}��,��l9L��֪rW>�_�Q���ʴͪ���������ds[��%��[/��h�ҿ�������o�@gRc��loR!��˭BF,<Ə蚥�C|S[�TJeK�=�C�#�GL�β��? H�+d���2��9������#���	��H%G	kñT:�N�!D"�KN���|;�S)�;��2-s�ʥ̙Ӄ3�M���n��F\�\OO}Cb4940p~�9�ZhT�����o�7V���|���i��
Y��V��/((!��F�ǚJ���G�>sCc&���	�1XN�$�\e�� Ch�������p��e�IΦ%�:�{FH�\.*�-�/q� >3t�рǥr���T�c˨��U��zZ�'K����˕.�`	��֪끹5hI��2���ɑa%�hhjj0-GY?���P�.ۆ���峹93f�X����cǏ?{������}rӦM�/��&mX�I�9y�J�.àƤ�@�2��}��o4���1O�n�j	z�6��:��x׮]X<]��lg�ۚ>�3��m�Օ��_y��7�t��5W��<��Llj�x<QMCf�j����O4yr;��_�2����\^�3�4�m�l�Z��xZ<�_:S��Ԏ����%c�P�t&�Boh�Zp����s����ЋH�U�Z�F޽�7x�����\b�������&C-�உlN�όZ��*��i>��輄 ���(ž4�3�`�*�:t��fhh�[U���'t��TV�}B�y",s4��@�jo�}��]6���X�x�y|��7<��y݇��� '_�-��r����푃�!�fL?x�������O|�w���O@x$n���a��P�
�M�t�`���xww�]�׋SZ��}�������ǀJW�X��O�8�p&#�� ��WM,�mcݺu���4�M���8�݇8F�2��~��ْ�J�a�{�����⎣��=p���a<8nD �ؿ��S��D�W�5~	Ɵ����;�y�5k��y^~q������ta0 4^���+�cb��{�?a����E�L�d_���z��:Ӆo	I>�x�R̰,	��mPϨxX�8�����s�(����@'P��=��7B���Hzv3e��:S��mZ�\r�;ֹ`�'?�Ɂ�$����`c>&e:�fb(~R�<�O/lm�TRW��Cخ�P���b3V�6��<vC�GQ���Xt�oFy�[98��|�K������g5��Za'�C*���2���q��z׻?�%��"ɜ�]�-.�x��rkҜ(�Q��jΙ���;�Ф�KElR{�h�b��C���5��F,�)�$/��ւxQ{��=nV�\��ː��<aP��ht�T�\��a>ŀ/�]�}鍭0����q�8��ʹaO3��yZ��i����Œ�rJ���x̼py�A���D��H��'k�s��A%��{`߾�K?���a�Cq/��Ϙ1c֬Y\��={��[,X
qY���?���K/ng[d�����W��1Q/e�y�<䋢����*(�kn�Ql~)��l�B!/Y��`�9�<����.%���x9o[|�ZK�]~�/gI��`W۠�
y�N�Ҭ������U;�R�SJ����>1kP+ S}fy)w�Di�?�/p�5�j�s�j��e�w-.�3�RN���9
�i�P�+'	a�X��e&&�`�R�7��>�t+H��� .�Ñ�4�|q�I��ň��7�Ҧ۠�/�Y}��.XPej��`8��Q�&w*�G�H9�p��u49Ն�'���",yŲ�`�|A��?��~���R����[�=���E���@ߠ��K1���ʌ��d�֜5}�	tŰc!���;~�0�v
,��Zw�ډ'�x��Y���D�����9s����7�|�0�e�ő���ׯ?r������E����.��Ƥ�����)���`�C�_x��SO����铰�ι���3]�^x�h8VVk[#�0���Lg�<v뭷._���׌yؽ{7Fx��Q����ɻ_ٓʤ7w���b��^�f���8OA��#���a	��u��RF��ПW��2�˧�c����d�(D5�f�����9z��X��L�b[�z����=}�Ѡ���=TX"�Zf�ؕqq0�
�_�aNl�x��;Y��kÊ*d��t{K���H>����\�̩k֮��_�����Tztp����rr�?`�S&��B�ˈi#�?TS{��`+��/��6�<�ښ�*����A*e�Tʮ�Ĳ'���HY�Ś��*��C�F5	x[#$�!Ѩٱ�آ��Ѫ���f�i�)��E0���Mk���{o��f�.�9}F�r]\��֖&H� ��dt9�X(h�τid���ϵ5\�ψ��g�*å��E�:F]� �d���bU0W�5�L8a�̐F3`cH��>iQ�W8(}(MG����m���6��������Ę�m�̘?`E�h���ލ�Vt�:�tY���X���H&���@ ���l�=JP�!*u�a���Ln���&Jd��(�* 6��S&wH~��\"Q̋�)������l�p�V֏����m�<	|֬�ݸ ��c�����ü<zp�x=L��.j��v��u�VL/����B����^��B&]�e��F�I�\ٸq3pۆ������r�_Q�s=ڍ0�+�s�:)�

���(��\g�!~�!�j
6�3G��R�u(���yv"q�*����)�Di���$���h&_"/ڸ�!nXK�I-�h}�i+E@�ٿ(�nxOD|V�G��5���|��˙4�S�Te�y�~q�+\P�Y�g�f�MpT�\��!�{l�����
����h3T�y6�0':$IjOS��_�VA�~������J �>��x 8��ӱaK�v���t5;�2K�U"��H��xo���n��s�ĩ�s%�Q��g?���~ݺu��3g���v�:�x�b�=9ڼ��y�1i�$���iӦ��K�Dw�޽X�W\q,u` �-`\[[,���z�?���-[0�/��2� ��}��������9r�̙e˖��uT�5Jt/�<�)!�3g�|���ӟb��q��'xSci�A���[��ųoH_�g������
�Y4����0n
����__�hf�������1���&����"�)VX�޵��(���uR¦X����bI���B-�ȱ�3�)�#�:uBDL������*_�_#���;�lŘ	=��:�kا~�G5j�п[�FG5C��Y,;::_��B���w�:�t��������o<�)�'"�n��.v)��f,�&�G�<�=��Z��4�j��Y�L��y�w�A�M�Q�I������k��2�����ՒLb=��������+�/��x�a�rX/-M����BL
b%cw$%:;���e�_�b{�Ä�]��֥Ve����dZV�����}����Wf 8�����KUP�Q���g"l
�����]�ꋺ��^�>��amX�Դu�BQ�#p����IT�{|�װ֋�99�ayՠ�&����x�)�aéV�I�8}����Wgj�4��%`�0<��OV�L���~p7�a>�+4��P��	PSLщGC��-�
N�*�ћ�[qY�}|��S�\�i2�ae�u�]7�p��V3�p��>v���3]R��y��}�cӧOw�wħ�g6�d�$Sk�Q����Q��[{ޒ��bY��L�I��Y�In�&���u��]����,<��|�`m��-}�?k?�`H^ﾪ�p�1��+�l�b��q9�ø�y��ˉ���w^�ͮ���O������N��=�����E��|	)�˹b<n3Ӆ�*,/SI{z`�-`DcaUg~�dk ?$�d"2��z��(�]�`�MJ,�����$���#Z�"�60�p�Ys���WR�-�,�*0�b()�n��������slG����E����Ų`>�?��?����o�=��t-di�����G>��]y��:����gh`C]�n���+w�؁.X�yL��ι�gL���+V._�hL� v�Jhǎ��!B��ۓ�o�����K�-_�w��=?�c����?�ַ�u������ ��KK����Ck֬��1	��� �]y����Æ��y��ҵ7���c8��Rm�q�J��lhl�0h�'��\�|9��G�=������m��,\<�>u�4�������>Ȧ�,u�K����T*�	��7��(���"-���|Q��
)�I/�R��0ޅ0Qi���~d�|]����X���h�8֒B���f2�`�\��t���ɿ��^`3�\�k���=n1s�5�,z&JgO���8iR�
cwvH�N��׸~��h,��/�KUl$�IK���5+O�:�ˤ��"A��U~�3AC5	W�P�VU����gh
vY 2�OG�o�!�����/�"p����L*�7�  `��]�8��j`Ē^�d	��Y2�V����9���K)L���"�G�����Ώ��o��=]��D}|r{3TIcC|x�h``,5j�$D�e����j�0k����ʋ>��E~�;�B7MYkP�~�#-���&�|>qU
9l���_.�|~3�ϐ��6GRE�,�>��<�;��F"�TZ�B�a����i@9�U�jZ����eҭx��Y�1ӻcU;H����X* 1��[�����L�,K���g{gG�diڕRI�(��WKOLؗ�XJ��>��ԉe�����Bv(9�Ϧ�0g͜)�k,U.�������bڞ�Xʦ%��S˦���V:5����ӧ{{��9���?k��c��d�1��G+�o/���"55�~��K�����[n����[�|ya4-��������ŗ�Ѽ��KXl�Pa���}�"����Lքu!k�>_KX��K��&�j':Y#l!�*�B��a�Q������AC9/��Y�Y�QѤ՞����`Ũ�������Q�	����`����èƲ�.j����č�^R��Je��1�Lw�������U����n뉋�R&���6Բ4�UN�E���RnA�|۰�a���,�{I�NH�v&����:���5_Ԙ8pM��$7Co���s��]y�h%�#�8|�`��-�-x���[:k|���j���]5��ԞLaAg�w���^ BڵkעE��J�_��_��?���6�#~�lv�#G� Xy�/O�8��>}��1�f�M7���������C/ ���F�=�i^X��f��ϣG��I�4�br�m3���Ů��
����߻w/f	�f�O*w���#����WE�K��(,e�9���W_�y����˗�p�������㚳gφ=�JcuS���z'@&q���f��g*D*V���+;pH'J�l�1=g��� |�E6ys�{������j)��,r>o��3��_���0��b1~�ىdI�\G2~J#��Ɨv����f���T_7d�b�4#;TX^��gY�Z���T��l�X�=3�-]RW_n����g�=�-��s��N�9��Y��HHB�Da[��`����{���`���ϣ�S���~��Ʃ�?��BȒ���RU�Jo�{��{O>g�����^g�P������:g�}�^{�9���K�Mu��N�@:U1ˁ|��ܵk��ɓ����p2�~i�BS�ett��C�������������;44�u�ֳ��`�o�41}�Ⲕ�֭���0L�,������h�.����ngB�$�����L��B�q[��CL����*a��:� ��ŋp~�w�;$)�	>8!X��=�tE�]Xԩi%�WXq}J$�6"l'q���4+�N�D��Z�˂f��עP�I������<qɈ#d5��Ip���1�Ŧ�j�������#?yn�f�hU�O��q87���(�Q?t�&F(�,���C4+�̸��w�yǻ�����=�V*9��J�/��򕯼p�<)*?[������������G�+�5�ڎ�Ho�>�h6vye�T.3��ъ(�����M�n%���>Yjp�~�f鿖�k}��bN%�2�M��v��+�o1 *��^�Z��F>�v}�ya�h�j�9kAqf�Aʊ�^~�8fN���k�̡��":�F Z)�:M�/ҙ@��(Ԩ9𴖵,�i����\\*=��;�'���6*�L��v$�������gv*#
�d�x��v����;��s�F��2���~;��?���mpp�o������/}�ر�7�t��@��}�Ξ����>}z8ovv��N��e3�����^�z�Y�ȇ���ݻ�r���tY�ݱcoww'����$��M7����D]�R���+���z@fJw�e���>/����@�H�紴�-WV ���b�*KK�GuW0��ab�<Bzv4�oY���� ��e������#�<�<~�=��9s���1��ѣG%W:'5/�y1_�M\�T���ȁ����:�K�X��J�u�8 (q��u::
��ޞ�����$�I)�،$��&����XZ�Da�ـɀ�J�
&�N����tc6/GK�6�Oz�T&��8�9=R��Eh�KK�z��T!��լ��Fo D_����3?����6o���Ҝߪ1��ڪK@��W����f;��d>n�P۶g�ߔ�+n=�L4Ze!�ȸNf\���:܄��p�@ձ&���ObgAG2�Z�$Na���*_�;epp`��yiޑ�����>��~�=�Ve����� ����ű�ѡ�ᕅ���9*TWkcC�W[Q2k-�LІ��~�S� ^�|<;���
�z�UZ^�����?~�4�?�����\� �v4�������q�kl�-��~è��ox`�~�V�jj���XS�%K�1���7`�cx���&����n�|�[:P���\n����Ryű�`��S�#��K=��`?�ۙ3��������*M�$߶*�Ʃ���������0���,[e���}�1�Vq��ѷ���l��/��uY"�O���4&��85)Q�F�ȱS�+�����>���O���}��?|��?��?}�Ob1�ܱ[�˵(u�S�������ܾ�����Z;oО�l!��3�=��#Q%�<�ԉ�����J;	�]#+�68��<y��4Fc<҈�5�<
�� ��+q�_q�}���H��(�+sC ����1����ΤŃuÐp���U�K�N:*22��d���Hޡ޸7������*�_KBʢ�\<R>b�0��d���0���LLL���H�V��l8�cJ8Ms�,��li�y�D�������۶}�_���_�������)�O=��ɓ''�F<��!��w쐎i�D0�=v;W4�uXX��܄	��z���_<�ַ�unn���.)����Pllt��%ƃy���BA���r���؟�ŗz�!���͛�/^����
�������$�gjwM�M��<���9�t������}�ӟ�����?��?���fȘ�����x:�6m�;A3N���j.E�/	�[\���s�����ï0!�;�.Z���@r��|�~8`_�Y�aN[�,M�F4wK��UI�AGڍ�����6dr����p�D�0XH���1�>� ��]eL"����Q��"�UVw�6犊�R�
3����˂�ccf<)��jc�Ӷ�r������y�i4B�+�.��~�[��^3y�^������dU����7�|�����'~�?~��[o�:q�DР��մ��4y�L[=����'�+���g녒e�}��Y}�B�רl�;A�:�Fd�WR�K*���E�J�Ťzْb>�M���1ElϞ=�k��CC0A��A�5��,u=����	!*j���t�P�xSxY=��Lx��/X��\z��:�����O������X��ř8�����d;}��k��P�ך�(�Z$��<iے���C�o%�|��H�'T��(SuBF���=ִ��}<�B���Zݽo/�öm����?K�Q��,�<�����7����A�nh�i� �}��w�u�/�ҧ����V>�_��?G3�/֬�W�_�`[�BN��%����VIS��鳆�@(�!�.z5�ޚ,:��X��g'�Ww�)4�F�����7ؘ��g��+��@=��(�7��1�5	...��I|ЗBf������
�թ��H!)�-a�è٪b_s�����c�=����H-q�G�vLX���l���3�;��x�@�@U=�L�Ѣ��IXܴg�,]�ȖpRU{Y���ꗬ��K{�Bg�5{���Ė-���o�<u�駟f¥�M[6���E7�?�m��;���n�?z�p�G����y��w��Wo�<NK�k���q/�߿~Hk��������V�����"m�O��3I;u�\>{�ȡ�'^�ɘ%���Ύ�9i����t	��dȴ�ZM��-�Ir&\E�D��э�@��I�I߳�>��O\�ַ����ށ� ��5�҄�*��b�C�'m���G6K�z��Y]'��BNXNBݎof�,��JE۫�R1>�J���OB�mu����;Y:~L^<��J��� a��lG��̤�
����cajj
Ϣ��M^�z��l�")!,����ʯ~�vZ_��7:;���K�~�j�Q���K}��������f�%�~�³�z�����Rs�2����:	� o��U�א��N��*+��Y���t6*B��=�si%e}F/B��w�}���~�R����G�|z���R��'���|6�^�x��o�ܯ�����]�Zefz�����32������I �0�\��7LO6�\9Kq!����@�<�������p~k�?7:�.a*���E�V�gK6�p���!،]n�)x��D��fᔔ�INc�^k0,(�[Ax~RJ�:��r��q١�7��9q��2�K v�s���eAG��Q�4a�!u Q������+o�����!S)׬T���+�)��!���$��w�m�l��J�V=xp���[���0�s�Z5�|�������8].W�NL�#zc3O���4#�Mx�c�#����ژ֎���X��Ps_��� ��,�`zna~Y��n��N�;v�9p�@N٦0�r��<��O�9s�����0����CK��`����;~�~kb�V,z(�a��6$aQ*�n�K	_O㊗�*�5��i{�#4�J+�`���~E�uJ�M�ZcBu��^�YD��b���ZIn��NNB��T��4=��Q���J.Μ�4Y���n�N6 9J���0��V��/*6��?��s�����%���c��8��R��nJ�ԞRU�c�v�U���jq���$�D��9�Ǐ�Jݼc���b+��+ĳ��P�uK�^�T�e�5r���4ت|�o0d��Ϳ������}���n٪���ʖ-[�5᱄����|gq^���0z�:u�Ν�۶rg�a�Ȥ����)J 8`���Y�!�R��e�+L�׾�5����(�	T�Y�Yf)i��H%���c��o�*�M?p`�����a%'cl�U�����ٳ�n�q?k0��I!���~�ϑV/��Y8M�-OV�:5��!����q�(L�،�%6V���e^\��5�B��T6Z��Q���kظL���o�g�k��y�7��G�m�_��[x��f[}�5kqY��v���|$����G?�������9,iV�.�/q����w;��z�h�̡�ԣ�jԦ�pm�^&h[�6����H�}s�c�a%�[�z�����z��>l%���]Kw}���D��y������?���_�G_<~D&ͯK�|V�(z�w��9lU�[�̀d�K���
Re({���*|g�z	(�:N�bUƐ�L2?��
	P�7)�IR��N�OQ�̎��E*�8���;���a>E�]�j�H=��U��`��]XZ�6Og�#P�k�&����8�rC�k��|�ո��b^��"/=���J��=�.�u\C��ï�t�M?�S?uT��r�<88��\�ʺ��0-IA��qb�bS��ͮ�m|f�^���f%�00���ۥqI�B��{��۶Y����=����_����ϝ;gk'�M��� bA�������Ļ�=�y3~�4̈7Q
6%?+p0���@釩���4b�<�R�颠�H�n�i��EkjQ�:V�(|?e�Iω(�<s��O-�@"�u����W|si3)�'��3;�W����V
�٫c�k�i%똀B���Sw4��R��ى�aV��d��/��4�sHFI�A���~�ԉ$Bm�-�T���u2^�Eڲ�<��Y�Ƕ���֪n��ؼ��� #1t�F9� �\u�1GM)|��'�f��$Z0��#��.V���;������>�y���ܥ�g'w�ލ����x��|�H��KK�sB_��3O���w��:t�uG?E;3?7::
�ETw�ĉR���Y�u�1�4�a��]w`Ϟ=@Um)C�
��~�k��V`��o_CSܞJd�Ê�U�/�ߒ�����Q��;�� %NL���h�޽G�a��lV&͖Ɨ��N���9}�蔼u�\�{\���!�X�������r�X���e
|֤�b�V��d 첪}�G�'U��w�R���0C!&����Cҝ8sb�g�l.�x�%��4_jeE�S-����{��e�pEw����9u�<��=�|Vb�.�zqq�X,8n�3&yZ�)�:��1<8Crk�J��-�=�Xу��������L�Xyo6癕�F� �2�
J*�l+ܩ�ʅ��jqi�3���g?�ٮo��I�Qǜ拹�ׅ	�]�U��I�)��XꞶڊa}d���/g��x�G�uԾ�c�Ƕ�_i|�%�z�g^��,�Tk��c��z�F��� ��f�`�T& 2�	l���G �2�_&-H�e�X��nl��A�� ���j4j�R8��0�J�+��2KW�i�&�I�a�0l'��J�Q6��啒��(v��~f�����Ϸ���������|�j���|6רCڽ�}��);ZM_R�]iɄ	K�t�
�W�M��U�f�z01%�����*B�63� ]���n�㮏�w���7�j����L�oE��T�'�(X�}���a455��'�Ʋg�>p=����7�2��s3V1�C�s��~�u+ʼ~=!dʅ��lr#�lNۿEOJc�Xq�8�)���(��Փb<e�i�n�1"�R֕�|>�oy-���@9��~Kڗ�G��|־��?��ܚ�ؤf(tY�P�9���u�F�N�NGK1{�� G�#���c$u:l��S�e�����	Ӥp����!p���-�:%{�ֻ�Myp�&축W�&����A� ���n����X����W)���Q�.�tkcN����^�@�a��ǎ����o�ر���������O��6M@R�b=z��K�� ����@ES��c�)�(v��3�H �J���!6�C����J+�W,�yXI}M�s	h��++%|qdd��w�0$�ƃۇ>~��d/i�*=UP�8'�
K:]]=�Ӳ	>Ly��l��mԹ6����|V��9X ��A ��Eɑ�H��ŕ�4�"�_��0�����0xi���D	�ہ����7[X7�&����>|��u�����̩Sg��o�9s�2_�C3 }��k�S���,����5�fv�@���$ ՜�S�h/�������
�J��h1�,�b& eD����s��o��_�՛o�1��_<w�`�[�'b���e:���5.�R�`��m���H��N<.o�&���W_K���6;j��,i�=L�?;���x)/#��o]�ȼ1��`-�h	G#���O�k-��_VvC�C<<���i�[�G��'�����$Y*�h��7!@��h��YL�?�|M�&A;Zb'�jE���ݝ]�B�����}W�n�����j�{��?<<8$�"�e�`;���$�"����~�U���4r��7�\������}�c?�s?�䋖�K��#�������P����
oE��z��١������{��?(\s��F6��� 'm�|<f��	��X_a�ny#�U����\CY����&��a�J�{[����Ȣ B��Va�:�r���I��+*�N�i.i���o��.y#|��M�lY�6�͊�D"ġY���Ҏ�f�����jG�7�U�+KJF��=0�����?�c�=ztvn
�KTc6D�����-?�:n�
�D+D̝��ryI{WM���R�-��X���v��F���7v3lEvF޼x�<��tW�s�W��m�ɻ��בq
ǎ���9b����f�.*�2̜��D~�U�::��BM 0���5�����[ka�{�� ���'��������y��C=t��o�Z���5������,���)�/,�"���&p�]�v	���w���.\��PFC#����no�>4ǒ�]JZ.����D���ŀ�U:X�x�Z9^�ҨK�2�3���ą.�M_�mi��}65;0�<Y~�`�Wk5�Pm�W��������F��l�C�#�[��|(φ��w����!�	vK#�g�z;��e!��\��SJ�͚�{�%��%+!:b&���4����*t%������&n�θ��!����mO�q%R�jM�_κ������^ܓ�[7m-�s3�0(�+�����!������`�ߪu%	��δ�9mս
Kk��uW�.	����4�KA�H�$��9aϒKE�$$�ۨ�L]ڋ�����q�A(�:�^|�-[�\����.@����G<�������r#��nFX+�J��S/,��LL������X���+xyLw�����A�)\��fݩ8Rf�A4�������(�ʹNS�w���[˃��^�\����LG!�Y��fԪ�UY�9kl���SgNO��]����8:<��_��?��wK�xm����H�D��b[^^*�Qy�Bq�}J�b���l�B�g���h�7��e�i:JȔ$��i�| �R�.�&���͉劚ð\a��Xq��<�|ƳX�^�./�@Q۶l=u�i�W�U��jUʆ2N����䍾~bߎ�b���ժ�lF�a+2�3�f��^ !	3e�r��[>��T)�G���G?��7�PZ��+��������?z�ι�A� 7�5����:�=���։��熁��u����$l���=}}�c�6)���+�n0��)ea��@�_{��8���طG�� 9��������o�i�R�i	��8OEπ;W�Jѓ&~Z��q�Z꘠��[Z��%3�YZ��x������G?��v.ת73�fy�Q-�;7������ ��$_�T:��z;O�<9�}��w��>=11Q��R�%�Y'c��Z�Z����:`�	A���Rk)�KO�^���$�-JU�J:`�94:Rm�+������*�����C[ϟ������y=�\=�qdt:�؏�=�"W�O��F�I9 T��=��j2��W&OZ> �j�]^��e�1E��cJX*�˂;�l�A�t�1P�L�@��q�*�P��(a!�k�[/�������o����A��7$��I��:þ���	���I<Mo��L��2�e%Z�R+�nmv�Ԋu(0��?.�{�J��葖0��li"�ﻴw��47;�� [�G����0E=k��?	=9�Xc�
�Xw��LH!�����fŉ����>���?���>����A~--/H��V�d����W5b��v;a܍f+YلۗǧeP%e�f�"���'���OK�A>��i�-G�dZ*Ec�؉)��Z��i���S��(a�����`xUtf%��h۶m�<�L:ص%@�x��ngO7{�l��&��`R��&�rU��3G��$��hM؂�E���{�vH#��B�s���&KG�<�T�ѿ�������~4� �}�bz��"[�;�b7��'>�	��w�x�ĉѱ�7�xci�
��Ϲ�D�K�J�$k�c!kLm�>�[c2��2��$���7_} �*��+� �����`�֥�jx��83�����c���ϲ*]º:�	"'��Ft�$�-Z��<V=�7��ҁ1Q��UA�P�������R>U,J�]!�����q��H>'&�I���z]u9'�C�nQB���" �?O�o�L�C�D\�t�M�}�v�����1��4�=22"�Z����(`���:�N�n�:������#�e�r��6m�t��Y{�����z��1�����&�L']GRST3�Q����
8|��P��g?�Y�3�P�bo��o���������ǐ�[���;::
��s������?�70�N�2�����U�Y+���bYC͋;��DXm>die�������8�0O--b[푷1Ѻ������f����v�s^����Wk�����暿��a#�����xZ^$�;i_��	�����F�6�։�UID!����>z��J�uf��}�r��e�T�$OYX-u�A�cE2[���%뷛�\���I�]l�}�m�tT�)�ܩM��H�i�Ʃt*�����^KXB�Hq��cMk<a\B4\{� �ձ�����k�ه[�z�/),���c㚈<g�V�j5e�V��<�����B gWʐ8�T)K��0�����l�&\'hEH�<*�fq	�L�~\�<� ���k��$��U��h���$~a���-q�j��8�����jH�b6�vڪ��\�0:1��a�����l0>#��m'���ωy��r�5N,5�F�?*&/��e�A%\�����F<AR�2�;��Vo��HI�;n��1���@i�d7�`
U��z�S�����)���9sjlt��������~���O�?sꤛ��N���f&`$��9VTo�\�	j1��ƃ��mq�*�3�Ä��J*l�\�N�_^�k:��|(�Z'5��>.��X��0hYQ Cpdx0�������e\�ܬe<���k��������*%,]�)|�W��m��՚x9�u�u-��K�X{�������yRmԛ���r�LH�[C�[�n�4;���dVy1�e_�v.ep�
Bf�@&tJ�WG�!�&e�[�{�fR�|��{���w�N��"g&�!����)���F^��UvI����;����ɯ��u�U*��.`�T[�,�O��5"��|v%�<ࡏ����-/.t�ڎ�-d��2��07tv(!�Ъw�x�B�O�ö��d���i�:I��X|��8t�}q����C��'���[������/~���y���e<����[޼y�>�A�i����{������d2�o��ᘂ�Xv\f#�٤�m����@��R����_,t��M�@+`f�aV��GI��L�}e�����c�e%��� a�LmSv����೗�P�0�*^Y襯����0)��Ga�����e~X֮� !-C�X���ĩ���X.�&��m�}ԩv�?K�Xf��T3n1��,M����*��9�O��*Z�#0²I�,�Qr/IMCW�3v0�=������Z7I�qз�*'8T�,	>H�T�ZB�`���\�[�e쐹���_��_?r��-���B��c��/� XI^m5Gi~COt!fL��[��-�F������D�e"�:��	S���sg���?�1���N�\q�k��-&sõ�'Fp~�K�)	v+�_�������	���![�xbU2�HrA{�Hպ
qYL��| ^�NQc+�i*'d�/�<�()�k0�I�
�lN��$pG�/�%M��������i��#��7�BR��~�J�S�����}�;̪�S/�0��[���!���#��wߡC��KFFF g�*���%!�&�琜�Xh�Q�yf�^ ��Jb��=��o�C`����⌽��Ah_���;6�
��m��v��w�fg%>Ш	���X�rl4%/��SF��%U���(9�I�W����^��KH1JH��x��q�e����!
�yfF�����/^��d����ĄH���q޳�ϰ�	6W�.K�?i�iau�`�l��I}�V�o`��1MLL�n,% �&&6�>Md�T6�$G���o22@U��;žܩNC���J#��9'�0{#�� O6m��7?��a�?)~q`��eiA�GF�D&�>�e	�H�kG�w���ːQJ�͛7�ڵ�K0P�h{�C>�����ӧO///B����ѡ�}��������i�f��ٹkt���L�����_����GI���)E���ii�dE�J��D(�{��ҘIAdn�o���	�:kn����OP�9�-��]�?��x�Wg��Vc$[C�6�s��櫍�7ϙ��Q�#	���S�B�g�K�x[㬢�*H�>��2��"�fK�n?3V�j��7z{��:�z��\^\)t���Y����-.��[d����	�B����F��G�~G�n�������k.��f�u&+�Q���L�#L��*Ȝ|>��̯,.v$�����ش_��?�����&�`�l�;����$D-?����\k��	��^��D�^͆� 
�+"��W�Լr/�R`��BաB=gz{�fg� p�%�}�r#){�X�<W��)�w�|�Қ��|.[��<�j�^��aR�9�L3�&>+]&vXa�*D!���d�\в�S��}�YI���Zl��e��IL���9��|�&T�����G�F���v���%�����K�2��������u����������kE��z�T}F�j�U�r��B2��A�&���E�M��j�f���z�|���tn��ݻ�u�m۶�����-d��bfds�=X-�ؾ�\֗�	[�;�t23-�Q�⿸��4-�O��R;5����C����ߐþ��.ʴ�œ��ք}���X޵mK�V�׫���s3�����^�opt!��ǏWJ%h�����4�j6E܈N�R�~�`->��ߩ|HI�M�:�uR�
���赹�lG��	!H0)nBXx�ٜ70�7=7lD�z�y��9K
�s��/B���<��ӝ�"�B�a�d���R����ˏmi�ˌN�<��$,` �ɗf�T��ذs���BI�������s�'����͸C�4A%�-�A�Ҕ���eq�RiYv����~��터1��� hL�O��x�7��1[6
'�F���[��^�p�ܹIWɆ��J��x�	R(�[Zo!�"K�%Ҏ������+��`4r��3/���������زe��[�n�Tl�<N&�3D(>���7�4�������0Rr���c]�n��7����P�h��^�ԩYԥ*|(��E�K^*ljU�+�il�$����X6�Τ�,@m�h
�e��Y���o��j��Ϛ}����ς(+c|�~oz|�jg�a�a҂��&��ԧ0fRа��H���a�a�iE��[-�Ȍ�0���N��I���BML��e����K�.�����.᷸�[IC�(ix�ů��ǵ֒;��4 U�Д)}��ᶴk0���+n8������GG��.:�&�6�-hN�ϯ�Sc����7���=����9�rV8��0 �(l0�
SO���0U�q"��ͦ�D���'L"�V&��2�Ĉ���x���Y�L j+w_$�ޭ E�Z���O�ڑ�\V��l|)�ɷ����!̵niT��Q��.��# �k��	+�ԭ���J2��ٮ�I�(2�8q͔�if���E�9+�I��~���xm'^Lf�r������o����]���%Hڸ$D#	��Q���-:�n�p۶m�sK���G##������{�'�x�Բ]|J�#�M�T�z`˵0魙�y�ǘ��Eb�tSLy|-�>(�j��q˖-���Y�9:2�5�k׮���m�&�KK�+��Y����.SX����Vؾ�e���v¤����Z�_��Z Z��5G���]x֦-[�يi�u�������[�ne�ɱ�E�� y�������M��i�o�SV��m�93}idd�)�L��G0}�`����z��Fa�|b�/�!��.HB�J<mc��oI�MvvYN��������n~����c�𣀧�3F@�=R�q�b�is�f��䴰�Ox���{�č�8q�u�С3g����/����޷�v~3���*�Ȯ}�J������5#�ה;��#���2a��r��%1٫XQ��8F������F�Ku- �J%��!��8�=
�����1penI���lN`���"?3g�!���
5Wnϡ��c�R�=��D_���A��+����1�4�V��܃����~ h��P��\K����aX�nn��_?�d�JUb0�
��@o���(�|6��щo��i��Q�S+KS^Mth����bц-P��r
�ńr$�D�C�٫ s��(��`�E�=\;����Ӎ-�51.E@9i��wuI�L2�
���g���d���ӿr��|�5��e�t�� /� �Hn*ږ֍g<�
��f�;n`K�2�2. A����{���TG��2��M�C��zmv~.��惂������jz��DYK ��ƽ�]���O�,Yn�./��Ix�sE�m��s�nh�T��#n���:��%J
<��� S� �������u	�+|)�'%�I�֧;�	��AW�mj�ğdi\����G���#?ػw��}��^�X���� �|�+@ר�������#-�T�+�|MbS,��4V.�>�F�R����ۛ�U�ƀ� -'�>�y˶����������{���𝝒��x���|�^�fi�U�&Y�f����r����*�H��)�ѭ�'�s<��̭�
��?s���z�ػ]��ҥϊ����`���76����^{�=��Ξ�}Ѹ�vm5ߨH� �]XX` �Rt��b��/�e������ɣ��g{z������P�ks���#)�~�� H�L^���$��k����#/4�E`G��p��v�6OD����H�������e�	�O3�Fnv�E�$.��e�9"Z�F�R��ca����|nԫ�_iyIR-�2W���-�x���ԋ�F��l�|�$"��~ҏ�;�q��������xqz�����~��?���<�1쐙����ጕ1mv�$zЙ�<�r��Z.-C�*����y5}��7o� z�������vl;~������f;�����&�CR��U��G��;�z,m��Q��ͅŕ���BQ�I�2�"L`�+4�¹"{�K�e.��um[q�Cܟ�2x
�\�w��d6��|�2hb��FA'�'2��P�0g�In��1��N:��gip��5 q� 6�*���J�aQ�hi�X��?��Z-qV5�ԦBZ�ɐ� K=� $�_TR��$i�L�!`R��{�m09]��
�-&D��Ȓ������k��Z3�O�����H͕�+*��\��5�2�f�ˁ�,��h��P'�D6sKW����2@lLE!����v��$�ܹ�-7������O���ojj��񊹎�*�;���Iq��tK�aOX����.�>zz���$�W�@��0��q��R7����	�I_>�b��քz����13���1#"�#mDc�*`]���E�/EICC������obT@���\��N򱶷�/˘�M}�\�݄j��Q�b�єg�]����������}����/���g5+� v�EE��/�������HZ�s��3�0YMF�2'���'�>�3�����W_�?~��3S����/?���C�+9:==RU��,T�G��n���ِQ­Hel����|���\��

�a��R��u�־����ӧuEI� �?�>W�%�זn�Vb��aZx�?g���ȼc޻�23����k�p.'�%-�$�f&.��l��;[*��B$��⺴T§BX����u��<��J:������&I�rEc��箭�#]��մ�s��ŋx�5��;44+��ڶR��F>����&��<Gd(��x"��K[B�]m��g��ٟ��?��?��������⇠�}%�<{��H-�@�;�J]O[$՞={�z�'�����o}�[��ۇM��3�S�q��dGQ�sxQ�c�����VM��3v��ؘ4��ȥ3U�Q��T��`��i�z姟^N��t�f���ד�e�u>�B"��ɓ'1՘�3g&g�u�����E�ߴ6�CVR��
㴳_�}go8?��> ]���d���n4��	?Y�-�����a2K|!����8u|�sǩ��%��Za=nG<�T�*[�cw�ժ�4�E��Œ�X��Z�Y�w
�=]g�M.�����}����8�r����cY�%_+	-�2YN�H��l��6:z��$�����J��d��:e8g||<��e���%܍Zc�hN�\j4�##þ��+vtҋM644�m�|��q�t�Z�������Z��}�S���w����w�뙹��rupd���y��S�{+ah������\._#\x�<۵�~��Efe��к^6v�Vju���8����/�݊�������f��Vmd3RJ�2�&fa�:��BGM	('�w��npp8�u�ҳ�e	�kjZ%�BV��(!ˠ��C˦�R7C�-/����T���r�mL���ˍ�N=z����C��ʋӴ��v�IK�����j�-$@�R�ܹ���2�4u� ��J?�m۶I�Ǔ������JFmw���ߺmi0��Z�2�l��fKQ.�7����/�~�N刴�)zF ���p����9I2��g�-&:�]YY��關°�(����G1]ݽ}���_����<���|�S�N-.,`��ٽ�%]���ْ�2�gP��Z����Ȏz���U.YXZ��'��J���[-�7���r�H�(�����%��o�'"��2h���
�ܦq�
�ea��,f<-���F]� �ު%��n�#��1�!1*�ef�Ç�wR�0e��k���H���w�k��޸�<�B������)%'L����{�RY�~�y�i��oi<u�"V������H Qڹք�6�xb./|�~�3Ҕ�e�y#�T�ZP�ă^��'ON~�C�馛��/�B�3X���ذR�i:��ϝŖ����[M�Y=#��+�9�N#
��ak��M��fffN�:`$��Kb�t��Ѥސ|��.r,����@�d�x��!��������}�K_�[^��[�N]�z����|g_7f&��k�!t�}Cҕ.��U��ťٕ��Ħ���%\9��u=��98<�a��(��S2������gv_{]�\�vv@3g�9>6���Ș~1����>!/Kn �J�}:5�N��d�%�Z`ډs]�j����/s�Y��[+r��K�3RO�΅r��s�NIa��/^��6�$7{��oi�fR�h%$�u �ݖ��:�(�I��o�j�$XGL��#ɋ�B����(��	m����oͼ��"S�`�[&�I2�8�#o��嗕PIYIA��T���E;��N:�MDIS���$�dqeF�%�ǐ�x|F��3�!��Uw:���$0Jl���k�M�6�����BY�K�ZjӹU�.1�����x�\"��@�޽��Ҷ�R�'��#E-��t��'*w��^J˕�>�/p��ki�ɳ0����FGG�Cԝ�}��{/��e�֯}�k_��W�f��q���m�f�CyK�����i�z�:��ˬ�g�&�$�+�74�ƴ'�I��:5��Ɠ��ZO��9���+�PTpI$�(�R�t�O�����a��Ɯ9�X� �l�4	�3�t�I�'-��4���(ޡk���ꕖ,Z�K��]���s����ܹs���h��&��m.�H��%�p�v|sW!�� ���{g��/�%z��K����o��'��<�O��O���v\��ڵK��fI�;%m@
��u<'鲅�Ђ,�֒q�6��ξq�`%l,fk�o�{�����J^���oy9ZL�+Tix(gٝ�W��(u��a��b��s���86t\�C�a��#��Ջեݻwc��ӝ�w?��3�^{-ο4?��\�\�\��ư+!sHf��A���n&:�7;���~���o~��]y+dj��F�K/������:�e�aؖu4�����0����)�F����!�P�f3Y�A9	��ז���̔ѷ�v���������A�c�l;�<�J���<�d�������>�C=�{:�*���x�n�z���6�@�+c�>�}�|�;�����[��ԥ��N/x�픍uD�j7��ۗ]*�P�99�V^�a����dŔb%`fd1X�ӌ��ɜr:�� ��3k#@���Հ�90�~���/@��o�A�I����=i�&�$Q�k�L��+9��u����hV�c�xca�|�#�$٩�#(jY	D��(���͜�ҥ�^
X�񺑱��I�&?FY�,��	���<v&��{�Q���GI`&I3����4�g�,���b�V�7�,Wz��&uHK8�d~��伮�+b��ڰt��E�*a#��39y�o`��0j��z��K��޽{w��366�\Z9y�$�a�<^�b��X��)�!#_�V+nO^�K/i3b�X�_����B�4��,�3a1�|�hZ��'��,Q�����"�[״(-K�\���V������q�	l'�6��+�6������Ԫ������Ȟ�N����V:�ĸBܹ�sX%�f��IrE�Akc���'�3@�(�B'�Z �J�fȼL��
`w�>$��S3�2���Z;��C�*��d?Zwr��r�ص:�d��S��Ǡ��l�{{:
����#eٹ=���Ư���o����y���[ �xxx���hVm't�H�5��K��L'�m,E��
ͤ7nN�B<�[i����4�-k�w-��b!��F]�{Z�j�7�F]�6��5�U��&sd�؍���х���2J�q'��Y9Q8H-ѵ����"?�Ŷ1n��,r��{S�f�ã�D/͸�s��W:th��iaW�� �����|�P�g�7@h����0�f�0��`��kl�0�>D_yE�1<��Q���iṧ��$!Dl��w������-N�ٹ��۷�kZ����p�Q�����S�->� ���V��x��'>��|F�tO����4����b)/O�QW#8�F;j�+�j�;4�{�ĉ�o����԰i8�ܽz-_��ދ�O�>{fC���hf�ҙ��7o���ؤV�K��..]B�E���dm��V�V�|��F9��5���C_��]��G
*l��.���CٚǓ�+�Q���X\\�+N��Z��4I]�gqj<��%�8)��8�L�ph`+פI��O[z;��k0���\���Y����  ��IDAT���R�mSv����|'f�x������C&���%Mcb�����e�fv�sFq.�M�+h�vXm'v���6m�t~*�����H�9p����F'i��/�굁�f�ZZP�J���T�f"�LL�A����oL8o��R�)Fl1m���
��}V�� �ԩ6�Ο�����cǎ���~��ߟ����b4͖V��6AZ "K���i=��#5��`n��o����f,k��CsM��Л�G�'e�
X�d�#�d�K�������aB� a*nj75.6勊[t��fVE��N
|�C#h�5��1flLLL$�9� �1:o���,�r����U��؝��,N\��v�l(�^����s�1�q��تN$���1��<�V=��7�cǎ����w�u׋/{��Gx���z�R*C���Н���L��.���:�h����^�#�H��Q��N �����-Ӗ��T��ʒ�u���U�k;b�aQ�6B�\<=�5H�J��U�t���ة��y����ݜ��[���4�IGd�N$���a�@�?��3[�l�䜛�W�V<�==}����!f�/��Ș�-����ĖLb=4�8�����$�a���!��R��
��Y�.O�{�@1B��U%�ĕ��96��1*B���d�@�8;�|�������ܺ}{������NE���H����|�~h�LVD����;���x�ޫ�[]z\{��yِl�rI2�ff�q�P��w�g?�k"�Y�9�~��Y���"k�ZZ�4&���Rj5k5[��`$\A�E��|li.&A�QW��wʁxI0�|:؏��m:�V3}i�d�5�Z������M1��*�F�!��Ȝ> �7����O�M҆��A���D��9�����N���뤢ZVR�$�:?u^�Xmjj�/$��R!9��	�[����l�:�LeC$���j+���K�>�ȭ��
Ë�ǑcϫK�%��o�i-��\�KU����''`f�&1�w�/t�He@u�P?� �M،QK&~Z������;k/�簸��9,,��ސ�ť�B��{�"[��q��m�����}���Ǐ�j�����\Ysl��|��6P�f�*[�`�F2]���۵�Ջ�+5R;�#,հ��&P��f҃Al4��Y�Ң�LP��Oj�ڎ&n�~�W�����O �۔#���j��%)n0FY��-Ɔ`|:�'m���M�5�����ǒg��)Eo��Z~��/��(\s��C�h'�8�T�B��)�ub!�k�0X����st1�(
[z��i�������:ё�!;JdS|/�4bqVc��tiO��~�v���@��	<׋��o�:�}۽���C��ۿ=���O�8s�u�K�g;�����R�a;<��s�ߜ����Q�wU88�۲bm'k�������
�.��yK@l*��5 �:PL�:,����D|)Z�zv��Wv��:�Cmʐ�&�c������nd��씞�D�Dt�#ܸ��(r6��(�5[���2�ن�}��_��r�Ħx�Ԅ�o3;77 �2�}����O�<	Г�z�� �P����EE�122���@C�{�pW��c��>44IH���ބ�4�>|x�֭aKjB�2ZZ5�u���b�V��f��<{v�Ν�}}�Ο�MB('��
�����/d��*yQ�я~t�ΝՕ��V�I"5a�S,��ff�ߗ�VJ#�ö��fS���dY���<:����1��r3�_Ú�N0�a+�es��ٹrI�����|��#�>�ַ��w��Q�@P�.�`W�����E��k��F"��\��B"��`�T����~�/gIlx���.��R� ��ŭ�s�.L���s��ә�H]�9xw1��:(�)h�6��V�4�����!�c�ݤxѣ��>�u��n��������6��|���V�t�:�J�Zӳ@{����L�0�bR5Ҹ1���zt���w�O�7մ�xYi�Sk`�9r놷�$U65�?��֩]�eOO	���N����55ڍ8x���b�$EV���=%,1�<��=�fϞ=Ĕ vR
���T3m����I;�k	�$��ReA��][VB��Q�����6'V�z�=w�}7 ��T�0��h+�>]�¼��cL����r�F��=?��R��^�b՘�����`w#�4O�J=��0��f͙@v�p[1�vӬ��x�Zw�6jtj(^��A>�$0]x�ܖ�%,��RI��ĝ��X���@7`Juc�A�B�I$4R��椗_� }�xa	ϥ��u*��.�?�^M6��9�r�e����D��>Q}��8{�,�1L#�+������w���� %�K��K����ؓOB��2[le����Ջ-�� =g7mڌo���������U);$����TG�'�s�E�_����'<�q7��e���u)V!�v(��R� � m٧Fr�k����..�o��Y����I��Z����O�#&c���!čW_u �/��H��a�9uqZqUM�j����Sj+*]�v��
~��,?Ě��L�45�!��K��$Jޙ�#RA҃�_�����4��d�,�f�E�Y��q�:�$I�e��y�P�GQ���V��i�y����<xw�0}B�Y�ٶm۴��~4��4_�"�)\���P�%���J�CC;v쀭�[��axx��'������w�qG��x\��(]�䱪��\9jsX���uW��ؚ��_��h%�W8��I��$���HVq��̔�B%��R�};K����1[�+�85L0ǰ]�I3$��L$�z%bjéHz��yF�$�uL�FZ��*NRl/rB�v�U�sƉ��+���a>�Z�q�ͯ�-欠٪J�G���%�)��#��؅q
R�b9`6�R��j*C�WP;��*��𹌇=ii�:�A�y�>s%��R��a���f��)�.kxmt��zYU��f�\�bgB����ٚNkI�-&r����r����~�رz]B��=�h�\Q�x3�-��ۧϟ�p���͛e�C���ҖD�J?)V"�5l��$.L�,���uC��H�iW�gY�\H�p�[~+h5}��v�B�(�Z}��e0�*��Jy���ɸ�b�3w��Ɗ�%���ei=o8�:q����uv{�ڟG˃b���/CT,�B�^�������Ev�՞$��k,!sث�M?փ��� �ۤ�S�:�A�\6V�2��5�=�����l�E��t����;媼����Y���B�)�ϥe�a|�M74����C]�a5j\'h6f�/�;39���ܳsWO�-_�6��"s݈�d��j+ڭ�)���סf58R#��'l�|ױ<Wn!�8�^}��,���~Mv{ I\���?����a }J�x�^5�}���r's�Ĺ�zP��il___�Y[^Y,��㣣���P���z��S1_XYZn��@������6m���@�d�H�h�a#c9Q1�Tc�_��6��<�/��v�ܶ��b��MNk-+�ީBT6�#�]�]�Uط�<���A�� ���P�Y�S�j�wK�I����`8n޼�����ttX:Z�^&1�p���������92�]�>`�zcx`0�J�T�e3��y�6����K��]���uw�Be,�+��v��h:Q�fw����|��|��R/+����g��у|����	�,1iXܚ:�%zR��O��&��͎teF�u̇,L����OcɯY�k�D��H+�5��J��Z�t�ף�,� � �@�liٖ�����6�0m<seÕcK�)1����H4���j�^�>O���g�&2��c,5�U��g�;��`jg=�߫?����l�8E�!{{�z�M�����D%:����{#l?�ұ�1,gK3�@��i�e�`{x؋$����6z#/\���\u�5��T�D	G|&ISv{�P�~#m�6��7��Ồ������7�]J��JyI(֊E�A���:,!�_�A�ʠ�w�@��d3x�eɺx�x?q�ͷ>|�+>��n�>�'������ɸԷ���z誫�r���m���}ܾ}��o�Kxz�ӧ��I ^�Quj�X�ģدKl��:L�v&n����$�0�	��'IV����]ry�ص�b�S��J�_U�{ݏ롈�ת7��UVG����G�Βe�%�j� ��� @'��hY��e�^�UT/,���	>/���Z�mɉ�Wx�j���F�Zf�FW�Qe�DR�.А�H�J�rb�T��s�"� Eo�2e?����9췆e�!����P�NOO�d���Ǳ� �wdy��`��|F-��H�dIT��!���F���@��֞{���GZV2;�(�G	İij�
�C�αR�|���e�����^�52=���ڣ���X�+��5��	5&w����`,��g�c�Cj!O���G��IV��Ď։��7؎�Q�~l�Ì4+��U=pvƄ�����m�|'������Y���|!k�7-����~�#?�_��q��Q���R|��ø������A���w�څg90`���xBQ�Q��;��V�r�L>#7��G��}�lie;!~E8�}�]�z���a�v��sd?��ꫯ��4�sE�J�V��˭B��]�����>��u�]j]���/�7�F�,�H�<�w���F�ya�1�V�.�t%�e6��m+�����Y-�JαR�����J����,$<nK�*-�_YcU���Ƶ�~�L�H/`3��'0��R���k6Dar��YR1%;��6��Խ�� �{_3?��6�g��m�j+��[����$�I�-�6���z;�9�w_�����5MBX�\����{�L�\�D�dC�[��[l�����K���N�m-���ly�TtY/.�:oۼ�v��Sg{|������326z�ĉ@G��<�7�� I˸��k U�p�B�)Y���8Q�B�n��]><���������ll̩/���s�w��F���t )�3���`ǃ���ê���8:2)���e��l�����Ł�^�Z�4�R���*�,��t�M�ӧ��������r3��s"A���C��}���y�Xo����RFCý�=�#}�WKne��e��:��`�9&�eab�V���t�M���כ_��W+���k�uq�I�H��ʞK���ÍcnM�`iE�_H^*]7�˕%�c$�z�W5��y��s��Q�T<5q�ZQ]J����C�6�fw��V�Y,G�Ym�;�-!��L���ѣ/���]8/�]���S'��]'���/-�h1���V�����٨wtu��Z��-�:l��R�x�$�f�V	4%+�^%��� ��f�_;)5��[:%��_�6|��1�\�.�9�m�D�
Pc9�J��zƥ7�b�윓�4uzT���%���8vز|�V�[~�s��v �{x:��S'���*2"�{϶}W�l4��S/aE-��esq�J�������j�0�+��8�c�wɣљ�rj6jZ��鳚F�Y֍r�K��$�૤�Fq�i��=v��Ep&�EJ'oK�+P��� ��F`�k,�Ewű��묵z�	֚hc�b�"1g�Q{�Z�V�vdm�(s��ͥR?����\qx:{�G����&�=*�ÃC�� �����t� ̩��=�����;q��S�%fb9�� �wo�	�ċx������]�
�?�[&luwH��cg���V�J�C�v:a���sss�؞����ei���"�5�,���(�~=�������546c���G�i�=8��0��5PZYl��4�z�\̹��+������wܱm׎���E*�����
�͎lJ��g���������WZ^����w��plx���?���]W� iY�"�l�{����5jV$��m�"�s�N�˅�~�\�D�F��}7l޴#��z-<��sc#�͖�߹�>�OZ���TeA�X�~�TFQ����B�P���_j������]�"$\��/W�2��/�,S0�9l��	\U�  fwQ�O���4�U@B����m1�(���epii~ay	x|���ɓ'�f����d�J�M�;�U p[ ��9[m������J���|"U���m�9�����a�{�|1ҬTA۽�)���2�ʸ�f�4�y=Jsҙo'EZAl'����Bv����"Q�e�z:j*�q<Մ�	�6^���Q3ƺ�TDF����R�r�Kx4F�wB�S9�&����N8�F` �S���{n���o��V�11�	N�����;7yVq�����[v���$K9��&&,ۛ_�o�[�0%�����P1l�����������ށ���a��_��R`x�O��>}���D���IF d�2/M����cS�w��?|�)\���Ɂ��V]2�<���쑅��+��xY�l	ZS;Y��7�ub�e䘚+������P`���4������WVjZ��%΃Xv+�1��&g�9ƅ�&�DD�;]Ҷ���8󂸢���,�[p̧�ug���VC��Y�N��"��L�RH���\����ڣ�Ћ�h��V�NE��::۲,Y�K3��bk#hCo����Q[x��l�(�Q��W/󕗺��`dG)pO���	^����#Z��bJ,�U:2<F�'� �+7�>Ǭny%e$Ӱ�m�뎁�̐���$����U�YѨ�b�D/�Cַ��+��8,��E�d�&�3�Zz>������L3��̛����s��af�rC��4�,�8�.�t�����O>���?��;u�$�4+��UW_�g��C���Zcjj��w��,�ͫoU��0
e�U��0ׅ�?� ��S<GTI�o@2�v4 ٞ={ �9��/b<��|P�`�J�v�l|r���y�{���o2�Z�=˒''M��������5{������.>=;���a+�~��a�r������޽{������[��|�9n�B���CC�b�wv)߯� ;���9�g�d�)z��5�\��O|��ýS�`��(-�]��|�Ͱ �T��?bk ¬L����Mf��$�{~���:I���F�]����J�/$�	k ��q�������]�z��2-��6�#uX���c�ڎ�b�Fa�J�ִo<S-:�כ~����O���j�i&��Q�4�ę_�K�f���N+	s��B�o�_r�j�j�V�Y>ԋ�-�L�ڶ\఼���,�V�7Zql8�u�)�<x;����Ї��?t蹛o�ւ�I�ؽ�zz�Z*�w;��wd�?�:M� ����&��VI��TN�<y��W�G! ��.O\�,�Z��H+Tv�Zf�[H��8�U��:@���^�n�		�AF\dlb����gϞ�B�����ܿ/~efj��c�����Lr@,�eEfWf
�ʄۏ�b����ZG��th�S%�Ox}���_��O�p�~�<L��Ø`�3���V���{�`K��L���߷�K/��Kݍ�@@:F�$z�B��������q(����X��a��a[��
Z�
;�������������������ׯ$ũ�x}oݪ�̬̓�9y�wr&�Չx�	z��l'��d�h4��d�h5}��м�$('�/�cg{^�������M�gF؊�$�ڎ)�������.]��7BO۽{�Ky��b�DwO�(��-ղO���������!_�� 
�0W�F��Ck;ADΧ�����UK�{�f���U�3LT�o�7�  KpaN������@��V�2��Ҙ���O��C*��dY>s�o��R��QG5�0�z���A m�f��VdIj%Eʨ�b'P�Z��T���@+���S�3�Q�E�}�GX�z�H�%�A���tu���& 3!Z#P�,R���X�sJD���}�6���)�-[�?����������7������T����K�;w�w��Mˎ�]ҁ�K���lsY\���������K�|�����mi�d���pZѩ3zd�^ww�����|Ш���/-��2́��U�u?T+ή]�$.A%�e�T*���q|��ꡐٹ9� �xk`"��� �8���l��M����
�V_�!S��#��R[�����ޔ��c]F�Y��������犐�h��˗!�-Y��b��y7�$��S���t`����]�h�~�|&4�-V�'�(x�S���[+���8��D���&�i�H��>?;���O.\�Ŀy�f���"���|	j�`���4��7�ka�����Ɓr�y6ƙZS ����#.I*~��W�4⼍`$vuգ�ָأRZK4i>���fׯ������I��O�}�4��$T�wq�jG̍�嵗C@�+�q��M��K�"�B��B_c��܃~�}�vR�s�����.�oY� �� E'+{��d���Y�~ ����?��ّ�idd�Y#1!1]1�Q>��"-�31��q�OpC"��$�9�� �n޼�ހ4�{��!![R�4/\�pG�.l۶W޾q��������z�-ꋌ9G8z4��J[$s��ɦ_��n�A��OO�n)J�?��?��?�o��HEHءY�"��(}QX�t��濦�G`���� =P�}���� �(*E�4��te�>�E�U��%8��O>��_CI�'��G��v�ʍ7���>A�ʛ�y��n��V�s.	ZN�<�8�a��`m;��h��i�C+�j��Z�o�O��wP��#�TE~�F��w˚�71�B�q���4h�tD5�U�%v��U	�!q���z®s#bB':����8�=��Ɖ`�mx��#u���jJ��W+�ፇ�^{p�/�:�~+�����`���Q�B�^�z�N�PS!ȗ�����n��O��D��w����p��yȴ�aɀ���|:�c�	y��H��?	7F͍�bm��g1X��⭂Q\�L�߹�Ye1�P��BpFCi�����㏙��
+E>'��j0�B ]QÌ
M�3<�;�s'����N,���V�.����i�GO>yO������6�Z�կ~�.��޲e�rSQ��:Й'���о�z^��R&tww�k=���G�sFXj]�@�g�%-}�JgJ��1�S�p��-�L��D�Z���Ɯe�k=x<#ٝY��LO� tI���*b����45|�lݺ��ٳ�h/^e�8��<;�!�*�1��S�P�	=��cC�l:K�+}�̭3��&���O�xƬ�m�Ĭ��(]{m�hl��V�6�4Y��&:�^�� 4��V?��K-�5d������S��T��H� w��in�H$�S}x ���ufvjp��ҥ�tzp����o�{rZv���V�X
�0�6�K��}T�N2$)�����.!P���'�ƅ8'-�^;v��X!��:>������w�t�+���`���_Z���D�y<OA�@K�D �pb��.���`�O?�����O�����O<�r"Yf)��r�ȼ�$�e)���h٪�dۊ���t
��lt5Es	�P�I���o}�/��/��|Vd� L$�*%@�B��b���v�5Vh���s�������=�J���x-*n�������8��(�7
;eh:~moY�b���^[XU� ��4g�mY��2��TU{�J��[Q2
������W�Y+����c�����>�eNԵ�Yi��k�I;�k�,�������0����Ia�i;�Ő��-eɯ��Q�P����0�;T�GI|eh�nl��ՙ�r�wAQ��$=Q��r=�`��ʗ"�ã��eԲ���5paP��k�3�?��}k�yԍs5�����Մ�b�������e�f��ׯ=����]n!�%R ,z���f�>9=30��x⇚�/B�9!g�R���!�L(�/���Tď�b�,%(0�����^6�4���,5� ���� P%�V[�~#In��z�E.�C���6������,�/e�[-�SD�W{�ߢ��#3?�I%Nߺ�����}���ڵ�c��x��S��,6ww�ܝji��G����P��8����l�����ٻ}��'�|�ڵk'O�W֗�-����Fw	r�B'�.o񳹼҄oE��~��_A!z��{�u��NHګ鴵_]qf/^��eyl�ڼi ����/u{��7%�\��>���H�}�s�&&A����s����?"�Qh��2��M��u��S���D�,�����_��=ՕX߃�Y	s��K2���X �t3�E�R�ӛJ"�r��-�k\�&ޤ~@�T�'�&$ ������?�cǎ��� ��ZE�'1�a�g$�wE�6��Kg[4?8.�dT�5(���b�p���CD�-r( g�<j����\���S�@ pJ�s�6��۷o�A��}w��	j���˗%Ɂf�O��/���o��oS}D	h@oH:�)�E��Lms��}�|�	i G��IVR�|^{�u[�g�xɤ���e�L��d(�2���^m��Bj�*�qwHϼ.z�0ASww�*�+I/сd�zun�<�]	����=F'�UB�wcbdf6D����|��Wj�	��De��ȼo��7r�u��ȣ�Ύ\���7�&�9�֒�X�N�J�zAh����e�p��Y�xrM)(�m�h���xW�b۰eY����+4
��p�ѯj��� ���N���ڽ+�&��V*��� 䓉��~#a�e�W�V3��ƱgE�4;�ڲf*��$oݺu��Q�yH׹�9̾W^y�z��������t�T�5c��+�$��bCK3s%���=fR���A�2�6�t�d*.�Pe��{��2�-�ݻ���z����k�� Õ���w ���6:I���'���{�!��[�/��5�U:f(��2�Z
�� �ny��ќW_}��wo��Hot��Lg󑯳%~V�;�����t(݀�XP(�>�J~��'N���~�o�ݿk/%��b�&�F����i�����n��F��lB�T� ]�>��������D�R�0I�,����h��$�N�N�2��ĊS�%��n&�ч>��	U����jlT�F1�[Iz��YTڃ��/H��Y+ůn��{�\�3?����.M��(���]��Us��c�X�\,ry!�P�>��|��$�(�(=�W��
eFɰ�9ٗ�g�0����L�)���YۖsK�c��lČ*��#����z�u�LNa]� w���Ӝm��활�_����$٬P���۶��B��6�q�nh�D��+g�V�,k�t�	OgJ���.9��� @��V/�S�	7�_Z��eM���gϞ:u
��FMLL@̍������o�A֥��s�΍��?��#.z,98�ܜݽ{�`��B�*dQm�Gp�ѓM�ƔmC9$�V�D�"۴���3)[��`T*��~�~�̙3xM�>�c+5F�*y�s���g�dBE˖�!���u����mW�#ɦ�(� M�]�r�'�x�X"^-Wp���U��ƖM���t~���v�ܑQ�,lb!Ҏ�U�<|���3�>537w�����Yq�b�󳳨�db�d��4�)Dk�U���P$y~܍U�*=�dvx�mZm|1�Pώ�fV�2�jX/�5&�Z�:�3ӭ�p����%(JA`��D*5��UT~�l������3��`P�$�j�$s���9�����`%J��G�B��ۆ٥��ي��u�|n��!4�q�5����]k�E�� �}��ZE�C�>�h��n���ք��h	V7jt���H�
D�v�������n�kW:�ĝ�ya�޼uӑcO.�KK��|N���u����v��_��]M�XTj��ǲ�a(�
~K�$�.* �S�����1a�]�� �䉡� t6Q�\�Z��={�a�]���*P�%m�\A�si�@�C4Њ'q��(�vP���eeia���mݼ	��4���Wo\�m�+_}ehێ[ã}�6�<kv1��Z��o���6��0�H�b݄���9���8c�Z��Gq.;�̑#GQ���o�9[�pU���C�\7�Ż�W�f�w�*��"0(H-9Qe�&"�W�Km�~fv4{������7����*�-�`�x����B�짟2�b�	k+vR�q|�E �n�Z�NA��}"Rv�e�^�ɈC*���b?O�	�Wk���:s����EDB�(�@����*�g�س��[Be+��;�ج:0��B�
4�0�ڹg~L�&��GNӈmV�!��'�@�(*�1���������;y�d���pFH��@hkI����V��9{��#W=��X6�С\���cB* /L楥|�s��\���ʉںu�8�)5C�%(�7�S���v��e���<�_z��w}��C����ӧO��(��=۶m�-t�qS*A!s�%O���}�-[��G���؅��U����Z�g����N{Uk�|�)�_��W���o�q�L��z�>����D�fU���mOM��J[1ZM7>����
��WV*�~��&����d6*א7n0�n�2�Z6�~��觯 �x������J�c�.�V�+4��7��؊�@}hn���uBf8,F2`H���9nP�Z�������&����fVʅ�Jֶ�=D���c
n$!fR�T����!��Gv�)��p��X4�C����nŏ�����+��ԭ7���-��h����U��C �_�c�.�������\�|��W�\������{2M����ۻeK�P.ٴy�K���������ĉT&�/�Hq7����}XeAǼ#-�q�v�u�vA[s3�p� �p��m�j�,R�|�g���+� �J��W_}2���޽dqT
)\@gb\��+U7o���ӷw�^!-��=Ƙ ���G��������o�d�Gw�܉k�S2���2���dP)J�%�er�<�|>Ų+�M�8��t��'�|��7>��#t9�:���xEv��:�Vܟ�Ў�%@����jG��n�g�D]uREO�k��L�-�8��C���x�_�m��R���-�33Xm�a��� ��Ʊ�J��L���MТ>Nu&��A"�ܩ�\-�+^,׆+��Q�T�t8����k��u�����L�Z;.
э1���H������h�$�R;ҭit���P��#�&���_Z��#L3��dM�@J�p�8��D����DK�UV%��Ŵ��<k'�
�._��%1A��;��_��J��.]��OPO���U6��i�ʤgg�Z�eJK.�d�v&%ۥ�G���ǰ�c��_�!B�kA(�+e����(,0�^�'���#��an�={V��r:�x&��wp���}���wn�V�'6�M�07m{��'6o�ʘ���D���R)� {��g�nh�ׯ_G5$�A�Za�-�	� y�1��v3��J�,�y�ݟ���l��L"������~����~Oo�ŋ�B��D�<gW\.x8���	(��n�-D1K�U4����˥RK[7(	���:7o�U�@��^µ�/2��aUE{A!.�QaA"r@Ԧ��ӟ~���[E�Z$�W���K�|�Z��$Kū��Ns+��(0�0�=�˜��4gi�zl^`}�Y� �_�ռB��l`�aik|�*K}�QH�';dS�3�cr}s�m���_i��F�Q�T��CyX
ӅW55"ob/�ƫ�6ώ�C��BI�X��vU�ޕ/˷��=sA���̧��Q�j�+Z�"�7�^�zFߥ��ګ�e����ʆ��^��Y�Α_cr��"y�n�n'�e�۽��c��;w�ĉ�}�k_kʤ%�i<6?5���˦���M��O~�칋c���1�����w��%?^��#O5���1s�	q������tp�zppprlS"��!q%P�!D�h�A �iFY����o�^�d	�����@���ux�&U?O�
�"�3 <J���۶cE�	|�>�&��
C��ff�˹�_|W�/,|�+_�����{[�m�d[��,�LV���vˎa�V���V�q��C��;��URA����d2�	�8�JMݺu��<�֎֧�~�VL��L�m�(���@�D�]�ژW�C�ϳ"�a��a� �~`T�e�؆�L�:_�"��F�.�8j�bi�v
�W���B����I�fB���ZF��3��*!��ļr�xܐA������]C�t*a������˶,3M��BI_�5�_����:5��Fp�k�e�U��j>�Δdڮ�)���`�$�T.��p�^6�FF�BFX��Cc;�R�Q�'�"�o��.���X`�1��a;�K�to�X�,)����X�{��刡Y��������Xl��](y����(�g�O��������ghh��j����O<!��M���:9���}�]H�/��ɦ��ɓ'�	�z@c�x_m��;ע�|���J�\�<���Y�>���ā�cǎޮމ�	�����O�6����
�_������T�;;�vu��_�.@ix��}%|��g��!���@���D���'�~�����2@�x��8���O��@��h�	&�c,ЎRNq`P��[�LKrz=��\�A�6AZ�X�~P"��y
K��$�B����B���V�@�υ��CT�U]��ݮ>�X��_M�RW4A�<��g�ޥ_��U˯+G���e�J7���C�V��"�ۿ��y������jx��sCq1o�B��e�� �@�Z`�c�A�▮.(���UD6fi��	|!�}h?A�*糸�mMNB\dSifP���},ےF�c�*&I�U�R �����"%!sP �7� E�?�5����}�����AxB�.�m5��&|���U�
�V�8p���R�`�v�"){�jKe>���V��^��T����U?t���XA����RL��[jW�)۱(H*��4�/}�K������Gh�\�j�]K� �ʵ�knA�n�p�Դ�uF;	pǓ�/5�2C`���iu��Ȳ$�R��K�r��]�#�|�A��(���%t������Ƿ"k�c�����J�)[�9/��;|���C4�s�Pڶ�j🙊���f�����M�d+��㭤(�*�Ex��� mјBb�Qd\)�^m�8�f�ێ��g�k�̺Jɍa)Mj�0f/����\n�<����'N�����_��_O%��X �����уO�V��OL�www:��� ���|�Z"A_*�D���xi�$%h���Ö=��ӧO�Ggg&��s�������Í78[�ĩ��b��aw�ҥ�{�b�����D*Y�I� ���C��1,�o����ށ����;H�8�m���ޙ���щq����H��P7�m�䂜�I�A(�W�\�ƽ�����b����(�B��险b����y��+�>&*�$�O�A^&���<���˝D�$�R>_4 ��x"�0�j�$���T(}�QT�򵣥g �̮
b-{Q�JybUm���2�	7�2X����.q��'�����{�*0�'X�p�8GV���-������.�����v�ק�}l��S�ju9��*��&�g䕩�=�����ٱȾ
8˶��Y�)���X��?E�1W6_r*@�Eڨ��Z+jKlj�v4��v�5�k�C�����c#�=����F��؈�d;�b�Z�Ο�p���RNf�?����{v�A�R�T�'qh�65�ٳk��]]��ϟomN�^irbč�R�x>�\�p,U����Jr�.,,�K�֖�@v�|�J�7��	-@q~Ϟ=��$	�l$�!�,���U��������կ|�G���?�����_�zmll���׶��o�Lϒ���GM�����G���,��ěZd1�xՄ%[���������͛7���w��1H���ٞ�����?E4&t�*�%����wV���ɩ��0c�m@aO�w7o�zoxt~n1�������~��-��v1+����S{YvP�0u��\��!�2B���#�
���j��b�i�P�(�Cp/J��R������'>�q]v/���FdbE���C��,d�s���"��ӡ����wU�"ɠT�jЦ�i��Q�� �|;"�U�������)����ڱ>���sx%��kń�+�O6)Is��@��2��K�U��e`<�|�������z���y����$�I\Ϝ9��Z�l���H[,,@����.�X	�-�M��[>�|o�da�B�"KY l�)���^4
�6���i9p#�"*܀JB#�p��mu�+C{;�؏~���#����� b����^ZZ�>|S8��#��z拥�� �\75LG4��-l��r* �W_}�CT��A͡������xM���oXP�p#�BK��֠��Ng���y�p:M���Q����?��θG�#|��$щ�{�|�f3R��M��v��k��y���(
������r�j'	�n�m*�Dn����Ը� ��°�b~ыP��Xج�����nf���k[/��懃_��^�ő"VJ�j�8Y����V)A! /�rf���^���y�v�z��b���	+���}õn�!��?����_�Fʩo�°�A�I̕���i�gfL�KB���B��ٻ�!D����g��-Ǐ?w������k�*)�����������Ho/D�mȺ���TB�����y��H⁹���,��שS� �~��w�ܺu�����Z�}�:> xA C��˗/CP�ܾk$t�@q@[F�F�$*\��8�K�W���WE6��E'@�>��3����Zt�Y����X��>��'9�B�@��!9!�Q%H{�����o������C�5�Z	�{�1��	7^+�أ�Nޮ�f��P�
�j�V%-�X����[C.{]����S�%!#��K	��NK���4���Fɴ�ύ�i�]�x9?���<�l'�f�o�h/���X���ii�Ǎ~�v-&�F5a��ᎆ�,�'�o!� 
8��`����S<_�k}%#=�a�$��*�1�K;:�����l^�%n�-.}���D,����1�wS��Id+�7c6Z��ؽ{
$����mʴ��J|�������w��-��\-M�L�rY�2��9
�1�1�������5��	��������M�F��ǯ��k�0�{�=	�>�tkk{:-��p��3Go���{l�޽f�y���ӟ���'N���6=z����w�p�Rv;t��;PyHOZ"�z�)� i��(ςL�gkV�Xj6�J@��2���O�j4�BG((�Ad��ю�<g���t5;s R�Z��i)�G���8AK�� c|������*�_�����we��2�bn�ּ>;���Xj���[�����=&��۾ma�%��'U�4[뫵RH�MOs���u"�qA�nk���s�D7���f�:�R���^�A��f3r<Z:�n���c _��C����l�cnP������j�r-���k�O�!M�=ώ
jDyk�8�ʹ��do�կz�qո��_��Ҫ��	$��L[*�W�~��v�z��!s$�jvƯ���ر'���[�C�+u����/�xf>��TD�Z\�U<�(fe��<o�d)dJ�j&���@%�ږ�sw���g�4��� d�-��zH<PC�~�ӟ���1��_��_B�A�<����PcD����M@A�,�$1�ŋq�o���[��H�mep
$c���0 k6��$�]� fTni�O8��D�iq""	��^����q]n�Z���ڽKH��W,Y޼y��=�F_�����|I�g(;�H��c�3�Z3�f;��vģaG�^�!�]a���E�Jݵ$5
4��u�]+��ܩ�?���OZ�d��!��~��A�f+Λ2�NO?r�hD�a�ǖN� R�[�XU��R+*p��Q�)Tbu5n��N�jLAN����=��$���e�ј�g�鋦�f�lf̏F�� b��5��ϸ�]-��:�/������2���pCe�۱g?���M��o�+Z[��k���� �@�CQ3�pݩ��Hi6:>�����MD�K<�Ƚ1fe&.����~xx�̙3����"�K��p�|^螕���{q=
���.�(��������ҡb j33�W�^����@�hH�c����7�I�ne/������Y��ѣ8iQ)�,`�tSӬ���9��#R���qq7�;p2Q�\_����GI�8�Y�l�kk�+Ɍ9+,�X[z �Sq�����)h�^�R�8���(��,�s\
��5ٽ��F8Ij=+b�s�X�0j��
�2��^E�ʾXݔY���ku!{���F�ֱ�������"T}�yֺ�7��V���ö�$�ְY6�]������E�NtE���-��8>�^����*�~�4����C�@�A>b��WnR47h��'O�nK(뗭�{&�ޅ�������~��g(B�lݶC�c�MW�ѹ���F_(܂�6��}�]i��������b+�ZH��������K�.�.�={�P��L﫸�=h���n�K�23;Yd_����tg��
mG3�R]xt��&��R"E��-�ك�D����I5�x��Z&�I�y萸J���E����q��Ǩ��S��?��-R�m��z1��L�b�/k�
wi;�K�IbK]C�`7�G�Z��]�AY��1��>}���s�(����^+�b��JkF�G�g��w�M{�߂	I�0k�CM��3�O����g��,X��;E�
Ѽ��� Q{��	0�mA��J��]-+2ڱ#4.��i���9='~Z��X�]�����P�eQ'�4� f83ھ��ǎ����پ}�8�����)���$��'`� _�Ub�K� ��ʠɦ3�4L��!#��dX%&';��L*�I͚����z�526��N� {�q��ar�&��b���܆�.�`%�s��J��O�X܎�&��[�>���B!���������!��l�J�)!*;jH�
��1Z5�e��/��ҏ�cL�64��7ߜ��&F��[�V��,�r�J�/�f��RU(�J�nog~u�1Z9����|���վ-M�R='�����U-q���zK�ߛ[��_��n!­�ѥll�f�̋)N����{V5d堟��&�ۤ��r�l x����W20�7�aB����?��zC�5F{C�װHh?SJ�鱤��,�sD���(Tɀ��X+��y�Ί�n��G���\�d��R����j L��:h`)�f��n4�!墸��8	롎0�Cݽ�b���X��C��DY����� <Σ\>f;�7,..��.����
�N��'?���;~����#��k�$2��eW�M��X©�7�&ƒɄ�m��CfzwG���,ɔ{z^x�۷o3�'�9�T��<8��s�A����+W$���׈���@2 c����)n5ܹsgk_�;�:!  ʾ��b��]ΧR(�Em޳O���6|��ؔ�&�)OB�9�� ��&��8|��B�g���a1\ZZ� �������!���߅�SRqSՉ�Bb!�21�YԴ����S�"�2`�^�y�9,ג�u"��E�Z�\nfzଐ������:[5?C�h��L�
��<Y�jY8�̅�"�T���q���+,[�	��{�&�2���@�HW/�ƳB���Ruh����,z�|���d��G�3�
���f�!���a6�T���*�$j&�H3����z��|䔯:B��JH�Ǯv�ڱe�L$�@�B���ø��WLD}���"���o�S�/�$�D�7���ؽ�cJ���oܢ>~�d���P�w�y�Vz�u��C"�3f�JǙg�̱�1|~�����I�٪zP騡��R>�����W(C4�5�2+�PC���Kē@T(�ޝQ��7o��axT M�n&�J���(j��zK%r�U��'N ����j�w���O?��dlx.q*9f�J=�X\E�A��������w���b|U)/�@Ɠ˅e�Dyߩ�CH)���5��%�iܥ�QWUCڱiٕ�'~��"P��h�˗�d�� �+q!��3�f�5b�P�дY��T�uf������Su_��7>h=��Y��/�kT�FQu��-�N~���(�BQ�n��VC��N�5�~��/Nm����k�Ўй�T�lR%6�RJm�s
"b�������k�K�D�?��믿��W^��������C�g/^޺u3�E�E�d����)\��3�^nS0���mDXU��j��W���O>����X�Dݱcǵ+Wu�_4rU�|��%����ɂ)��"�<�@� �QΩS��t�-��ͩxUH0@:肪��T�,a���S�j��rh��s�T�."�ɣC�ں��R�;�@3h�m�w`pa��|��
���Z����̊$=�X+3����QSu��z���uV�u��	3x&�o��A���FgB�c,��	,��B���
�~����!N�_4��?�Ry��R�ʋ��U����U�"�{�ݢ>���4zb��G�x�V�,c1���г'r��#������b6�ZD���0P��v�+�w|7�߲:�˧Њ�n��N3�ӎ"^h��Uvo�a��9���_�+�rk[����,//��%�JVKE�\*�v����ւҖr�W�_��zC������b.��e���10��ijj��O�r��5{������<��Gҟ/.�b��[o�{��qT��{��ھu��hI&��l6�LMLtuݼ|���-�ŅlS���-D0��&F{{Q�?9	=o�����jin�r�dWO{K[�o���\�׿���SS�g�|����bK:[���l�x�-C��;�R����LoO�ȽQI�i ��ٹ��#c���uo||�
*s��B>������	9�LHo�T���9���͆/�	�������-�Z@����\���$Z^*�ڵk���>�M5ۉ�1�x󃾾ބ��&����O��;r//���h5p����n�"��8+9�S��=�R�\>����˰��r�⨈'[$eܶ�~�lj&�R�MV+(�>���-7�+��Ԏ��|I%`z(ߊ9P�[���b�Ji�g��i���L:�I//�aV=�Q�\Zҙ�nN�>�WL�5�J�Ѱ�%V聴�*n@㶠F�ӑ$k\��8�)��z�ʬP�՞�0�_�����U���16���j9j[�����{Tv͖ƳԒ���Ŭ�e�[��a��
I�$��H�S�*Uo�c�Dsh.�=��^�����!÷���~Z-g@m�n����*?)�#d2��da����c�)Q���/	�Ŗ�ގ�N�b��m�~�䉹�	���ףG�!��.�t�wO�M��to|�ر+�o�^2��̛
oug�� ��\�� �L],�Zu�ݺ���-�*�\������R~˦Mj=)C[�-�����$y*�����oo�}ꩧ�{�Y�J?��"�;�Z/�dOopn~1K6e�*^ HWr�hdɏYe��W��x�ZqcqtV�����.>����[�&�v���8�$�V*�x�󽸘�=[%��e��&5�$d���ń�U���ӫ@�,�擮�k�>t��B4z9�ֻxi���7n]����8�nu���*�U{��P�qNڝߏ6�����H n;ڑ��ed7���}���p�]U͔"�"��K���(���R..�3�J�\(����2������U�ҕ��^$�<�sm�ɋ9��'��
����#eI7;(Nh7�$E�Z��Γ܌-l�)t��j,f�	+cքFrSl�7p+Q9L��UO8;�I/u��H�q��*�aG;�<e���Ͷ����A�V#PZ/��|۶m��uxxXx_���e�$no�i?3�&���{c�wu�GwrzS�$��1i��P[[�pO�1�CC��}D5������ڶlI�v�322���r��!&���z�� ���������'����x�"���
U��ж��a�Ie3V�S�+��M�W�\y������;��]�6??�jܻ7��T�
Y�9ʑ(9�D�
�B�x::�NQ5�*><Z n聬A��۴_Z�SAy�ġ�p�#&?���tF` A��ΦeQ���+�%s�+U�����Cw_/�V�@I���h���ԥ��΄���c����Ӵf�PSJ_��ljd�H<����4V^Db�a�����Xy9ͬ0��g�WRڪ&�K%�̗�b����T^��1�׊�kS�!��6z�f�_+Kݬ����&���F476^𠖿�[⡿���eSP�����9P�4z�)��EoZ�i*Y�%5��C ���k����?@����;G�=x��׮uvvBz���r���3=0v��|�J�]-���U	�]�JХ�9�TXؾ}���(m�n�t�@�9sf`p���Ο����pF4��yU-��4@/�����X�J>�mڴ����$&͗��s���hK�#z�œI�c����"%�e�fa3сx�|���XG}���c��dm��P�g2b�sb�NPg[��hW3�[F:຺�2�=�\����=�o�¼1�RQ#�*eZ��Guv6+j�|�C�S�(ɣZXC_^u��i�?!GyBs�04X��]�خFy��k]W�w���6�AQ07�s��X6�N	��.'�5ђ7���p9Đ��=0Kcp��R[�m�VT���e��2��2!(k0A�Z��R��.����ިńIvvv"�//:��9��ֶ�|�9R.KH `������$ ]��t�^�T޺u+&<fK�Xܳgϡ�$N����-�[�gryn�2���͛��M�7�Z���(P��J�yd{�W�'�����N�S52�T<������Lr)�K�.�[�f¨,55=ay)������Mnzv�)�ܴ��%S�u�\]\ʕ�E�tZZb����i���t ~B5P�0��N%Y�7o�}�6�K�ؗ_~�J������й�6=I<<⫭�;w�0�&����?�#����l�xaf*����ܛH���K%1oؒɌ|�VD�熉M���xN���㑧#�?]��G�l�P�夻y���}�q��P�op��������v^��~X�s�$��6$Z�W���} d�+��Qk7-g�8\���i��ϧuv�E5��*<�  �",�gf�+�"d����ah���w�_�*�T���Y���*���x�����ͳ>��өqR�B�-�ݘJ�wT�O�])Cu2g����٪��@��r��Ƚ����ut@��x񙧎�޽�L�/@+���(�����KW�����۷"T�]���o+G�Ŏ�N�n\����l�<(�_Y2+�
d��{I�Fמ���؄pۿ��'�bMI�3��6t|�\��:2�c�
��l4ױVZf6n�4�ž����������7�x�lG�?���m�p�W.������a�5����uȃG�ٹBh���mXQ����j�Z{6��h�zG��5p�����>>�Q"Ϧ3*�qc���&VG�v�6Q��Mn��ț�U�g5|F�!�f���J�@QM}�G	���v��>�Po#�l�+ǜ�5|F�
�����P�<��g��f�P&=ٹ3�-�
�k�ӷ�t�=�ଌ"qU�F�\�g��+^4��l�*?Y�mѺ0Q0r����R,���}�wGQ���311q�G�! )z:��?CCC���$��a�M��1� � �C�Qf>�CG7(:�4@u����&V�g��Ç/�����`����*2���%_�~�w��ȑ#�tdDC��������ף-�6B33��Wc��{2;+$@��L���B%m��RSK��$3����G}��߾p��&�>�^ 9�n�~��g��b�ߗ$KV=�W����CH��"E�&����7�
>S�fQ�wh .F��IZ[���I*OmQ1-KY�Ć���:�%֫�T85�"G���t��u�,}S\#��/s9_�����6^�ƻ���i)m�0n��~�u~���W�u�+|t6r��>z��E˩�bH�|�����x�X۽{��?~��œ'On�6����yHу~���޳���/|v�2T͠j�LLLQ������*~�Ų�:M�PB*���B�>����$'>@4ANb	�D�f턔+���|�̟���(j��AKw4�f7���V 9�<�֭C�ٮ�'V1���9�W�n|��1I^,I�&��{ 6��⨽a���
6��PJ��R�	 �d÷Tڲe�_)�#��O<���ױ��<��픢���V�+r��[ S����
�7O6V���J��?�?�(H�A����˽��O~��/�ϩ�4���vi�3[��L0�%��G��䯿F���Bac��[(�"�4�D4~���&�}�#欤����k���ׂ~Qm��`Th�R��]�,oʣ�Ľ-��Ff�����۵
h-M�ƪ��c';K o�U��I�ղW��tn)W)W2��x�������d<�*MMO�:u������^�Źbq|bJB��{~��[��=�L�;w�i���_<�����}ӛm���㘠B1,����'�*2�M�b�����͛g��s(�$=�-7��6'�����݃k � _��EI9�Ǵ�����?{��ݹ�y���$Hɉ�@0�������D�qm��gu��BT�&��ם/,����{
�d�YT�J�` �N�*�գ��?9�׺y�P"�D3�@t�̭a�A2�%r'fzr����dVV}Mٯ��x����%�lg�	�s�@��愪[�\��4�W�(i��K!�����M�S�Ă![��.��~E�3hXf���c=[�}�goH4e�>��|ݙ�+�9�֪$��A��h�/�A�����oեq�!��n�.m�{P�7:I����|� �PP��K�xlɱ�;��f�M �N}|�¥]�v����v�&����|k6s��㣣�|.�̸�}Ve떭��i]۳�J:��C�cP�T��Ȫr���Yy��0�����O�E}�˹��)7c~�۶6�utaFCtC|��g!�8����O��O���{��F��+�V�Ӗq ��B� *�c����yB��zUr%o޲u�ж�b2��y��mm�b9�N��N��%�	+�v
}@u���P���%�zxӦMSS��d�gql앯��������sˋ���U�V�^2��z�x<�W�����K�m$�l9u(��kc[�e�|
XKx	�3f'�/^������ve31IcZ�Mb@��Q}��8f`��g�9B����k"��1��}�<�hŠ5��Ʈ5��J!�B`��Y�bא��~���7�lj��UײW��v��[H�q�1,������rt��y���7������U���A�H:V[�~2�����T�pW�P��
�g�W%��P��M�V(S�G���;Ϟ?+��� k0��c?~��5�Rq�J�,)�u����� ���Cɖ��CX|��gh�-�56.J���J�`� �-sttTx�U�ZZ[+岯:"��#A���ش��3g��$� $I릦
�2�+M\ X�P�bL4 �)�`��W�'�n�\��SV�,)���ܲ8u}����I6'�� �����BcF/�p5;C����F���*P��&v������#%Yp������"c�;* �-�2��#�dÔ|�Z�x*M�e�� $���)j�/��.[��?����(^���Is����~���n������e>���Z�������]�ЍZ�>fg��Xsa��>�N=�(,�!|.Y'9٭(�f�?�(Pt;��!gp�ƍ[�a�w�>��)W�^�U~�D<Q�D�pPT?#�)�d�u��a�ߺur��,.Ṁ8�`�b�G�0|�w������|cv��ܲ�W,Σ|��V�t!����ވX�3�Պ�{{�SMjL($P��k�6�Q�o~��B#�(7	�A�^���y艚�|*�$4�����^,<~�!:�ҥK���EP.$[t�6,��b�1�3������#vz�_w�X�[���,֎���婽  ݱ�ѱ�- �X�����$�ʡ�VCs� �6lfԨ�`�QCK���h>?ZԳ��'����mUvը�+�t���G̼�6�����x^�J[夫C��S��O�3�E頝R��f{L��d�:bQvD� V� �\�A���B��U��|:��!p)?X'\L|�3EI.���Č�v��w�����_秧w�ڵ07�3x2�q�M[s˦� �+W�`���@x�-�l>��'��{����@-�z�pႰ����u�#�H���#��R���g||�Q�b�>�b!&>�����Yo����/��Wr��-[��W�%ȑ,@؍[7����
+�iONNww�*Ӣ�&^���	&PBIl�ਜ����$����Η�n<�w�.�I�uvw߼}{ay���n�P̱���A{t����������&���X)�P���'��Q� �u�_<���`ѩ_YQImK#�3�)�:��w�#�Ղ�cA\r6;v<��$^�h%өx"���a	��)/c��*P���Z�Y��T�o �Mٮj��1�����8E�Z��:����i-�Tu���~_`�m�H�`
��cԭ�B�?���k-u&(	��|����:���U��9
Y��ՠUt��A%��uѫT+�ݱl@���9��$L��R�}yvV؋nߺ%փ4���� Q�@_�'���ܚJuM�MM�/J�;62���\)U�$�b;�D�پw��Xկ���[wnJ���a�]�b�)��c��ɶ2��=�K����]���4q}��u�eB�)��Tf��ݨ��۷�mEC&'�QHGs�W^R�Ie q�VC"�,,*��y�_�*��|��cG��6;���c�P��e<S.h𢣋�ocQ�<��g�?�:ZL9���xsj|�)�t���vbiX^�c�M��r�9�&��� '�Pe�ĿԐ�aF2�ԁ$�����j�_A��{]]��W-�sϟ��hmmi�̋�O%�'��tмd9�/�ʉ� �`+�hsk(mEeB��51��m���A�	��E�Y�J�]Ceb�� ,$���jT�6'o=>#N���:}��+x�<�׋�ڽ��3al��̺���:df �F���t�uF���w���d���܃��B"\��x(Q�x2I������@����_�җ0��9=y�����ŋ�+
|Щ�-`��[�b� �aVK��r�OG������̙3?��������PȎ��7H����7o��� Q�ϐ����/~�)D}�F�Fe��s�$t���W_�vC�P ~R4cM�ҥS�lk*��Ro��U�����QT�L��]�r �*�v��
�;�����3Ϡ��G�E�<t`��q_e�<(�dVc�M�P�Q���9�ӊN�mE�*D�-���ZC`�4�q�*�RLe@��@�;*�{��:N�]ИKG�(|$��Ԛ	��ga[k��dMs���<Ǫ��F��yaG��%�)��ȍ?z�+� �3/h��Z	�ݵ��~��.i�=�'u�I[��\��(�OO@K���#M�	�\	�D�"#7�s�J6dW2��!$�|����Q	�T$D����Y������2e�Q� ti�s�.�ڊB&&&0���W��P�P���A\	��@:e�� � Q�lr�	蠒A�W*�w�_y��g�p���x�����jWe��ھ}��?N� �[�)�r��U�o������r vV ~�(������]]��,��h�l��O?�4ޫd:��@�P���	�����ٚRް���o���<�jsu���܅`��$?,��?�я�y�2�s�G�q�u�)�t���ͭ�֚�X+�Lơ�!�m���Q�6ίUZ��zgֱ���O}w�&�pE�x�`k%��ń �Ojc<�Q�Lv�TU��}���|�����Ps��o�����w��sH���d�W�x"U������P�����d:U�='�bz��Si1,廪�rP q3Ƈ��o�����1�,{������0�$�Sg;��*��ȵ�W1%��Ho�+ɿ::1��[o��3�_ȶ4C������~�X N�ر��(u��S�=W(�����;w�<u�4��7�� ���.IR	�\� vSS�{uۿ?)q�V흝p��_�f��*�Dm��7m��_��Z�(1�^��4m�ڵ�0MPR�+~[�FA�ܹ�c�6�# H\�_!�֓�p��%���H�w�+Q`G�0��0###: ��e��8�)Jjo[1npd��t6�\N�ܼ)D�Yq�c.�bcj�c��%���G<���M����K�K���֖�M���������*�8�}�PYkk;:���������.�h��5�Lz���Sx��y��z.���2��:vi�>љ���eFW'������uO4aY�z���
���Bp��0�2-��y�Ǳ���>����Wk�gi��Z����E>PǷ6�I�����g���$�1��D�P�N�z ��GƄD3&�'i'��\�=q-H�3K���r�T*{�֩���oP�����>�9Ӝ���3�a������t��*F:HZ�^���0g��D������rB &T�=̌~��%���遌����-,AC�1^x@$��m�H$�$SZ������];���ߌ5��_b�S�zn,���5eR�H߉ų����y!�D,�Ғߖ8S;W�~&nh����,|q�[f竑o��[u��xt����֝��˯�}=z��ɓ-M͛���j��>D�D�%�)��8�r3ͅfE�oS3�Q�Z
�н$�bu�p�L�
�T@��/B�5�Ύ�j|�P�9V&-۵�=������������L:���S�a ��e!~��"��U,َc�>z/���5wm�:��@���J��A���(;���\�����ˌ���P%�mYU�e��Ǟ����4�镁�B������,��3��
�]N�4�ݿց�~�#��G�X�E[��ԂC�DT�r	�,�sf��Nt�=U�����s�5O�;2�@�CM0�AJPyT,����Ie h2--�1���{��!��]]]�̤�G���!1�� ,�F����! A��.��o~��G��k�F�maaI<��0�qKoo/��*������BK?��c�lSOdwuw���	C��z�q@"@1|E�$�T{;S��*�%��-//ߺumGA�0��r�
p/�+��HL%]߀�pc8l���J~B�F܅k �$#��2 ח��e����c��Y*�r����7n�{��:u��d2"�������.bPE�-nam�*�	��y�&�@E�r���gQkD�h z��g �;;ځ���D�eh��N�P�:�Xlk�hZ>�l?��o1��F�q-m�u�;�֣�y�cu!�Kq��9��ɵ{�y�s/G<=h�J�O�4gMS*I+�R��L$
�]U_���،,�U�v��M����p�oӱ@�ҏr��2���� �\���������ߜ>}z��6��r�:�	�"d�8^~�e�v�S(|`� dD4�{w�q��eB���aQ,&�I�QT��
Sj��R�'�M���W����M�	�fTd�↵j˫�C��:5j��Bbk)	�u�
3"�X�*QeI�i������u�dƳc*�ԭ�W�?m���P����W+
��T�I��G:^�uǆ�ydC�|�-*Г��@����}�װ�5e�#Ӊ��mEB&[^��V�@�=JMeL�Ȕ��T�t=��5�j��@�`�b,��7r�s�<i��p�i�"����o���+WLm���G�lBp����@�D���|�&��k���6��W��Ô �I��U��PT�ռ�*d�D蕉��Ƞ��h�ŀ�����ĄT���IgW��T������������@f�R!�0�g�.`���QE,�z�Ϥ��<��|Lu��v5�5�$��W�>cV���رKY���691}q��b�<>/�@�&W�^-K4Σp����|��ГH�\.�
�T�so��G�5W�\y��� Q�-1���Tf��Q�D�T�"���[\��\.�G|�R�������"����߈��$UQ%u�Ν��aȬ�[�Z�*�ƎM��`2rcT�[�LNO(C��ʤ�Y�fA���<p��Ç�����r��Z}�m�-�����[& ���t;�϶���u�(�צ�@�㈠ʦ1�+�r�����[nkn���A�l'2�a�
]8�g��B:W�%	���ڎ�?�#�x���������(�Y�)P���z�*�n�L����۪�k?Tߘ�x8�����У���3��.�08ސF���
�%K5���o�h������$ӟH���m��s\Yw�'�W;���K)�B�խ<U�Ed|b������O�Tf�Y���BӦ�
!	q��hww/��djbTh�%�4�b�A`��-�*妖fT+� I��M�:t0���$�J��>r�����tgWWPuf����ܻ{�L%��S.T{��H@�x�Os���Q��	�]���~���b����M��K$+Eߎ�>|띏N}��L'S��}�Ͳ��5�R	�ce_R�eR1��~�UWV~�n�. EEOyDl4&Y�Ս�6=2�"�V��Ǐ��yt���^(1���^e|�މ�ޙ��&�؁������@��Kj��FU |.�$0u(���ڣ%�&b�+@��t�L�Y��e�m~
�5����}�5����j<�$�F8R/sʄ&-�����T�6�E���ͺ~u��a��zG�"S��JO�s��#��GD/*���3n��#$�ʵ���X���������ьX (���	��ƀ&��o�
ԙ3g���^x�%�\(vǎ(�&3�~ڶm��믿�Ҁ3$0Ӳ�l���c�ɔ(����)(WB�|�2n?x� J��鱦g��={��<�X���*����b.)�pcOoWD�������\���+ 
���E�}T�.��ࡤ^�Am!�:;Ł��U�0��F-�at*�������Juʍŀ� "�C[�h�e�v�Uō�\Do�&Q��{�����d�j�s��\>����@���[�����+ÃpI��?�͍N��*�<����̤��"�*+ *3�l����L���Tá�7n�5Ԣp�����=��7ך&q��{v러;c���k���z��F�p��>P5������K{P�CM�������FfUu}��D��ʐ:
jJ�A<L�9�&2l��N�j5q!��Σ�t�?Q�^iZȲMM=��|��`�>��,f�8�@C�\�p!+�=.Tj]��ݾ}2����������Zq��Ԥړ���_���m������Xի�U�ܔJX2��:�;6��,�Rj�Rָ{�ޫ�`
NG�A���[+<�}��E�$�	%�Z<�0?�ں�w��I���?�G�{�MYnA[�ߠ���RqM�ţ��'JN;+�� ��?1��\��u�38KEwQ��)��x���O?����������e����:��ر�:V+-|�|�d�Z6��
ɏ���Y��=_��l��r�N��5�֍O4����l��9��q��56V�R�[�$ګ1X�0�ފ�~Q%��L�w�*��\*aert-4��|]?�lv�j�u ��R�Tv�d,�+o��p ��,�N�*��BQfiU��&�jP������W�20cgW{`����ʎ^s��(nٺ���?+�KǏ?q�=�R�8F�ݻ��7߼|��E*��)�9��{������q/�9��!# _Ć��E��$�P8��{�o05��vp{����119��*�!��jn�8�)���I��6C!�������\kG;io����^{�5ٌ���٥�D�%��Ν;��-4
�e����)!���Wa��ݝ$��Գ�w��^+쩄�7n�@9-/��@K��<�������-�i2�\@��x�}�����@��Ɂ"�p*���2�g�9�Ҥ���SNc&VO��B�|�`�m�ہ�����!�4�tS�$�%���������*:��4j����'�����T���g3�����Ύ��g�ڑ�mW���]ZX\^\�vue]RJz}��Ϲ����}q�:X����0�T�����)c�Q�ieYu�o�ekݻ�u�{�6x<4t��Gc����x_u^h����<P%h������s��{�ܦѥ\��%�҂�W�
�`�R�KbV��-������#>�[���}%[�x$�I��+���K�͎ىt����9��5���+:t������oSP_]wT�q!ש�]���&�ss��H�!� �J%���v�W}����_x�Y�(	�ť(���e�XS��<?;=�ٔ�ֿ�����xiq�V	��T���\�\�,\D3�e!KB��*�l\�:6y�W�*e$���Z����Ξ>������W��% ���x�w~�wR�U	��"�U�R1�p�W\k��#g,^��UD���xwt�FR���&檃�7芴��6VE_]�q�7���֒vl�C�%q�P��Tok��c����� ��E
��5rzG���&��Θ���Q����)��0�qBg6��2���4�#��F�����)�7�핚�,+*�9�����tw�Rɼڋ2/Y������%O��. %��T��JIF_"�v;�(�k��a~��-ZV�j���VUX@����eOSe¤�g�(��bL�e��G49B���f��g?���S�|��aV�l��|Әa� XX�Ν�z/֚d�W�� £�P5=��u�]�-[� u��[�t���K�.)��lW�����b������ť��ѣx��ӧ_x��s
�dPԄH�׮]C�QLN��=��jP�]�T:���P%4ARtv�n@r(�	�&Z��P����)¨X�}��������'�D�W�4�rP%6��SJԠt��a����L���bܤ`�S�q����]]]b��%8g�J� O$b�����_�,T�������?�*�C��H�55HZy9�i����J*)�O% E&�F������j�[1Uש��Wk6g����:�������<���H.���8�����mj�;To G�J���s����$W��{D��ݷo�gVe�R���"@��ZB�Z�b`�/������`�6?��Zf� 5 BU�Q�T*վ/����{�����ﳸ{xl�ݗ��q�T���Ƿs>?~�my,"k3#�5�����P�sD~ �Sh��z�Q�8���+� J[��j�U*���4�^m����f X W�ԧ>���O{�ێ�;r� _u��Q��������u�>�Zi������� �7\\ZBF755jm6fg_��������3�<���@mfѳ� �b<��~���䈛=Y��"]��93������F�"�D6��Ta�sý�l��
��{4z�?0��qq�;��	����j��#����:��`��d���pX|�Б���_|����������^�V�ψC��"�菳�jTp�Y����F�VJ�����dk3�/<T�3�XB)���OH�*@��dԊe�D�q���ri���E�KhW�n��?-����~ϱ���*"�+'&v�Y�����3�3ƴ��"Nٻ�*��qM/l� �����`V�p�!<c��շmMd��p�Q�ޕ���{8Î���o������s�3o�<�o�<��#�^r>���@�'��/_>v��s�Е��ʕ�5��	�S\)�@d��}mffJ;t� 0�������w��3�s�Z߸���R��$x)�F�~�ee�qc��J~�> (���V�~ux���
L,�!��@F��]� s����<���CC���s����7g��)_�0�-:��m��C�^;�:�����G���p:��[�[�܈)�&�C������C�)
�;37ˡ�R�a4���g��j4+����8�=G8�gkq�G�P��CZ�{]@�0F4Q��Ņ~�8�����0������rHEAs�jxp��vb@"fr
Z�l:3�kD �}e��Hy��qI%vcWS�Y�ΆO�BJQd�P����G�&�NeX�[����u�����D'�S���Y�$��9��Z�ƍmw�� ��>�� ��@�9�ό�^���ga�*?�4��*J���� }.�0�o���}�&�0u�s��E` �X�8�-���}�� 5�w����7 ���?\�G?~�E��`#;w����������=��#��w��Re�Q`-�ݍK�إ�F���O^9s��g�X���m��~񹕃�ssb4ܸreqey��y~��j�^�׭7 ����
Xk��mVaHR��j���z뭍���S��{��}����h}�+_y�|���������A����$���-ωh�(����r��;�� oG����d��L-��FQ����;w����{�f����� ����:��4#YT�5a��_����!��h�/ܭZc�TM]&�`H0n�H�Ye�������������9vش�n�tf�"�I8,�;"B߮e���������k/�%p�8)�>��]|'��wabqt3F���e�E٦�v�5k Zqg�q!�S<WXZlOƗy�Ʒ8����߻D}^�1�gf�yn�\ߦ4;7���������.�ǝ������!5�bEh��n��?x%xp��� �`+&)\Td�~��l�;���ٟ�t��w���Lth5 ��y�E���1��3 ;�G�����~�w�o�[�����������&t±w`L��0������������z���_}�U ucs`ʑ#G���_z zq{�G�����+�= �/ί�-�*�ٯ~��P�p�w��?��?��%𥁅�Ev���O(�M	�Ʊ8�|���L��9 �����3��!�

9a�8ph2��cDľ�����c̈́Q-�t�mǠ~,{ꩧس�k��J�W����|��k�q9��j1��P�*����gC76���ڲVe5�g^�v��bǢ�x�����&ndz+��1�}i����'#D',���K�[���a���d���Zw�*j�Fh�3s��&�5�6����Qۄk�e���1g`-;?��Y�:v��k��o}�[�����v��C>��/���8,j`��9d��K��_���_�^���Ϫ���������lujjkm��ҕ��/~� )����CQ���z�����'?Y�Ԁ]/,�}����A�..^{���'��Tc0߾={<�h��%}�V�j��°�q��{�/�8��z��?��_���F��h�D��M�AA�>J�Q4�+C[�e�(]9ˈ��G�ˡ�A�@'�3��侊��z~��	̮ �O�������~���u�-���]6}yq��	������ng�)�R�$"��d�P�(�p�#���Ƌ*���-r'-#�m(�<����)Ǚ�r|�\�:��3<z&i����y}dPC{ �
�"Ǩ���91�!�l���x)�8 ��6���o���5|Bu�1�Mَ�bLn{�W�}E���̱{��U�#��!}t�T`;�7��~�j!��3�͐�6��=��v�QG���ShX�j_�ھ�p?�gϞnw�����ۛh5;�����������6Z�ê�뮻�����¹sw�y�W����{��{���t_~�����O���~�ٜ��O|�{��k�O�|��IK�r��� ,!��Yo�*>q���|�?�QXґ���Um����d��N�ܯ���ol���?+9;�5N7fϽya�ŨJ0�N�|�#�(����心yˑ�3S3�o9��Ϟ8~�Z�?����remyu������E�)<9�^��ٳ���[[w��.��[��.�/�-�"���Et����{��,,�9�f4��n�MgN��GÃ�g^ :?3���\��xjv�7��O�>3Uo8p�{��;^��ڔ*�����������̛�� ���o� �CI!�z}*�b� T��vzx.��/@s��VV� ګ��f��Bu�䙍K��j��;�p�~9�&�������g���z��l����W��!L���H��p~qh �V�UEu���j��N7�o�j�����v}c��bt`�W�r��,��?3��8.�k��܊��V�gڿ6���s�E���Q��q�s,���x�`��'�R�v�mb��	��5<�c;
�r8�H�q3p\�ҁ[1�������)l��=��_�Q]֗��&$�㱪��J{��ba�С��F�1�G�v��6ySZo�b�Qs��ހ{���k&ڜ	�m0���x{ZS�!aH�ҡ�x:�XL������6��E�tm����+u�<D����� p��gބm����S�Q����/��(�w�wآ�YYe������t�97��\[��܊z��_x�η����O�l�ac�h߾= ������df��'�h�?�ѣ�b�?����s�̀��~����w�`{��;o9�W��51M�����# /�8u
�ȡX	;���!���P�>v:[�F�3Z
m���o���/|��|�� ;j����z«9��03���7A��MF����=��3��K��x�"E<T�6`m���|�����tS�e�@Ȍ7���H��LA��hVE��O��E�54Di�>����˝+o.,�|k>���˫K���lnn��ػ@j�	�^�������X��6��x�=��6���w"e��V{��C��=��Y!��#�&<��;��Z��:6\΁ƚ ��MQ���
8�B��xd7E�����m%�>����J�0f��شR���YM� �aO2R��8�qB�:e���W�ĳ�Kd���U`j�,T�>��N�r~�H�O��}�q Ȕ� �+�X�f�m���O��>{�ā�!Ct:#/`�<��fI�&��Rz�c/x�{ �{�(�9%��J�����k܇�z���ȑ#���':��/f
,ˍ����˿|�;�O� ���o~�F�C�,-�a���/s�r ��sϩS�^y����ĩ� /SS���'O��ȯ=��Ç�H��+�����U��O;v�B{D���_���}/�N���۷�8����÷|���^^}�ĉ?��?}�m�}�K_��v���o {"'=�)�[ vE<������M'|yػ7�M����%�O>�|��a�Ut��S�YF}�	{��0die(��O>�$��ٯ�3D ����0�p�>��)-;E���2�=���Ю����:���#��Gp���vW��΄�@�
6ʰ�}�g�������V�]__���K/<��#� y{���_���i�D2�C�~�����Ge������gCo�4ӌ�;�� �^:>�����&!C:V&�c����(�ܾ�W7���v|�eɎ��p��H�$�d����^���˗�u��ߣ;[x F��&�eiF�&&�1Y{s8p]��{��^Gםl&� ��(P�<�|���O��5����/����wA���Q@6��C�؃&,k����Y���K�AW4x���7趷��q4��
<�LO���SO�;x J����hr����v�4S ~�a�y��b b�̽{��. ��-�e�#HF�y��=���AĬ,཮�&j��\�ϵ�vQ,���v>CQ�
�@�Rj�x�� @`���!0G`�hQ����8���2⍋.'��z�)���>�o���NKd�o����CO{�ym��C:�vR�u�6Ą�8rLw�H��{<'�?�{'D�ǈJ9x�ٟ(�	,s�C��dk�2�����d�$M4��o����O��ہtO6�q,��X�W\�\)3^w���[���\��1�z�Kl����9��Q~��l�F���P����`���X�@`��1C?���d^imw;������e
1�|�������zࡇ���G������ �̝w���{��髟��������uϾ}�{��sg/|�����>ФZ��>}fyeϳ�<�������~����g��8�l>���:/����	�r��yhN�(^^Y@ πc~���-�j�z5�/^<Ϸ>ad�����g?�k����?��o�=��c0�o�z�҅sO����� -���¥+o{�}���ط��چ��`���$��F��n�|����p�rp�x�`����x�W �A[��r��_�a�*`��/���,-�������n�4�D���.]�x��gg��<!����Μ;�|�}�{/ �˗/�۷�|��w��$���jC���/_a���	hP2ߢ�彺�G'N`�,�a�.�nQ�������~�|m~�4��n�͖�sU;�4jCs�:��!���D�\>���	e���#6J�y5i���:4����.'������e�o�gQ�]��7W���t79�ԓ���{ˎ\���
n<��]W��&�IN6w r�l����.��,��ϞW�;�i��?�֨�D���9}�tR$����CO?�q�V��|o�y���>�����4 �]�G]�U |��#��;���������,�C��u���9Eޭ��Օe@��{�ێa�����Yr����Am��^�
j������fo�P&�(��B]�smc3x�����*H0����/|��FT��%A�����z��Cju����l�����Q��у�����!��o�r��k�����Ǩ'Ѓ�	���N``Pڐ,��
AUl8·W�-���G�������;ݍ��;���4������I�%�Mu�y��bchxY��3�XDv�r�q�c,6�bJP�ӽ�0�����,�w%2�iF`b��m"y�dR��x�������]J�V����R��ׯ*�v��2Is��^�L�MQd���D.D����r��a�PC_��$`:��/��]>s�CȾL��fLw��Z�p���dʇ�&΍�=��B�#�ǆg�ҡ�eVf2������/^-���K@�3�<K�3���?��?����O��,(��w��=�:++{����#��ZX����}��w�����~	6Y�G$�F�5�x)i4Z__�������v�m/\b�
@~�ֱ�E�������p8�V+����7��:u��?�1���nV�1/��@
`FgϞ�������o{�۾�o�۷o/�2�E{�ԩ���K](������۷ϘX����'�䷿����P )����]Ԟ?�D+1J�+��h�-�P!ZH�z��g|�|�ᇀ�h�ʺrla@���P�4�Ä!�r�>����(�`(���#G� ��~��������(��/��į����E=w�G� ��a�(Tt�J͊_es���a^2׈��1�ʩ���K��e��f�Y�	oۢB��>��tw��F���X�,sFgf�7f(��ez�]��v|���c�@4�q��+o_۔�N�q���������%25V|�^Z�lgC.��}����5��Ņ%���W)���U6-值"|t�?;?�C����3���� �Ҝ��O6rg�T��F�\�"2���z���\\�w:����>0U���{�k�d��g��f��!K_TF�o"{������"Z�q:A��z�6߾�x6k��d8��bۭ�����w����	u�]w-/b�\�x	��<d�ވ�9EM">}#L#�,����<��})X)Ȏ�Y(C���{�#�g>to/��fll��J�x��:����/�z�u&.�r[x�#bE`R�a�
͗|��kkp$�v`��ܦr��L�gB���9��������$N�7�'{Mj�RU��k�LXˤ|����җlܤ�z��*�^���UR�?���@�����=��cT
��a��]�nq_c�@n�<������
�jy4E4������x���Eh���GPQ�i���|�x(E �r�{��M��W.��|�� ���W��7?���������_�? �Ꮋ��~�ܹ�G���-����ã0^Y�3���<r��E�����{衇`��ʧ?;*������菾��7^|��A�.�!8�z�É�y��0�a���
�N�� ���W^}i}��'��;v/��������B9u���*�!���С��^g���������¸�n\��>?��>����g�zrcm���0w�ѣ���[[���^�EÁ_�����;�S��o�}��Ǡ-�Ν�9�=��m��[�+�����:�����w����?���s���t��:^]F=%�?����F�Ё}����lCO�Φ�1������3xs�x���f��}�[�+��+0� ��5�߷f
nCG����J��{�6k�>��{��[��_�n�S��V/��@>�EP�b��A����j�W��n-.�7����0�]8?���)ٙ�ys��ȋcXC�Ner�o3[�=.��vg�l7:��$��r�g�W�./N�aR`������I�?��'�d�e��I���3������ki~}m8����+u���m���̱��8���<�	{v���b�&�?��n?��ݣ��V� b�& r9���E�2l�O����{�%��{���m?�����X ��|�q����������C��OQ��JՇ7�i�#�k�f]�:���M]^�B����g�
�p��Y�^:m4���P |;�֯�h�R�u�66�\b2�V�GÞ�g �7�V���vg���Fq�}Uk>���Gʑ/�FՠZ2OB!S�T��lB@����⹩:Y�t�"B@:��!�t4r���M��bܓO�B�烰K13�v{��q�.�x�4��B��T��D^n��-D*q�Z���g-l��=�����.>�	i.@H�����Z�[P���Ykv�+Ʌnj�h���1h+�L�����m ���ҡ!�l�\,}�$����5�����ڌ�fl6f"��_+����
��m��a�P�C��	�c#=_��O*�v�&��&������m]��@�*�`X�r����_~�K_�ҁÇ>����}�=�>�h�ۇ��/��Z���d���O�K��M7��_IRA�=wm� �x��'~�:����9}�+�9�$�t�����1�����C��|��{�{vv.��I7
a�&)�)mh�a��os���0
ʅK��u}}knn��/.CQ'N� �p�ԩ�~�������K���x�x%Ƕ��t+[b�y�VWW�g~�W^a�(�b�k섂�4�
�iH�� 3A��Whcw�0[�A�|���ǨYg޼��[�HC���v�P<��Z45��;�]�%ZvحQ��w��s�T��wK�4(�=�y�������,-����:P��O,,�+5��_��W��6�) �����W�	��շ��,XphQ�t�]I/���@�l{��[�>M"�EFx_^�`�3r����ܸ�Q,9L.ΰ�P��dU��r�}va��ܼ�e����=����bU��e՜��K�ls\%|&M�H��9ӱ�/� �Vh�*l�,�����O� ��<dS� 7@�At���)�J�e
^o��D�ml(���c��-@(;9b9���gO=×p�6$��J`�{�ҥ�t�����s��W �7*�>@ b�J��ӮM�lT�g|�@�b��%��P/���&���S�/`4���A�P{�g�l���gE���
�����h��I��Zx��5�>��;j�qI%'����9����3�a_5.��dQL0��w�駝!(�)�x)lh��g�.��#yz��������@`d���vz�c0�Pq��rQS�W���l�Hz�g��h!GYuE	<eX�lV�͔�9��ǽ@�}���Ӱ�G�oP�{��������(�C��0���10׻�>eCu]�V'KvT�$�3:�����J�cO!��ڂB����J��i��(/R]@�Z������N��$Q������w����~���8@1�s ������ J����@�1 {������������o���8q.,�����y�!h��/��ʘ����˸y�OE�>�Hu:�o��A�՗�m���Ӎ��wNOOU��Z��]�K� ������֛��f���_o�����=�W�W��ϭm�>�6m��g�*T��l}�#���SO=����������g���Ο�����)
}7t?��\<{艣Ѡ�]k6a���o>�w��[.\<w�C�̧�~:���|��W=�{��ag��U������TF`ey��g�����������[_x�~w�� �C�����M�5����s�����^s���҂���갊��Sd�wk���W�z<0��ܹ���:|�=��<q��{�}����������Ź8��YY����?���o�x'E�8�֐�l��^Ǫ������D�X�����v�~%bȀ��>�l��`$ʓJ�4B��&�m�e����i������s�I��%[kQu������9�*�R�ǲ�q�t���;�a�t�.ep���L�9�o�֞��Ei�}�XL�{����+���pL��?F�ŧJ�,�-ɿ�2v/|��7�;�5[�R�#����Vk-���/p� ��G]�VGݰ��n���a�G�A[�s=�%�Lll�倲3�S�p�W�vױB��>� ib�*����Oͩa8�ƶ�m�ա������
ikc{a_�ý{0��`��l��?��>I�I"Ə"k|N�@L�3����XG;N5����>����q��_2�N�J�M!F�1�e}����no'd�q�����t* t8���0�QEaP�����A� �&fФ�T2i��0�fe������H��,v:)��������\&��%�z�T�"֑Z&E�N+���>���a���]�Aa�����r��*?�h�3l]M�=�d�%���(�X� ء�4�աX�2Ş߇�w�
��+<����`�m2�Þb�Q��;T |��j�2���0�������(�z������>m���\s��i6k���ۀ�5ּ��;��^Vn	:&g�� #`��Y��P����<p�"jq>���|��_^\Z���>�T�~������� �q�]w�8q�%���;d�=�޶�ux����&����U�F�@���_�+�ܷo����u Q⡇����G.U��k0��޽�ly�̅���M�Bv���}��ѽ���K�`�	�����|��#G���OC�0���-=|�0 K �M����!`P��q0q��I>jd#}����K�kY�"�C�G)���_�={a}�����	���t	!�/�8�WWW[����,�a�r�vf�N�Xz�U5������G?��3g�l��AK�AӮ���={�\�e^Y���`a����ח�Ma�qf�n������g(J�����^v�L���݄���er]�+u�^�d�^V�{3�mu^�T��<W���se�d�uU���l̽�_`hiԨs�\����m�B��%��W��06b�H}�E;E��6<j6g�)�>��=ǉ䴸���N
'V�K:Kb8�+�^�Y��Ƌ���+]��ᑷ�����^�E�]��S45���nGR��0�u�8��fg�c�>}J;p� �A���E�	���#�y#�g���*ܙ�R.��<hgV�.P�Fjx��t(�7	3!��X���};���L���8�#����X��úD�Z�s� t���E<^|��j?�1���d�'w5�P���f�(ϧ���P�CM2�6ƙ�'��"ş�����ӰO����c}�,��d+�����v��1��s���C�!�JYc��M�b�3��o�M������?�Z|O;|������N�����o^�ݻ�:HJ>��~duLM������O�l�5�Y��~BΞ{[�6,�)�W��S'ވ�RI�= v���*� �2�/����#��Vo@���� ����;a$�hIMI
:-U/>��ϾB�"x���%�g N;th��Ę��~�gQ��m�q�m���o9�1�������_>q��IX����j� O\�xp�����/��X���z3S�=+K�vk��Xnn�����.�ӟ��w�;;3�S�acسg�����p�#x��w��Ϝ?�X'��a�w��wøPX���B �ܿ����}�<����ʕ�n��h<�@���{����������S������a�gw�}�=w�l!���ޠ�e.s��!�F�ʶ���c��E\�k�a�G$0������.�_�(�fg�Ɉ�P�2{eT4!�Ѽ*<�ǎ�u�F_������6�B�(�n�6C�q�*>��^�R�.]j6�|2*%�\�`�9�e׶���S���_�eW�E+��L_B%[M�0�=c��-���{M7���8$��l�R[�	��3~tǀ��ƺpX'' �����Q��0�y�⦼`��S6j�O����T�iG25B�*_��a܋z=��3	�ÑS5�I�8�/aK ���))��m�[n��^�n��icc�xN�K�q��՞q/�G�G���_%����Df8���;v�[�A���Knr�q+�s��ezj0���*���033��ڂ|�~=�Ũ�xd��^��KVڰO�FѨU��J����@��I��d�$d8�?)�~o ��[vqE��K�wJ�s27܃2`�xB5"�V ����/�h��/�<r�_G��tO�ˈ����P���:��U��h0�\��@�R�.�F*laE�E��D-���W��ъ9����=�L�	pPP�'S챈��2�(�Bz��x&�=��|�l�k*9N��k���Ҫ�8*�t,��}g2�dS3>�?H�y��Zk� V�/��Ut�P�� ��<���T�5T������t�I�и��7�t��e8"����'(��~e�$���%�+,�ˌ�@��<{yay�$��c��0����>o9�^� ��u�]�Rh5@1��"�߫��ЬJ��t��۷2t]���������4;�	@gya���_��O}�S R�j���W�L�i���-Z�b?�����v�"�u��9�w����~4�E z��+�,,-������?��� x:��Y��k���B�˼m̄����Q��g2�U�5*�������*%n���)L2>�v�̾�;�,x�B�)��9�b�M��HP��)�ۣͽ �����ύ�WOB�@�QmU��õ�{������먴�	���
w�����t¤�����w���^]ڱ^�K�4��B���|r%�2&n�v;�c�p�����g�s����*�k���.�/އX*N�z���qAϸ���Sa��Bt�c�$9s�$FcfQF���`H��]v��A9gٜ<��B�QЖ�N|)�%�����'���>��(��<�G����c�9�Z��9�VZ�Vk6��c�G}Q����N��d/	�$S��E������i>�fM/����6)xa�|C��(�{C���ޫQ�R,+��:&G���k+d�> Ȏ�;������+�`g(�� \��-@�J/+r�L<(g��p�b��ƴu��*j6S����M���&������)���V�J��?<zdD�����lmmml��,/����	eB���*SS�6��b0\_[��D;� ظ|�A~�HY�"8tp������Kqa�^�Tq뭷D�Q�מ��ū�feI���~/�a���7��3x�]��Y�ei��;���7`��/
� ����k����U`ܠ��.9|Z��l#4���*QG1o@Q�f�m8�Ҩ����|q�g�%��*,�V	���5���.�0"��Q,-�'2"�? ���d����2��3k�U��p�k�5�r��KTjc"u�iGLc��
�L��9L��@��ɲ����߱�BMյ�y��[�+&*�>��S�9+4=
CA+W�E3K>�����O>] �)�����ha�sd�$��'��5~�*߁t��6�9�̜s%g�ExS�ܮSB#�D�g��fS��7�V�R���bU�j�)�հR�R�\\����V�(hA9��)q:?i���ݩ"N4�R)�ؖ�'d�\�O�] �	����WJK/�y
�_���/Ӳݎ��Kr�1��aܦ��3S3����Z��XT|�X��-� � �ȷ/��0@���333҄�b�
��w:�V�p�N�C��0&m\�, j���(F��*��x�!� �*t*�'k6<K��'^��J{��c�L}��O�a�C{e�ӡʪk�����	{�x���E�
�"�\���Ǝ�����%����)�(��/���G�.\X\\�_��g�hi�����6�8�Śc�f��&G�qa��>C��vL�ʮ\��m9s����ÇO��A �.va͠�����׋�2��$*w���:� h�0>�����)d�������L��@�XP�=CQέ�:����䌬���EpG{k>�bk	kMap��[H�j�U�vӜ�^��g`��H,���Z�l��v�h;�<����e�Jm���J��Zܟ
	�}>F��6>��-k��+�2��&JʜmjǍ�t�g�ξ��L�*P(:=L�̅ 4��yvG0Sḯ͙'3V)�&�6+#�\
��>�؝�[B*�3g��N���t�n��+%xS�G���Ʒ�l��<]BI~A�s#�ƭ�A�W�v��YԐ|K�/i</J.@���������O��h����̲��<D�^h�utr�,�O��)��m�����pƿZ`�-�Y9�j��+��(F0�Q~I�_�[ԎD!ŏ�+^e@���E�����]|K���6{�&G��A��0�w�k��^
�'����7���T��^��+�^�U��;8C`�pدx��*~�Ru���7	�O�j��S���֦����hB{��_�9aX�ӨAN�f5���}��s��,--����tSmG��k�~g�Q��Z���M���z���B(��	���FC�E1@�F��koG%�Ф�LX-���i}Z�)"i�I�V��k�b�T��
��k+!_���bڀ(s��NwY(6G���UT����f�3���=5���;�	m0U��YVwY޸D���q7���|����]�5)U�sJB��9��i�b!�,��� S��1�,�]WW����[f&���W�ԁ�������D%K#��]&�������Ƣ*?c�..�>�H�'=���u�ei��WI{eR��h�r���q
IֻC�p��z9�G)F��/����X'�ό�v�,����E���zkg7x:��Nd(��un�&iDhZ��la,��IC��+Q�g^���f;�I��/��� �<�Y&N��u��hVC&E6c*����o�?��[�=�!s�©�cl��\1��P1���	�c#����l}"	��H�3J�c�F�%V\i�	��@2�i�$)���０;�V�h|��1� ��޽�M�06*�Mv�6��u�t6H�ܹ[���)��P�FQ�d�n�����3h���Z'����<<��6Z�W�:�\d�7(�Aq����u	����ߚ���)(���� ?F#���7�1p��&�2�j�� ���U8I����Gy��68�H+���=vY1׈=D�<�Щc4 \O�ұ����E��Xӹ�2���#x��2e����5��1�B��:wuؽ�xk�	�H&��ve�I���i��T�����MR�[���.t�q�7z^E	e�e������]y����Z��hʴ2CY�n0�[W�E�B*�'#���e��H�e��Tr��wD�</u>+�!�K%3'Uz�	g\

ɩ��d���r<7���V���톪�@i6X�r�<_�nyQ�s�Pl�R�-?�4���]0�	�&>҄��kO�X�����s� (|�����|}���*^b�s� =q:�f�<���[!|ȷ|�>)�0 y�ǝ�5�˚���WkJ9���
�*�8�+*���B%�[�x�0lb���,�[�|l��a4$�%?ī�B� ��(��"F� ��CG���yo����������Ⱦ�f؍nnn2x�@y�g�w�PZ�Dw|�t�R�(B<���y�0 Ƙ߳ͩ+���T���_	� :�EW`�5==�����Td�9�G}����Gz�h

qF
4@��{D��b�<c� 6�x��"���7��F
��������#��S��v2[t.�2�#j��Coɪg����˱�	q�dUN�쮗kOʀϫ+p̢b����#2�L��<#�M�e��l	'*����fB\�c*�<~4�K�.I��!�{u|W�yG�(��4
�d��<Q�t�R���������hѤLya��#��L��-�Ѣ��W��Tr����#�ļ�]M��s'�������9&lZ�H,�濋w��ԟ��yR������i/kR��R�^������8O��guF���'�T>K��؎��z6�EʦhG�td3ӿ�3�I�2�%�(wje���2�,�1.r�3��ʶ,(�.�̃�^~���=�y&=���7�sO���z&6�6j��[���7�M)�[�S,0hDR;͟,_�Ņ֧3�W��ڠR��~j�Y/�B]�xUj�"B9�(jcccvv�T��g���(��`%Z�h�T�!!Wt�L���2��|���3~��	��H�e�� ���i���l�=����v��Ap���(�������z[!�9�:�m�%9�!#?h���� `���p�AF����*���im�YkI)�]�����"7��gv�稵'��3����54�uiI���D1Hk�܋�R��)˻�t/�3�g���c��	EK���K�}�uG?ט��Q�ey��N��nKeN6���%v�Әz��f��.�ߝ$_��{�������2[x	�(��GP�~��)Dv�QT��}Qa�b�l�퓼�Τ�љ|�ݽk���.=j���y��M����%c-�ΨL���[x��F�۵v�	stQ
�MH��xˀg�S
?��� Ώ!o<�-��@�F�xs}[B�u�"����H��`DGA���6j�����?�-Kh6�V<����)v��A�����^���(�U�x���pg����rT�Ui���H���=)�'���^������DQX��M�U�h����4�G���ڌ�ތF�"j��Cw#��
|>3ӄ/�}����yUo���a<ԃ�8a��F��otg&�D��2�j0T��G��J)�U�MU�qDUx} ���nk�Y�V��,�5A[;5�OX�[{��6��كF��צ�o��xQ(�ҸJ�	iI�9�}�䆊z�'5w9��.�dt\��=�G� ��j�\�)\�98<!cf�^�2�t���fٟ�TN��b�e�l�Cߒ�ΰ*�9#�Ŀz6٭r�"��|M�,60al�.��&�KW�k{��X}��K�t
�;O$�����ʌ�&&��K*9%�e�,��UbdZȸsծ�$(MZ�GlhP��:S�-R�O2�����W�S�T���}��h-��j�=�3��=�Sh˭q��h��W����8�������K��{f��XDi�,���<�v/Kb�i���F�٫�n6����>X��<�J�I�D��'�׈���(2/���rz��y����8�7:<3�uK5ص��R���-�M5�iQ1��=�YzxD�����ֳ*�x����;ƚ~��X�C!��2�xn���$�����0TF%P����b
��ȧ����2�σ2~��*8�i1�a;#+��*J�m��WO[x��U�fMc-�\9�FX�Z���:��`7J �����l^��)/{i��J�s]D��^rW2P��'�r�pel��F$i�x1��"�����,��(���,�0c�, F�&��5��7��r�x�T֙o�4~_ǶآФT(;!�:u%�))�:�o���6���w�,�c{/�ƫ�3���H�~ڡ����
�t?qv�8g\Qx�]K�Ȉ�.&O�@��q\t�pzd�d�������ސf/X�ͤ�lv�P�j��%��8�T�y����J�12/3_�=�9�Lڠ��ҥ��߅wM]��8�l�]�1~N�AL�҇eξV�2pA��`e~���#�
�QBa	>�_��O��d8x��M�w����_��ώ��23)�o2��`�c����~�W�$3�qxw�4��ߜ�ԯ��i�PO�7�?��J�H����&
6qU��+X�d�W�!�9Z/���e�1��'G�����3����)��ٛ�i�Dd�^Q��[J���Y�HOi�#Dyg>����4	��A�9�ɛ7�M�E[�h��O�P����ǈ��W�����?���x�\�fl���UJdA��`CciR��ϊ:"��EH� V��(�N�$Q�f6����C�fο�9�'�:}Z5���<
�0���
�SF&�8E�%Ս����bl��kEz��Q�p�8�95���o�m��ҴH�z��u��2��<�l[�7�7��q]�Ks�\�0a*���a7\�vN�d�+`�[H�(m��xd�u��2���g()���9?E2e�'C�f��%��N�aw���E���9�k�-+��c+59S�[�Z�c�bl��g�4mٜ��g���21�o�
�!&��o)N�+0�y�X(k�z;3�2�ǳj�}�|咔z���-�)�_S��� W칐���g����dI� V�%�/ωClj�q�lT�1���t��ɴ"���V�3Vaj�	��I����pj,���k�r�-X��OH��
�>��4I%g�ɝ_u�uRP�r�ʐ�t!T]V#e�Lz^h\�����rW}F?�`�Vd���9l���]���IC����>�4"�iΈM�k���FK�\L�8�2d��#K�'Kv~yf��?�QPw\��kt��heu���G�Oe����W�N5�2�Y6j�0B���+�cZ�[�i"2}���E2^���ҟZ�2� e������@��gȓ���*��e�l<\Z,RB�����V8V�����f΀��,���WT�,�a�S���z��̜$\/�[�C�ͺ�E}�Z]%_&�9��bkzr)�Vψsw!�g�|��l�T��x�i,m����ފY�Ly�v�ϭˬW[���a�����3�^��¦��e����ή�ɠ}a�8I)d���R\f�
�ӟMNa���W�����������,�-��ӎ���+)������w��^�8T�Y�����=��b��m-�]���a�e2&_~�@����[�yƴ��-�88Sc���Im�����>��ԒAed�+*WNa6�fc�CY!����2�3� ����cR��Iz�b i|��)��N�Gw�˷P?��ht�����p5��K��R�4{��{~����M��R"�$��S�鋟t�O&wy�o��"=�e�v���l&�Ok�iZ�Li�,�g曏��7�L\��q̟u&d���y�ݙ�1���K:^/iN�M�SP'!�o��n���`O���7�;�� ,�ΐ�X[ۮ�}}��d&x%q��[��F*ߤD�dҾ���c6�?��7��G熓�S:;��kvWR'��r5[z����>Od�dC��e�������%���ν��N(�73Ɣ7~���\d:!��
��t�����(�lf�pE$�m�s6����]$%;�$H�X��E�]&�Y$���D�s)�������Vw�_{�����?]�n	u�FmF��~Y����w��R
���$C��G�NJ�̒^3�����Y��.y�͓׍e��I .�I~���T�2 ��ul�p���<����*�y�N�2�\?g������+�w	x^����e�{'�?ٔ,+U���oʣjw����|�d���ŗ����H��aE:¦�N���h�$,� m��ƻ��(�s���&�]��IR���>�wGt��3I�;�3�a.�0��W���帢_��x��v�$��,�Uɯ������@��r�5d�N�����NvNaQ��g�F���ꌓ�Dm�h?)$i���-J�ü��(�y ʕ��(��cѸ��8�gL�Se��rƀ�LrC���bW�6f�pF����2�A���X���G���-�(�g�|�ȉn2j���MSn�'��I�03��Ƥ�
�/��E�ޘ�B�[�ס���3]cb��\���OӖe�cp�U$���l�;��T	j罃��4���Kq���J��� ��,% 2�*�|ٯ�n��Sdg��g3ҟ;q�X���v�Үl����}�4�(�O�⍊��?q#Ms�<Z��>���,�q�HuI��~n�������� �q�v�/S��K�0�L���?M����.ً�i��ϲt��2#��|uk�@���$���3��M��H)1`);9��I���ehR��uxi���豈'SɗW��g�P�5ũC$e<��]��v�����L|g���x�l�E1��������J &H)�d抙2��Y�g:]�s4��O�ͳ4dD]Yʢ���"�;�T�g��H�6F ��77!q�0�	�lHI}��~.ܖ�Ֆ��0s���ڗ�jǴ�)��Jv��b����N��K�-��P(w�I_���l�9�oǐ�r9��ً���^͇s7.��d��7�W�vu�'��*���̿#���1M.�3�l\�����V��/��\����!�&S�-Y�k+R*�|��L�"���r�X$�PcKF�ne��Ζ1����A�=nS��?%j�c���١
�$vX�,�B���La�ٗk�]d)ta�HO>�I�`���%i���>��.���S}�n�h����� ?z�}[J���$R-��\�t;�2[��j�9��zH��B�`D�+�n@*��T^Z�Tَu7H:��^��?�H��t-���<�{=�k#���/�D,�=�A�^�!i�����{�<��ʎ�b+ے.��Of����ZJ($&'�.�-�uɤ�^�W���/ǋ���Ϸ<��3�Y2�g{�-F��:������mw��}�BpV�|����F����I�+��>m`�L���jIT���
qa8��~��i�UL�` �U�������O�v�c�� ?�ϒ���{�Rԅe)t%�Ԅ��e����-&�/]������*��[/�30��nfr�(?."��Uz�Z�Պ"����2�VN�R8Y΄U�!L�W��A�N%;�tw�\�{6�ϓo�HDa�~-�a�o)�թ-'է���h�Ai<N�伊��v�g%c(/�q�{h�"�rI����ڑ��I�� �Q�Y��&eg%���?�A�ӰB�&̤���a��$Δx83��k*���!e~u_f�E�&��a	4�n7�"|���Rߦ]��	��N8-2�Eڲd���V�hJ���5=C�X0�����I�gi2!s?�kr���|��4��0v^@yAS�r�]���̢p׋(��j�R%��_�� �o�L���z	<Π��|�����(��f��Y����6&#?�?�-���~��ͱq͑�Н�0�H$Z:�s.O�?#���	ي�X��&���_F���1
f8��#3eb��]��Si�c�j|���^߇��r�<~r���ɡ��P�H�<b\c�_&�;��l|�
�>/�,>��텴u#.����R��b�K\&󗬞L咕�n9�zm�e�E~I���9��TN�)���O��Օ���!��f�գȵ�����]�1uĆ5�w�����;�s�K�[J��jIn��p�}Ύ%������K���Ֆ;\���`>q]S�Jt��($R�}�rW��ax��f��v/�3'�͙��l�З��>)��%%��q_��Jg��%�Xq�$��!�O&[^�����å��ңoXY�Y�()�SM��%����i�n�d���~�@8��e
�/��8�Qɮ�h�������^���s�+z�27���:.�r<vP��g �w���*��}3�
����^�����|��s�ĸ����%`|'�!�vx&���u�qRPϿ�8�W���k\�2[�G����x�p{�ʆ���dr���AWC��b�-�H;n�d|ӘAɿ�ִ{�LL�B!��d�Ty�ŀk<�s�Tb�(�?܉a6`N97�K�W]�d~��m/��-���|���^�i�}�S9>��ԟda^�� �,Cv��I�U9I���5x�bv'�:�U,U2��HB�Ks� �ۡC�|��Ӻ��� ���f���k:�3Q	i��C2�f��J!���N��Mc��&91G�VsP�����O�H��߭�&�ն8�msm�4�A��<y��^<���4�/DnZ'E���g���pa�3��ǩ����6>�DJ7T���նIX�u���I+�������ծ�q���r<Y�|2�;�X�A�W�o�lI�2��ᙖ^��6��l���}}SYc'��ץ��C>+�Sy���&gC)4�q����nu�5;c�c�g)vaӘ=��~٘I�W�Z|f�
|�Q��Kz~	�і<�|c��V$�S{C�E�8D��utde��24ѭ�v�4#۹�g�/;�ѹl_+}!�fR�)7z���Š©9��s�怔�v���绊����L	�[�����e�L�HY�P-�c*|�ۛmЏ1�j��9lg���@bZ�;�\��m5D���&[�����㑖FF �As����[G���+�.i��[� Œ�X�Pee��[��\�3c/tq2���K$:F��c6��R_�@�Ҵ�XI��K9�(/7��:��S,"��Rd�$�M�KcG��J:��:o�4΢j���P	������m+���X�$��2�0�^���S�Q��-�R�j֊�k&�Vޛ�^✚�76[B��1]��:�
ԫ��*;�MN��G����x=Z�W�L��^���#��8,�c����T�dN��X�m]�X�p8��j95�_G��մ����L*��|��f��+��0
٤��O�O�b@Q[��$�+�^�t&|���U@^��h4 ��C��� ����,M�С�M��ֆ-���:�g�	=f�~�ā�b����Fj_h@��N��+���l�Ӂ҈�g�NC��R�?�������ɫbTl�ǚ�1�Q$9�Ge��%��G_�zFi�.�Ѧ��.�_��FE�6�/#ꮐ[�.�=��ڿ)FG���J��V���6v����^��i}基˃�Rγ�����@	���*�<�M<ad�@����r]�����#��4�#�!ɷ���X�*�yz4�ȫmt�HN=��O�a;ī������A#�
̓X(���
a��UlŠ?���O��x�`9D�?=��ۖ�՛k���*b'����d�k�aF���zqu�@V�z��,��7�Bw��-Jò�{ǫ�Y��_�<���?�L���U���m��iLf�d�v�r�=�n���_��%���t�m�mC3\i����܁v߈��9_򘉝Ye×���S�|)w>�ϰ�❉����`g�4ɺ�fqE�\�1���ЈK�>Z%/F���z�M@����#�����I�e��N�y��oX�Z�� Fa��4�����:T����t���-������>�v1Rq�ʻ�������W��׾��Q�Ax(Y������'t��z�>
`���{������&<��0Ԥb;��C=��D�a��q*�G�;
c$����.B�W� �%�g���T�Ɇh���U"�^��w�4x��{O ��C{��*� �+L*��0�?�@�BK[Ax��A�)���(1|i���U�W?��@��tCЦh�)��]yD�ox��@,���2�$>U��������_y|��h��>J�H�4?�� �|V�r��zczzz��]�|��������0�	����!'�u	Y��ֻ�a����]v�fxZ����}���:Z�.���"=VLk�}o	a��Q%���u'+G�V�b�.�]y'5�E�5�������K��H��?��[�����(I��qgh����~��2v����۽J�t��c�����*ڟ\�R��'�#y=�	��nռItz2s?7�'#z�[2p!5.��Q�c�[cMJ]���K.w>@L��r��	t����%��N��e�>A	Q.ۋ}>E�8����46s�']*��
1@�D�8m�c�fRd�zɣK�S��P�Ng{iV�Ef��
,V�P�-p�$Z	�|��s2ݟ�>�b�/�C��JK{P(��u��z����	���
�e��Օ�v��;��>���?��]j�*�3(��ŋ�`���?�� ����X��#cD��S������eN6>�@����k�)4��R���;U��J5��P���2�6�<�T�Z @dޥ�k ��۽������Cg,�{��Ņ�
����'��P>��KK�&���9��� � F�h��
��t�������'V��3��������qU1�dő�qp	�K�$
�D0*�<ɔc�x��x�)��g&w�<GO��q/�	D*V����K�IV䙻����<:�{@��^�>)���Q��B� ���O7R%f���o$<#*��~�+���pB��op�yק��QN�V����t?�*P�Ϩ�R	h7R�	���j�]oT��N��t��U�j��YJ�����^�3777Ӝb�8�v;!�|XV�c4�:��<��I�G�SUڊwE,.乡d����Ĥ�˜��"����%��IwI T���W4�^ܲ���Oi7$��P"ӊ(w���h'j�gW�1�@���R~�WV{����ߖI��۔�dw�Ƃ㫯.�2SK!�($f����I�bligK�s�6p��.�	i�#Փ�	YTTvަ�hN���+2y��źd��Y�lT*5�y2�y�Э.�����X���Т���@rY+�R�k,ݻ����؜�Y�2������+��b�d��io�T�����_V��w;R��_���I�V���2��@¡^��jh����o�\�_�<�fS���������W�}�=?�7Ҭ���V4��t��C��f���n����D��X��^�J,�LT#�$�g4���0��U���y2$,�U&��$'��N�������C���R4�*��G0�h�ilcvv6�ӡ��]���㱉�=33M�v�@C�T�����1==�j�x� ��r�������~���v��92<$�<t*ځ��{��LOq������<,/�b�Cn4����r����p�}�^�:��K���{���A\�<F�,�W��q��;ĩ�괠d(�;���N��C� �ȪG�y=`�˗/C�P��Ç���Gg��L����7.���Gz�hv	�|��W>])��$B(e����t�n�E\�6Op��)ٜ���+H
ٷ��v��K�A��2�������SHE:v9�p't=$�����W�-ZYn(g$B!�BE%�'64��.K�8y#��uVa%6�7'�e���5$�6�vШ���E�w�l8W�
�����┾	���f`V�wߊ|���S�q�si%zA���&Jί#�%Bݩ��q��V�)Tr��4��/C�Ҳy��_H�%#�i�z�=�<ò��(�W�YC�N�9��̦��^.m6 uҲ���SS���t�eE��%,本�5yp�,�Jq!��Ho���!&�$�ѪTc�7����l���ޠ���9r'|�fs�[XXX�x	����R����ET,PF�0p�&�و����ǲ`4	���k�P�ŕO��"�ХY�)&U�0����F�"U�~Lǯ�ht���+W�������%@�N��W_�����T�S|���$��_�P	:A&����zS�RVOXl$���"4[�A��h*�'�O5�0��lPx���C.��ul� H N2�!�*��V��iP�3�������/��K��Jŵj�iJ���l�
6<5�m@����uz|L�'�V���[�����=�a���ٞfj��j�^�t`
�^�.�Y( ��	��677{�i�<>)���<}nyq�A�'�z����8a�=�0��/�+� EU���qv���y4 �#��Ֆ��k��@+ 3����={�D��� <��|됆T&�.@m���#qI��ba��F.uTk�0����Y�{a�kvLy,�����a���EX��%+ܘD摜K��)��//,|��a�N�Y�s���<:� P�dOC��Ǿ�W�B�1$��q�&Lf��`��%$��uL�>/�¯�Iu��mp$�=O�-����E�����>�dW��>Õ
)�����J����%���<e�N�-7pu��C�>��}�wT�f�]M֢@9z)K9�euH���V���b�.����)�xm��-=�>�Q�g{�/��A���� [�p{ H@d2��<�*t�	��I;J�$�4�R� ���}؄��Yb_���V���Q��W�{ƥ�QP��¿ �k��	�� ,�Ξ=�%@���@*_�t	�¹s��ͱ��~�&��O��"�	A&q��܊��WxFk��4�ׇ\DXl�O������K�O�I.^��P/��VTt���X V"C:��A� �¡R��W��7;٠f������mc����0� 8��f��'n��TG;�{�.��'�/�S@���L��e���X�1J�.�I�.V�ؽ{�ÿ��_��]	�!v��qf ��Ӭ��ei'@���M$w�k'��OP,���n�]Ȑ��*�p����XO�J,�L`�K�uY ��ν�Io�Vun�հ?�M=�9UoX�HE�w��6<,�	����"Tal+5>�靪��w����?m��(KD�N�O=ۇŖٱe	j�s4:v񁯕�*#���:�w��E�[�Ͳb6�R|�*"��uuL8�qhBp�Y��\=�i���W��g�xM��0���{�A�^��yM�r���9���
f�U���*"g�6�g�7�	;_���[LF�o#��m�������;�vJ�	T�E��_��gl.]�H�����e�I�G�_���J��\1{�3�*j���Z`�M/C4\�%6�^��kS�q�V�E�w'Y��?�%���jf�ԍtuJ\�Ѻ����qǅ�p�f�`�?9L����#G�8�7*tXE��d����g x=ؖm>	�(�{^(x�������������1�5JC:-"�g�T����<��]!�� ����hn�GQ 5���D������J�HAN(��G���G�A��ڮp���7z`@��*B����5�b�m���W5
���ᛨV�L9�D0;���<��J\��&�Tc`8h���P >�
x�sf�	�^�%�M&`���l0���XV��<���1.�B�}E]�|�4�M����b '�d� �20�a�$���A��\�N���x�qլ����X�F��6���I�_+��U�(ǩh�C�M�s�����g%�$�7:��aO�,<��}:(�.�ٻ�
������	dܬ�e�ؔ[o`�p?�����'�4IF�����0D����r�ZH��dv��8�	L�&_����A"�V*������	v�@��=?;;=??ߘ��]��� �j����ju�	��4�IKik�GWD��+��CD(��������3���\��4�f��{r��U'��̿��N.����%%W�����x96�xz�ӓ|��T�C�,�Y��L�	���H	!���� �1��g�\c5�l x���C��H�zr��_���W�5y�W�#�O�������]7�ZZPzOO��9�!ɝ��o���'�r��\(�ƚ�s̏l�|~OV\j� 0�����cKmm,e<&e��1V�!�16���7�Zls��D�Qf%D����v(��2C4��n�����X���M���x��
��r�޽{���g���� ��V�%s�X�i��k$d�
u(��� �3A�������b�/��H#�Or5:�:�mL9���o"be	�륗^b- �o�� �{�9:M�ٖ ���\�T�Z �
�+�j�K�F���74�l��϶L&J�S�*��{�[�?�z�&I��L�w�%#����A")6M�L���ed�ѫ~�<��iL&3Imj��$R ��BU֖�k���|�|���*p&V���p�˹�|g�xB[�8.�U.���d�@q�x�0S@�\w٩@��0��/�#��O��1�����.��ԍ�����Ȑ>��I�#�Cbq�Vl�B��]��w����[L���TٵxH�yt�k~%�]���T$Zrq�2Hț�p�R+�Ч�㡛���<P��_�MR���%�I�c^-f��d=�B���)��[:u=�����T� ��k�\��`�� *�q[I���-��v6�[��C�y������V����P,�b=�=&	˽ʺ�,~k���ʞ\sVI��/i��e�����F+�5�'_|4jZg����p��-�w�\�\��<{����poo���s��ʜ�㝫����Cq���-�*���S� M58C�e�J�&PS�I�l�����O��ˣ&��}�Oc�L�/��/��d0iVv��۴zb� �Z�Id��|[�&������̼�\������J0x1z��"v�>��ԓ3JuU�Ye�U��06V݈5g�(�睑�gU+A���\K����a�5�1֙a��V����ɘ����6��)�B�x���^��.�fd�I�B	�����P�/^���=܇=���e�U�LUe��}[{M���?�.�s-������j�*�V��=���2P��1z:	�Ao�J���JN-]	�j�8h����q��z7������ײ��^r����؎�$�I��b�Y�,2uh�Sf*|�\j��<�J��뙳�[oW��L� lw-�z�&�Fr��]�1���
{�ȡ}&��*��>� ���_!�V\X�@?�&.�t~�;o6M�夗���hB �����\1�o���;�(3m��]����G�jH
$:<>����� o���%�ޓ��"xn�����Elw�ܑ
�܄�u�zIJAş���=1�����P�q���܊y�����?����9$����j\>����8G`2"�+1]]�ಃ�\�E���6�rR��W���'h���k\C���o0n��QC�Z��af�#�
�wn듐�z1�H��S5�\�'�8�ڟ\��I�@Tuv~�a2��x�p����p���	����b.d&%�����
�v�6E�)V*��|�p/TMP��r!f�(� �I$R�C~'�k��X��֚%~��7@LYϸ��l<�3Af|�P�W�ـ8	r<�H��0�G�y�GXաJ��h��.E�A>v����͚��@��rA lG8�-ZA��;D~�����]N��zِ�_�N�ؗkRHM��uP�'�	n�(N�Ȕմ���<��3����	M��H�rA��s;:
�m���3��0��j|4�)��K�Hp�(-HA��b	h��	sxI�7G�\Q�Lm�&vB��n"D �LGl�6���#y.�#)�5�<{�,�S"\5���R}�S�+V	��| x�&��54���ԧ��g�Տ�����)��b?�����T�ps��-���)�q� ����...� >���իWT�pq��g��
�&�"t
����֧����'m�P��?k��İ�������.�A���ժu�Tw�l��o#�x�]�XG�3?::�L�L��z���9�#!��W�
���%9s�0�z��5~�����
�d�]~�������60e�)	Y��-��ǆ�$�[��&�r���*�@��_�ml��jJѪ���ݻx4�K�8�Ǖ�����1���&ID�k�JLN�aD�K�r�F5��S���,�b�E)*m��U]	��Çi�`d!�]ub��A��'Z
�Q��-f��J�q9�[�򍭸H=R��sG)B&�>#D#� ���)8�Hܐ�DTP��o���*�Vm�;C�Px"�%+��%��$�N�7t�h&O���~�yVU�>'M#<���$�]o����	_V
���5N��k�l�ZE�ԑ���ؼ�8�I-u�O+x1�h�ܸ�'
`�sj?����wied�\^�Y�Rlf��K�V�ǸE��A���3rF�,�Q�����+�DmL�Og��NHj��mks�ZC��� uB��@��ci+��E��YOc�p�o�#2�g��֦
m���	�N#D<k#�¦�fD}��zT)t�D2�V�؂�^;�e2(}ÎD�S�����+��،NH�֘ #s$�ZoA%�f�:<��Y ��}�~�������\�����xaD	�)�=&���O������6��Ƽm#�7C���>�A>P]�p�e�1�3Ҫg�a�7�9�:�x�$��S˺Q����9���!�hiK-�GA#R�!�ẍ���,ګ@a��P;�N:��A��o�ɉ�=SG��v�6Rn�t��>@���)��mLTK^A ��PG�vC�l4]pV��`X�Nj��4e[��y��θ~��d*ؕEx������=����1�v����H#eaj_��6�S�G/h�k�$/��j��e<KU!����E��P��Q����MAU�;c1ѫV�P��ꫯ�����`8�,˫�Tp���?�L�{��������7��` WW�t��ѭ~6�����ZMS����.Ը$$�6�uA�[JϪ�N�q ٷ���_r1��d�W��͠�5���.9�*�X�Q8J�A��ϛ�"��,q�W����6\��sE��Z	OU3�fqcۘӧ�F�.I
�
�޽x"��8})8ʹS�O��Zm^�|-8) �p`�1#�����z�+\���AߚM��{��l��� �?�췳�c��ة��L�������r�!��9_/__4^���,���I���I��s���_�A^e �bS���k�4W׻-d+����*4�-���˩�Wn-.T�ƣ��΢Ѣ�O�<�$&�=�6V�t�LAj�5�M��j�b���KR�%��6��#S�2���zN�R����
'�*?B#���[��r���^��&!u���\N�ؗ��{O㙀�Sjv:��<^hl�4g������ʮg�͜�����(A S�1$�5�y��O����J�͉u��˷���F�7��+��遑-n@��4t8�!xVZp�>Q��d�X�m����5e�& s���b�׸���>�!b,�qSY��BԀ��E���X��r����O��F��^Va�G�z
o6��1�x�8M�%��a�Ư��Ñ��ʪ�����M��/�GFR(��Y����9P_�����mP�&�g�����&L�*W8���{�P�b]J����㓻�%��:����$�a��V�$2�5�1u��é�ݴ'�Rm���4����
�Ȏ�������հ��'%0AԜ}���}��P�z�o'��Z)��	�j�>5C�5�بDre+�FHoo8Nf���u��T8L�&�z&סQk:n��Rj�d�[����-mm�g�hqb�YF�*�-^5R����8���`gSuC哛{QUVŦ�l5�^U��<����O?L�w�.3-�����o�ɔ��A^�ԕ����qA)F�O����ƉҪ�)Hxz���� wRj�"H�8���*�U��Z�uQ��Ǩ�&-D����0*�uo95L�ٶw9���5��g����V�%��9B����q����\I�*9��g�z��L&�"�u������B
L/�|r�}��il�BF?��'%�8;;�6I�B���?����?��4��_���G#,Г'O�ɨ?�l�l,.D)���̀E0;��0�p9��ή)˩�!�gf/���c�:�Q}́jl��o���IҖ�t�d�l%D��O܀����o�P=� ݾ}��<�!|��KmXM�+�8L��޶n
����X���@��{�~���ӧ�'�ނԡ=����p��b����)L��Lm�{�ܜV���o��Ϳ☞N�К��I�nL�i
�i��g?D�'�^�j�eb�Z��  zO���ĶeA@��6Í�k�>�q�U�g��}|�2f��>�F\�e|����Ǐ�E����*v�F�^8;j@5&
�Q��.OTaGE������*	��N�0h����=[��ђ$B�Q��:�^����^LV����q$��:�m+S?�wv����b��l�t���jNӎ����塞xv���j�Ԇ-��j�2��R��O�pӚB�a8F�� :��l	x���Q��m�+��e�@�4�Q�v܀��	ݤ<���2�7Ӫ����cx�  ��IDAT.<r��m},0,�5�s�Ne�� #���vp���:��&�ԉ�*�#ގ�d=���h0�D����j<1ϻ����0��m�c@��-���
@�B�C{F��E�Ԟ=[,�'�B^���ْ��s�#"i6�~A~�2y�	?7.T��(nm���G��&�0d�,�=�c"�6�Һ�[����[c�Vv7�銶4����c��X�����L���o%ݶ�ϴ��!r�η55B�ǌH�J;��b%��8������3c�a4���)��Kh�=��+2ً�Soh���$�YWR���8��nNB}��x��%.���D�Y�H��I$�<��k �)�d(Ҫݔ�Njj�Q�÷R����o'���s;���� EZnͭ��t�j��A+M`��{��f��y����(�8��=�dc�F\
!���� ���\P���Bh]�%
���\��^�9q�\C.�p���.��K�dc�Y�tQ^-/0k�g��l�����W_ab���̄�@�5D�Xr=%l0�ٔק�X��w��D@rAO���Q����,�/ 9��m~�ͷf�&����g/Z�E����?�-ѵ-���7����	"�	�A�Vb�� �4�|�jc�I������T��k���Z�{V�raI1����@�l�7��K7ea�%�
��9�AH�X�_K-4�7��� �ul����9�'J��1��|��g4�z��d<&�G��}�~��l1u�GO��xyyYkE� #+�E_'e���z�>�J�``�$�����5su�g���aq%��x�s��C<�F�PYF�� :���BL��|�J�#%�"~��ט�v�I +���\�2���ΆD����}ZM�Nv�e���6��Xg)��~��� &N�d#l��4��4[QS=>q���ґ�D�����r�l�>Z/튇�2>z��І͒�k��`�sฏ U�7%���8�uQ
�`������4j$&)�ّ1�t�b �-�������Ql��ߔ����	�gy��ɉ%�*�I�g{�3+�:i�(��W�+���Y����{|��������7��vj�8l�֋m�U�W���q�H�6}~�P�	�1�lb�/�R�V�h�^֨b��A���ф�%^L4�WHZ��ad��j�4qi�bHb��ִ��I|�����Kg�����Z.�t�[�!@�cd�3�[��8�Y�4h��D����$7EB�W���݉OANUa�^���I�{'�����\.M_�з��mcR UC2~UQ����)���I�]�m3G�ȩ�*�q.5�����ֲ�8,�$�����*c��'�[���`�߆U�X)^TWI-��,!km��Q����dF#K�l*}�T����5���Y�,��Fq�c����i�Q�F)h�(��|=%�҄dI`a;Q�e�W�X��ܿ״!�Zc��<,�����c��H�A>�g@���05������ DF��`���Tb8%���8Ǒ-n,�*��J�_�\=����/�&��E=m|o8����jG��B[��>EG{ܖ�i�4iL�"�a�\�"Y��rzzJ�,�#���5K��$�#H���s��N��6u�5eg<~������֭[���	\�fEi��zJ5�D#i�L�8\iAW�E*�&dJ���]Լ�U�c01l����+���_�4
�K$�P�w �.r$�D�&�2�ۨ29��&��Z��D�8?��l�e��i�Z��gP�u	m� P)EHh3��'��ħ�A~m`�!9c^�z�#���&��޽{���������.x���_��T�	�U^3���6����wtt���������� ���o�Ť�b� ��bu�S�PK�f�Ȉ�h-`�2ՑR9x�20@آF�	�#Dk
���K�A��)���8ފ#��M�i�s����M���j�<³��Z���7��BKC���TV�����,j�xV�=IT��I��i�y�@Ȓ$��FU��8�],�ˬit&�U8�����vS<�L��V��N�mGyC<~ഋ�|�9��y����:����.�0xι9,�);'����A'�H�����ԌT;�"}���}��~�~���8{�38��۔#�����~9?�s�򂪬iY!�o;���;��~'��,`�nzw:����s�����"e���I$]��\p��7������e]8[�˴�l>1nC����8k�G��;�ӳqu�$젛~wo_ݲ}�����;�p�\C��J1�3EB'8��[G-�l"���LRΈh�x�U;J�hfF�5;	#�<�EI���߱��C�m�Y`�$x�a�C��6��8��Ɍٙ��o��jy��v�������Bp0��<�RG!E��an��k}�|������V�0�M�F�ق�adV���x�jM���'�Z��5�4&���|	y��0����d)��i�3f�Ν;�!~u||�+��Çi�"K>Ç��J��)yC�����'� ��{�=��	,ف�Cb��A?\g1���m�Y���OԚ3�ׅKA;wS��-���]s�S��̆�^��G����'%�Z�4����O���R%�h<�`n�_�����٪S��&Bv�g��޾������x�dص!92���/����E�
Z��&*����⺞M����^?#/K��MU�.�p���!������?��'G�t��ϟ��J`8��#��C0�|q΍ƬkJG�бW89�E	�M6n��liuJ$ko�bh-��m�qf�c�<�#LN���9��F�=|��0�n4�ۭ����o�@m��6g����.���^ڶKz�(?R��Q�����(J��7̸������?�`c���dǅD�)/�����_^�Y^HT�P�\j�Rah�j�����ͺ��,��� kow�W-?�+	Z_�Y�ׄ�9�u��8�o��q�0�A/�'{��X[H#Mj�#A�=u���˂�C�Z��9�e�>t&�LT�G[�ܖ;hD��|����i������,$͏�3RV�11
S�$�c�7
�Hl�?�����dce�4����2�8O;-�4���3�~=(�8�i�{��!i�G�VF4P�)ե��\&���]?��2(b��}2� Ob&��O��fC�Z�j��w[��Ë��낄�+0�ڜ<[9(�G�֡v�s�Ss���9��y�	�׻��b���dc�`��^v��A��q�3�#���q��:����,Mc�6�H;I����6SC�ٮU!���ˊe`����V_���%=��n�r��x	�5ىw�αƤ���K��dF��=��&�������D�zy>\,V_|��o?��|�$Fd���TW�?������lVk����2�C������bmj"���?#)��!�]M��h������vyj�`�oK�:}G�Z0��ti�X�`]4E�:a�����MhWJ[3��H{
խ�=���G
��.����)�k�e�|0�У�r�٣��)C5��c�${���'u����U�B!�-�ۗ�a���r������ƴ҄�S`���EC
�@�T��k�'9��@ު��Di�*��v���1;�,H4KdZY��������4/R��X�r��ݫl�8�@?g�f.B��9`�z0��&�p�6����.�ˣ�b��-�̊n����g���?�x^_���X`�M$ތ�TiR�Y�``q���a?��u:�d�%ǯb�)�q���E�я�`���Y��I_���Wt>`�LO5jR�C��t3�t_��=��K�j���J�.�XG�o�z��?*��x�C)�B�
�Y�y�s�Od���@O��IH o(�3>�L�S��،�fPbc-�j��w�Ƥm�b_�
�z`���T�7ņ.�ڤ�G�m��И�%5Q#4Jɨ��')i˔�FW7�X}$�C�$C$��J���
/��1~nU��v������G; J�c�K�4b�W�B��'rj<�Mm���8K�&��K�
O⌵jN�ONNN$�k#���	z���N�sEc��b����q��J
	���IY.�}�fL�¼�~����@��JA8�jmZ�lʇ�a�c�?��c��dʮ�A`�0���L��4P�"�ꔭ��Ì���d^�05��l�O��4n�SWT�ߞu��Z
{�i��<+1�K2e�\w���୿̷��
�m�KQh�:H�1o��ئv�t�E]�2����m-��F��'
�2�p,������cs�����ߚ���T�R5�K�倯���V4��~"�d眼��zv�;�[��m��u?&,	mn5ק1����`J����8�h9�
��-�wlc�m��q����n��^6o�Ϣ��$JHT[��ױrѡ��)�fQ;-�re�-��&ݲ�l8��l��?��o��R�Dc[�X�`�8���D�P(`�j���s��i�� ���sM1�H��r�p�&5G��JF���~G���O$õ�¿�����������ĵҚr�����I�����g��'!��}\5/��,`�]-Q�.��J���ۉ5b��$��BV���4z�<���Pu)6���f�9��{��p�N�߿�'p�ã��,��Ðe0s)J�A]"ה��JɈ-{��ɟ�����C�yj"�5d ���+	��W�Qm^�zq#&�邂	#�����2�q�,ݯE�4�-�ڟ����n��nb@�������LV�����Ç�~8�I�P`�9��x��|2�HK ��N���~������ޣG�>?��������?�����sĿ���^�R�Q����� 3�Tᐾ�g�u6�Pi�S��?]�cL���������_{����#��ߝ�x4e0�'��̶���Fv2A����'�=/{���PlTaϦ�<�Q��#����`瘘��X.+q���M��� �6L��{�7�M�9M�L1=��F���M�cx���`or$�y$�[������C�9qC�l���
HD���P����%�^c����Ò,u������S�~�?��QN��z�PN��C���Ht/���3,�Y���t�2,;����Y�+N���Q�S��f����b"�d��=�%�.w��H�G����~��AZES��^_-���In�(�(��{�/+�Iݞ�ڀ�D@�PT�E�c��A�EE�O.'�KR�_�������#�oww��2������z�r&����H��l~CSJ��g��A��e*�0F�]��p�FI>09����tTӲ�x
7o�	됺S�2,�+2P,�>�|��3be�F:uŁ)b2�(/���D<g� �^�ǄR�`wr�o��z��	sA��L�%�h��5�FBg�;£�F�Kݔ;�	��j��s���s��k�5��*E'�uO��g���}
��|:����m%�`k�SV�+�3�!j����,>����
堃Za�p�j) ��!����aJ��Z���X���z�k���S�>�<n�Ɖ2�[2�զ��:�OI״�u�e�ʍXn4�{A�i�Mi.��6�HU>Im�����C9*�a3�	Ŕ%�6[�,�!!�7d�H�:&�I�u����ԜVl(��j���ên,�$i&y IODl(M�&ioy3����� ��gOE#d��gՔ���/�TG#������0M�5���D���<��5ǋÚ�.��*����N��ŋ�a2�m{#�I8P��fU�t.���//�).��}��ɯ��?���o�������C��Ʃ�D��Ov��Aq��޾��ڲ�5�e��H$k_^H`C��D�lk�G����g��|��H@�$�AW�W���;*v�G?������zu��]�=�?�8�2�~��h�M�2ʊ��>����-�&��m��#1~<w�Y��/ܺu4�k�z�3�D4�}J�@0�s�ɲ���o=�_����T��WP?��K��q�K���y�\qI@I˅I�ѪXƜ�6NSmLQU|A6_}�������ʲR������h!�)�R�������HG�����x�����Q[}�3�%X����iLx�bQ��#�?�y�V�e������(�
Q�����U��
x!(��W7^> �V��(C��/� ]�
��r���������w���t	����6-� �kzW�yA�uym/
i�`=B������{~kZNK}�4J�0�
�G+:��Y���x����n�=8=�����Q�B�z�YT��MZ����uW��M��#�X���	P�{E&f©�#}aJ80T}NNN�C�O��E�n��2�X�7S�W<7�����,��%�)������iJ֪H#�����ӗ�M:�:r��jQ��{.0Ǉ6B��2��r\k��/`��[�c��������0�,���[���J.��kY�5�Mc�L�"�"�I|@Q�y�F�&O����X���3�$�R�T.U��
@z*�f*ֹ�?�v>����u����iqt<�"H��J�\�S�H5���u�t����m�b������!-1��<������2b��1�)pK��<�Tm[SaUz�*{e�+cD�r3�F��H���Fxl�l�9��V�x�]^^R-�9�f�P�s��edbI���<���?c�B�GLK�AhRR��9��&6%K�,�ҵ��Qp�5�e�o߮�z�L|�g�AZ���G0�����&B
<�6���5�B�dc��jj�ߑ�*�����񉨓�����[&�66s�T��2��1�2Eu�(��L�*Q9�;�#�	��}tO��]m&)����he��|�q��1��J�^�Q}Ҕ��)��(�4mA�3#����h��1��t�}���"��N���$�JkJ�˂�\ҧ"���<k\1��=�@�l����9X�'���Gˑ�=Zq�[px]��⋧O�➒�?�;x������|�����n���^¨�7�_����g�������o��>z�H��������D�}��������@� �i��n�G��4�>��8�� SK& ��?��ω�U�2��T;i�S�,�b�@Q�y�lƲ����vo[��>d�cBs#!a�Q���$~��n����q�.3�L)��ɓ'���\���EU�b�p�.&%�	X6հ�����ڐ�V%5Nw�8���=.��o����&ԇV�:|�d����29���&��?���?��?1���6N�׵U�&�Nl� o��Y�^c�;#3�v��.��Z mU�|q���;y.*�����pd���H�Fr�q���ȡ��z)��xwBm�O�-��D�m�s�"Z6�F��T�e���p�������p�Jݔ��q*�A���`4���WI�w�&�D�!&I��.�wp"V��+�F�|�P|�2�0ф�!9����A/��b�`��κ)7��~��1P�s����#
Y~]�j�>���A�fS�RS-��RU�E"�}���m��r��X�^�~������o�Z��>6�G�oEx�<Wi�4Á���.*L`�X�f�H�A��iK�\?JzI6��ӬH@��w$9���a���_HO��TuS[KVnC4B�0���l�'��)ܖpY;���b��v���RU�pG������VY�h&���c�-�%�/��RPr`�8]����Ձ+Uyq1����T�q�a>��%�hgD�������E#3Rb�>�D��"X����|5��+���i���hE}x,E*����f}]���A>&F��im��ğ&��>+S��������7u��j��i�v,_k��
�~?������K��p,�l29���Xk
bJ���|l�Wh�E��©��k�Z����b��4e��jF��,��R<�I�ƶ)M��	G�P�4[�QQ4��i��#�q������Wg����8��6�."�b��mZLqڎ�&�S����/�]�y�f�'/��"� ��!"jU4��F4��)�'�`�\1��9�;X�����҉YS[�@p��'�RS�	��Ǐ>���)i����i�u%p��w�`1�ÛN9�pz���=��g
6)����N�Ӝiy#����<�7?��Oل 7Oz)u�[PذVx.�\C(:��㉃~�@��&����b���>�A�������Ջi���X����M���K�m�	P���f>��,V�X�� A.����BAɚ=u�Rs�Ě�;`1�A)Cq� q��و��kZfy�x�Q�n�atq�%��p�Z½�,|[.���5<��MM��v�w�
�zx�:yL���;�v<+IxC���hжCK�-���̊/j\ξ���u�,Hl�d�N����=T6�ȷy��x���Q;�U��~zN4m�����n~��_��DM
G6PD?��Ǟ)�]6�>u�����*��U�T�>s�N�X%��p p<�s���Lt�|w�-Q���l}S͈
���*�5�Tߴ�M��R�{�	\T�Ec$��ټ��+wc����C�Rg	������4���b�u�D�kD3  Uߐ�g��ȶ���ʳ�ͣ9����?a�M��N�qk�����B0a%��II�*�E������5O��Ȱ��P<���h�.)TD�ЈNrJ	�_,
�u0E���ΙH�����֩���]c5WD��e$J�o��QYڃ�J��#ÌG�C`��UP�� ���Y=�*^ GSiڼhrt��q���X̈F/F�ЖFHTK!��;��U���j�a�d��Ms���Fk>��ׇ�J9má��f�T����ۀ ���Ɔ$��� ~b�5f�S���sH�e�\�D�h��O�MwF`�p��:�Tٞ$�-|Es��Y��bZq�m*�VJծ�	�VB&�	�/pq��q3�i����
ak���]2H�����g��5-g�2b%JR9��R� �+,��6����9:*mm�xZP�}Β͹C7��>V��`������s��c<x�d��f�]���eW�<�)��|��V����c"����~j�����w<w 0+�ȉ�����cR;�кƊz�M�d�>� �3���⼲��} z�j��F���a�	�jVfg�#�����۾����O��8#�����Z�W5��" @�Dj������P(�ցE��}nlB�)����2�8-<K�\��ŨS��b/�ū][I���	%��v
��V��#?��d�hH@/���$�5�0S.�'�|�=J��f3
�?ȓHYνv6'w*�~�Z��a�\gb�Ɔ��6��dY��V�wL�ƿK}%��	�܀w%����l̬`<6v��8�M`k��.rPF��eJfDUm��PJn!��O�*�jgo��P)�U,�fA��%�=#�1��sS��60ԙ���ۂ6��[:ޭ9n`C#�j;�b)�*��ɇv�`Ӽ���k�k)�m��j)�?	��?�9����kφ�����뉓3��B6���,��Av��8���v��g\�V�	�Rm(^YhV�w����98� �����L�R�V�mU��U��S65iv�ã���j�<h�팓aD�w/�ډȋ��$Ql<)����$�1�D��S_E���b�m�6^SV�'��,��)�0p�~?�:с���XE_o@U�$�^�0��gr�b��>����g�q�˒TRӆ���%���Pj�J{)x���~��N:�Q�"N�~.#��H��z�Ժ]i�4�w���(�I��V�H���L%�IRՀ�[��qo���t�Rò�&ѢSˍ��Drm\]3*�Y����MQ�al�<��p����c����z�WeM@��c���&�i�?m�B�)��KE���bA��Q�_����s(����5�A�1����b������zIJ�(vu��׆g�/��\���>+ڟ��j/�T���ͯK�N~xx���[�@&�B���נ������m׹W�^y��1��Ʒ�~�� ~����"qr]\���%�ș�/Y��f�2U-��_������Pj4�HLFd�W�U?x�������g�(�l֞��B�����{%~����
�&�簌��t�2C��keM�Hߴ�aU�-F����^_<=}�ryP�i��GΨR��W�1���{Xտ���"�������}���������_���I�Cw���*�~�b`�S�J��T7�1�Ǧ�]�gϞᆐ1�!�7;��cX����G�ѻ����|��_����Օ���ex���㎛�:U��֪4jV�0*)���+�8�Z�'bN�;��nvEVN/�TMi�i]����	�㞶 Ʊ��nR=?T�]y�C�χмo�s�8��r�Mh��Ŧb�����e�jfY��e����0
0�R��Eշ�Ș�C�N��H�MV���,-�dT6/���h�3���Sq��q��wh���2��ҹ�vD|%A�E"z`��=Sǘd��N�%:k����塍�ҁM��qbs��ܸ�&�0fs^��U\��%���!�b��L���	����i��9��a�����C'�Mil��ݦ�Pu�e��Q����9S��Zji�U�]��~���Lq�ʍ�Ţt�Lh�^������&�	9��c�|s�����_����8@`�H:�6�:׉y<��_f�|ww2٫���d(�qo��dRx	���Tc�Δ'<Z��Y	������WA�dn��<wcQPp7��t���X��cxE�.6�$�� !�� c�F�X�D�#Ɲ�=�s9`h�q�����y6�{�J�y�%^U_�����,&�Ʊ��!2�����4{�L��m����*�J�dD����P�ݜ�����n��E�A����G��mEr�V%�r�A�+�ST3�t}�0 "k�bΎ^؎:�N���F��ȕ�\J����ӑ:�y�`�d`�I������P��ٕ[�5$k���I1����S�0�6W����4ΫT,�\���Cf�*s�,��_�'b)���h�._�X�� ���M [$�G�	�g��;<�y÷�,���}�,�Ls<;;��G{a� ;mu����o&��JNN�����޹s��o�󢖢�0b��w����
0�
��hg���pg��q�<şL8���1,����ŝ�;��?��1�/^�~�>j$l
��NҸ�������E��g��<��E�!E`�3}5I�O��Џ��|���;��}qq�6_?�я�§��ϞIy��PJ��!a �W�|a2/<���b%��������������_���¾�����Z%�a���L�����%ޔ�`���W�[��_<nT����8��y1�V�xj�Q�)n���\�|}Pjb1Ւa]-��+D�*t�$fJkr��D��)����j��B#��S�3�
K�ޯd���S����#�����y�2��T��w
�!�ਠCje���h<.5���÷��m�唴��|����1���\�Z��.��e�JZ�%��z6���K���
��)���P�m`"_S[b��I-�t�����{���3Ɍ�9<m|[��v)�Z�=WE�7�D����,��8E>�)M<��z�.E6�#bu��4�qh�-�������:�BSnsuNjm�5� #u���i�X5�p�Ŧ�-}��A������e�ackWy��K��uz�����;F�j;&��t��΅�nnՁ����w�O�V�L�Z$�_]O���Opo|)�	/�M�m��w�U�O����=;c壝\�t�"��^ $&���vS�Q/+������7R�Lz$G�l������w�>��i�Jak���n�>4i&q>m�Áv:%K��h����n<����	א���Dգ*^�����f����u8ޓ /��?>8�����i�Z��4�ƅd��1�â�w���k�X�� VJ�����jFD%{<�$Zv�.��i?O���1՛�\"-JA��[��ARf�/J6#P��F���ō"�Oa�lF x:�{Jq�8f2+YH@FU�M	A|F��~�,�i��Vk̲�<�Pz�(Zh�o�4�2���������>�9���_`:X\��V����}�s�b!��GR+�"8�W`�X҇�c����O?���G*��3� �S=saH[��e�Rk�.��y ������K��RJ %�yrr��}��[�Z�$�w�%;x�����I�`�M�C�/�*� �;.{���mo%�P7|sv���b4�
�"Q�SYi���g�}�o>|Xj�3�9����`�'�O��:��W����g�'x
v
�LP2�Ԧ�q��l��v��@�O�H&�Op��;&(�l��Gq� )Qj�\_Ij��$��������G^Tj��_Lt���@��/����5���g��ႃ���m��Am����;I,�c�����P=�k� ^oϵ����f��	�Bh8�\�fe���
���P冒b��^I#�(Zo����+5}�v��k	�;������+,+"���A�yUJ3y	"i���+#}�]>�4�^I��$]0�Q\jH�����u�l'�lUu���"~ ɭ�z(��q"�I+�*����7WW7���h�Cjצ�rfSI����V�s�����р�1�!�C�Xk�`"�Xy!)-�cM'[�[�2g�=���j��2X��52���������Yy_ʞI{.��(?��o(q����T3Bj��h��1eA?��U	�T#K��2���$��lNU�^�gǕg�DHy�k����^7����pZ4�3�*��Fs�6����1�E5`g�9�A%��C�>��[��a���jmOB��Na�Ɩ�PìL�v7t�0r��!U�H'�	m���+yˌ�}���s�M�!C��<�,��e��U�?x4N�Q��4�s�+%	bw��MY�o�s��PQ�)2��{�����7o��������}o������>&ƺc�ϿC��5�
Э��M�$�Ș-��y��`��r7� ���LM���������'�$��fGGG�pH������|���p� l��_�k҇�*���.Xm��(�L��X�C~��?��������=4��R����.B������Pc]�_��/A��Ӏ���'��X����Q ]\��^`�Z�*��Įݺu���/�q<��#� �IO�6�&���oX��{ϟ?��{����� w��<��u����g?�s#���E�r>�1_	+�fCp}`#�]���U����`��b^�4���ة�A`0��� h��cc���/����?�����Q	���0�qd�橥�#�*[U�S9��w��D�\bz�P�%J���D�x���30��K�.�x�V<���җd�~[{�`-L�M_s�q�8��m���Ns�rj���]j���� �V˗X�#,K�|�y�#-�	Ӧ�AEH��Iu������҈�&��Ⴁ�*${�|�s�����{��B ���?�ܡ�;�b:'u��&��� s{į>~��T���ёgY�S�.Y��\�� ���hTJ��=�Lp�.h�`�${6��:��49c�����T����;�������>���A>a^-N/� �+ԯGw�:�${�/�b��ϟ��I���t� ��~��������#��h7����)�/z�ϠX<��V�M#>xc�?�����Ő��)���bSyJe�>��v礡�dF��>^��jq��k��(�aS4z��)��fy
%Ƿ�9�	4�P�3��|0��e��.>�ݸ ���ha���}�K�fJ13����<5�@0Sc�_�xT�#-I�G')5�֖������7�&�B�K�/��t-%\=&aĶi
Mt��1�+���C[s����b���b�[�����\���H5�y�uӖw�0}�סM��$Q�xMa�L�a0HF2�Mx6[���TF�����[�Eq���K�j�˃ct[������W蠒�&�]����aWWל����剁VH����VL��L�k�k�i5z߱��Wc˅tq�����:�;qG��:�5 :0ؗ�a$!����a#Cz�)h�|����.�c$�`��df83���M��&Qi���R,��_��S>�/�����K��}��;w�ˀ�tx(��$I�������c�(��Xz��9
?2�A=&�)���}����Hb#z�|��.�Z\Y"���kS���R��.M3o-<[�zd[���2��q�?�� �������E@I�f$\��p>f@SLd�Xk�ly����0�q�'������ik̪���2+��=~��D����ZF�@�����fq��Ã�]����k�� �#�Di�W�-p��['7W�����\�[ϯ>~�	-v Zi�?툗9�o�1� �����/o��>�(���t��f-�%��`g"V���n�����]q��H��7���[V���p8x���FG��e�⛗b�������޻�^���6�zs)A�i4��<{sr"iM�T�ڊC�������z�|�ȼ��o�w���a
�����t~~�iahzF�L�Ŧz����dGR�n����ymJq�a�O>��3,��Sb}��ݻ���I����7��}sq����Wg��?���5h{>?;�P)~8�����W�x�h,�xY+R����h�pz���g�/vv&�U�X���u+;X��BrG4νd�Rx�HnjMxd7����Աڝ����sZ�$�3��E���|~)QS8ŭ�"�����9�5��=�	��N���� �MaV��I��M��WK��y/�W�_��ؗ�?
�^?cde�\^I�?$6щ$*��0�-�����2N{|���紀�����j}���V
Amhځ0j���_-�6���`<%F+�����V�G|"t��+
2� Zeq�a,��|$�S�y5��^�Aً�w';{�BiW�8¸��`,qo8�P����mW��rC)[{U'e���:��ђ���<˳�L����F������`o�4��h��J
S�W�3fq"0�/�����0���!�3bZ
���a:�<�J�P�"o'҄c����:�	��˵��H��y��ym%7-U<qqui��q���M��b�[����	gv�'ga��vR��L������X��$�������o(]R���J�e2]��[m��Z1�dg?��D�ű~�Z{@��E����њMkX�T�\�9��<�1Jej:�7�i�ML@���T��]�� �B�1��|M�e�<�!���J�tV��Q-:���^�a�Xa�u�S�D�Ě�m-(�6�2�ָ]H��h6qǢ6<4��Ɔ;W��Z�E�a�=�����|_=�RnM0�����Ϲ�h�C�?k��ݽ����&��]f��ߩ[��ʱq���h��@go..w'�q�-Yo(}��(7�"�����)�~��u��q�J)�2N������Ȯ�<�m�u��;�L'��!���w����O>�dgg����P�L=*q�~\�� [�78�E�w}՚�p��Jhh89{�j��l�D�Tҭ�S��v� ���V��Pac���0�U�A5����XH#0h	��>&��ֶ/^�`�C��Z77���H8#�}�EE� /��.Nn�6nHC���.��Do��|t_[[���|�Z����VЮ�I��B̗//��TV�=�������驈��C\l��R#į���s����*m't�<xp����|����r��ˋ��L$"֯���X�1ӊ����Ļ<�ZL�z���t�����&�X�9�L;���3��79=}�^��_)xe<z��Wo��FϞ��S�SЙ�Ć�دF���b�ܜ4ƹ`���=ɒ��n���Dʲ�򗿜i˼`g�-�5s�A~WW7tdc�,�@�+#&k�{｛�c�5���9���'M�=������`7!tY��l�C�������ۛL�DV���񡖸L��8�^m���+��֭[Ϟ=s�����{��9##G����/}�����쌙J��M�x�fj���4���e�5�,�5I��AL���G�E�Ѥ`jJ��M�c����La����߽���W�o�R@�x�R��j��`�i�L����w�4l��H$izr1;̽0�Հl
�^Ҧ��g[�n��f�v t�qcdM-�Τa
���Fea%�)Di� �}w��}����3z����'�(]���t�'�Lnnȓ�"X�66����K�����o��p��<D�I�4���*��
�m�DN��г9�ԨC�WQ�}�q���9cFW~w���0�����]����ڶ�sܕ��x�pr}Ѥ��Ӧ���ӵ
���߀�i
���m�������m�߉���9Ӽ���������=�]���*9�ݡ���V�m�<u��֣qg֡Ig s�=�1�� !g��^�>����=}@k'�.�-�:R�ȫ�k��E����W�]����\�3��/��= 1�"6�w��{�-�Ŏun"tٵ@��+���z��=��C2]�"��P	��;�j�35	��ʽ��;��Ţ}v�x<(�� })��(�f1�8w�jP ����N�˰�P����Ҕ�<覆̅���I�I�+�C������'�&X7�i������RƩ�M��$.{�7a} V�(��I3I\���仔�D�m���@f�D��Q �#�5-VK\0ٓ�X�o�}v�fy�޽D]��4�M��%4�WoΎn��Ov5�%�o=�e�v�vYfb}s���o%��dY̯攔Q�`���l��jI%��i�,X��P��3�QI|�'�� �(}^|�7�R-%��ʺ�&�>���`�پ�ڶ'�X(AIu}��%�LʪI��_���R,�O��܏{��͜�5@�fMz�y��e�H5��R"�����>��{�O��جQ����bT��|����O~l
���z������q���<}L��Ear!=�� �M�,U�ŀ�����E�����/EY���C����deX�8����a��bk4:��	�mm�x~H��p1������,�|ws3c�Oϸo{
�P��7�J�9�ia���N�z�͛�|�%R[|��V�R�x����ͺ���K��^�ǡ�d�!7?;3�?֬�0NR�>%�G�_�
|q�0)��N�fa���U1�Op�&9ͦ��L��g/9;ӫ1�׶���1���3H���x,�I�K-�P%4�r�'쏈�F�aD~i��}֋����	n��|��$#(W;��C6.'rE�h��lş�Tb�A�U�n��]p<@��svss|��k/-]����Ŝ����, ��r	uZz��/|�#������SE���&�.�_(���{N"bh�vR�I��V�ly�C�²g�`�]p����.r�m�C��qQ(�Ǉ@���
�=����^T��jk��O�5�}Wv���c�)��x�o��쭻9i�q�Xf��4@`X�k[�e�/�����Ԝ���W���ց�:��ϰ�y�u����lt��#��i!�	 33���.�tw�JVw��u�g��aiu7���l����zg��Y�.�d�;�����ht��hű8M*�~�iYF�z�}B�o��JؤlvPhll���g��4��F���?���뿎����80�Y�u��'y�B�jm˼�4�R��R�6��; �����F�#
y�*��=�r�3���,���DJ�+�jx����D~n�_`$�� �M�%���תEA�<ym�虐��3�Xs�q�L�c+���s�1�O&R��j� ��Fo6�/^����?$��U����H���6h��L�̡6���4�w�ՖV*�(Ph�X������)>aK|{�/��|m�@�s�8��Ɉ�j�>0X�a�_�58d�Q�s���Hz��Md6>3+�,�{�X0S��@D�;���//�9����SL�������l �g5����'A�	�DN_�Y�$'^�)L�w�#�����F��#�
l���1��ۧ�4��0�Q����zdB*w�ޞ��,�~�����h0d�.����F����-�YU���Uy�ݻs��U����uϿ��[�����/..�z o_���!V��|ˀEv���1mG1����sĂ��������V�� ��10K����x@�Hh5z<�4�;1O��e���\�T��j@�Ր�P_��2 ���x#��6u�!U^�5CI	�������N)Vk?�M���r홞W�-�D �8h�H{LCq���6j������` ����<ў���Q"��J��0~���FCӝ����'�{tUZbP�o��JŕTM@�F�"�h�:Q�Z��յ�Y���Q@8i�֪����w�\��j0�ncK��3�OZ��;�J�d�8�y���wL/]������6u_]���S�<Ȯ)�f�ŗ�ȢL��I��ڌ�-�T�)�(�~�ؙ�r�m������`JwF]��Z�oùb��fwtۀ-�w��n��������nC����ZD��D����	c	�	G�ۯ�G6n^]�q��}��M�m���(�+=�]�Tua]������7&!���1ﻔ�t�=�a��iW`ry'�|��@�k��j�χ}����<����ݛ�FQ�&T��.&����.5$���U�����@�FS��{���nJ�)��q[�Q������t����2!�N}��)0�� ��$3�$�yS���rAQ��ڣG��
*��5�egJ�D!H��0 rZ�z��͙���*n�^��$�L�+u���Hpޓ
�,�6G����g�gުG5�%|D<����V���
���x��R6�����t��,[����0y�v	 �U+?��c�6ة0Ǜ���#>ei-��uit��>z�m�Q�i�L�7A�������,ϳ���K-֬Hj�C1˵F(`9�ܶ�b6b���kЀ��KF��L� ���y��Vi/q)KwIIը2 �������>�������2�A��`p*�&�Q�e��d��=�}�>��X|v\q5�x��b����D��ÇR���r0;<:ɤ�:�]t���r�Y����׳�\d�������7�>����y�f��Ս��ٵ��/��`%w��������:�*�}綫�r����DZ�&���L�fQ&���^s6��yZ�6������8X�����1� �^?��,��+	$���4��x�Z2f���}1G�+I�O��N}�|0n;�I��t�R�ZiEE��iW��f����&�-�-UW���<g ��v�4��$n��TQ۲ھ��G���n�I�ҽ+%]�0$�x2"S����e���/����x�FK��`i�d�KO�%�7���Ċ�*���C��M�鍩N�^�q����=����
��X�����\-}:��.ttB��	x�t��T}�S	e�@�X���M���%{q�3Y,��V�
%��c%A_y�7��XF�fݽ51�(�x~,9�6QXc^>�'tzKW��x�ƶ#��fKs ���՝�ɹ���e�6�ڔ7�sYe�FP��z�m*Ս(R�'�$^O����ie��l�R`_~��W`]����.낉�%��� ����:��|}���-�m�%,f�v�u���4�x5��YC�����v���I�|g1461�m��\{L������;V�. }gݾ�g�'oõ�.n:V��u���1�l��g�_�k=��b�M�ݝ)�S`[�ua�;~�$<���Ui4�b-ͯ�~S��.�i�~nD���\���B=Ƴ�Z�U����#m/<�֭[89�^\0_���?���o?������|��8��h��7N�Yf��
T�p7�8�SjE4}�見f��O��C�i�&)+���*�}.�3,�UBУv2�y�C�ۀ ���K"2hm��h�1A����VAt���?ĸ������Ň�黪��z�����
�SfĒ��,6��+u����`�6�$�4�j�j(59Y���&�s����@n�ݿ�gU�l�3b�hU3�"���Y���1\%!�У�M��G�*8��"�kz�,<�P���hؗ�����Z@�ٽ|���O�޽�V�c�Z����D��+���� sx�+Q�	�b�&I���@`Q�s�4�	mh�W� �%��J.5�*I��X=��xO����↢ׅN:#(+��,M�
:\"\1^��9::b�2C����ZYͱ$�y{���t �m�A\�'��:�JANL
s��Ϟ=w�܃���0���c�}H9��À1$�9�
�4äX���y����#]��7oLO!�� �Y�U���=F��AӔ�N	fLU�v��\�Nb<q�|��?��*�ϟ?g���f������l����<���Qh�.;��H$�H,��kb�O�����Y� %ע�j�G���wE��V��I�����<�!q;�Ʌ��]P��j���q���53��-�?��J<���GS�\s��x�����M�A�m!(g��y��lǑ��w�d L�L>���Z�1�47�a�w���-��s�m5����w`��:����;wv��u�N8�g��JL�	v�\̜-�;	r3����\ԝ�;v4�vB����!��Fi�1ݫ���w޻����4;}����I��h�� e�C��EsK�>y�~�v\����㳂��~��3SE��i��4&TF��ö� � #(�r�u�~�Y����j�g�#s��	X3�)�'�|�W�W>\lĆ��$J^�6�園��A�a@8G $�(.��3�cI�Ҋ�N`�Fs���^���Ҥғ�^�-�ˢ�?K2�` �A>Ҟ��˫p��HkEJi�2b5�	���SV<�񬛹4H�x���R�E��SM�F�f��#(X)Ʊ3�hl/�v��5�p��P��djE]����z�H8�B��X�hj�a�����ӧgd��8J���s�m4(]���-Ĭ��:N5УZj)N�i"�Gx��������W�k2��S����޲,?�����&����`,���H��Օ�[��)�(��ji ���*�>'��@�����:
C�DEnm6��J����TG�US��a/F㱴R�)�>{6��������o�X��Cn�7�<PXA�͖ �R2��2�R����kh�^�����X�{"�����~�Z��SЪJPq�����ys)�m//�a{���������RZ;y1�e
� ����fVx���^�a"��e�����xu��Ý1~�򅴙����y�d��T�{�0��|68�X��"�HN��G]�Զ�x�`��=���*Ix��9c�Lu�:��b)i�88��$��L�	fu˓��R��n��5����H"��˕�0�zZ[z��A�lߢ���_��̲�J���s*WuUg�@�A檨(�(�3#8��;�F�3fd���#�GAP1�$*A2=D�����]]�+�S'��ֻ��v50w��i�O�����ֻһff�5�n�5�4p?3S&8&�'�
������N�t��Iş��S�դ7p�Ơ#mG�)� ��0a�@bЍ���H��}I��h�Wk�/U���?,ҡ���b�Xl��LL��N�;����`C�y�RnW�H\|EV�s2��ҭT��#XM���.Di�'����*�����	����v��M&�g[JXe�ۅ�5��$?Hy']7��̅����I�f��#�酺kR/553X����N͐W(�H(��%?Uc�TiLЦÀ��-���,�z1e`��C��t����$[�g�X'G�t~5�%��	�9�DNZQ�'#�v<V�	^�Tܶx�n�/��£D�����Z�UJ�I�5{q`
&8�D��R���G7���q|\���I���8��";�$h�����<��!�$lHB��*$������-��p��o2-�-��h��ۮu��HN���Zp%����:�����GK_"lD�B&�]���6���L�37wM��lZ,���F�Q�9����7�z����ۼy�ڵk׭[W(�����&���8��Z�4(��řb ����%<jL{<�
�ph��=a�h0�F��_8+��hV��=K���6�PW$�K�6Ҧ/�+罪�S𭶶"`a��9����i:\��4��'/�)ud�`^a�t6.@�=���Yq�U*6U3y���[�l���$}%R�A��%e?��1�����JUJ+\?29�h���-�W�Ęl���/(!'�N�T�6�n*���g|����,ŁG��\l�U��g:3�����\*������{�u:��݋���� �~���X�"�*~mKi7[[u	����@2I<R+[���U����NL&�SCJ�~�1�q��)���qÑ�>r��E$�#%��z-[�lpp�)bx:�u�����Ο�f������Ȫ��408��ݍ��i���9)[��Ҏ�2����Z�:���O��T��t��<7Ca�^�,U�-oyˢEݘ[�x����v2 ��}~���f�%73&s߾}40� mS-��Za�(��p��à�i!!�|��=���)S��>憳�nCy=�� �X37��V�3o���f���%��X)"�J��L��u�)S��QF1v��W$�R��b/�&b[�2rP����Ԙ���m�=�R㹴|(�Ld|�U��UP��h��r��a#��`�	D"iU����OH'1@]F'��,0i�)CD�l���d�	�
���p҆Y�b8����3#0Dnq(��V��$�8�)0���"oM���I�o0�Y���:N8k��2��2�79��f�C2�R7$��˜�z�O�,D��Ȅ�
�$hHBW���/��h̗��B�3b4➧zk|��y?������d���d���y��|]Q��p���"	h�_�Q�yMA W�W�c]'�}�����%9�掩����t�y��ѭ̉ǘ�b�P����r�{{%azr�9��X땩��v?�e��\�@kM� ;zj2����.,���k��j�昍���?�� N�QG)^�TZ*_]of�"�&χ}���f��1T$$j�F(D"��M����PB�^䥽4̸޹V�6$!�� ��i�˦S4�SL%Y�(�V��+ԣRJ��V�`�ˡ�3.f$�ep���E��ku?�z�W���Q��S��%�8�OOO��z5I։��VhgsrM>��7�JY�\�YZ��OHsq�Y�͚�(R�cҪUU0��Y�m�[����>:4�ʒ-��1J����T�P��2A-�-�M��]��ӳ�z�b� d�,�����q�Į�E�����r�U�Cøg�  |{QzE��<���:ff�wj|j|d\J�%7njzʣ2�ZZ���MN�Qd�AK"��, �Q��M���ј���$m8%�/>�@Y��|kSq���L�q��;0�BF�H���0�t � ��ҙ�R+�
N=h�UN��X(b��!�͏h;�t&��� ԕ�k�,J�D�&d|E�(ڻ::���n��e�jq���H���Il���}��&�`q���s�Z����7�g��Eڳb&w�؅?׮]366�,�t����N�+��}�^�T���Nڤ�q�ʌ 0�l-�߅SS���H=͒���j�0�<`��2x����ʳ�T�j�B���3�j�:�bs!
}��RQ�� o�Rj����j�$�eҹL�����\���O����yQ�֪B�Tjn��Ʈ(�H�	湻�7���4�SN*��8ZM
kĢ�Ԗ/_��48�O�٦�쌫a,�j�YbČ�����K�3�+V,��T[�ۇa���L�OoooK��?-x��+,vtta����0X�'J��Tu�2+������h|d
��҄]T�)p�Ԫ�*BC�ߴٮӿw��i�����,�695#6���Gଥ�@!�A��\T�7�e�m�c�c�S�/fs�0��,6����/���;m�]$���;��K-�m�R��.LO�{u֤u�D�� ���U�m`hîENg��I��lkS+V(���e���ל������;I+�a}���ݎ��J����i4ZZ�u%��*��r���4N&��i�ڤ%����M7qאH��
L�%˭�/Ѹ�������:Ҧs%���I�@T��D�B��ZeK���TJ�ؠ# �uo1��Cq��L��k������]e��`�g���|��`���͇ۜ��Oҋ�Y�x��Ȭd���i��ڮ�������0���2�H�"uϔ��1\:��ٔi�Bc+��h�Դ�R'���7e��g�ӂ&3������5a����]����2֒��8z1vqC-Õ�a ��FeҲ{��5e:p��%q��(N�m�ojS���a��[�d
i\'�����F�:�{ϮF}6�j�9/p�Z��N*A�5{A����"�}�t�h�*	W�f(�lP	���0��i����  � R�k�o��;�� ���6�p!k�? O ��W����9&�M���	�$��YPE�8�ԟ� �����\��f��w:Tu��2)�8s?b;d|B�\��)���b���fn�lY��$N�ૹ����*&�T���g:Z��D�'cBS���6���U�M4 į�RNIkE�#�"K�,�3�<ڣ�:��$��0(�(�� }lI�M5�(�k�F|�����m�	А��<�6�@t�4v9]и�O3�3Ąp#�&��+eŮt����qi���lm��c��MQb
 �h�څ��v���_.���4�C�v����w�D'9�8�&����r���֝I����mbo	������/^܇�ٽ{7]�Y������)t�Z��V��V������8�BT���b� �	����k���MMB��wbFךq|c���һFZ/j#z�]���'�D3ω�N��?[���L�Xssh�Ds���k�՞]L���֘U6�� ���D�&��t(���el��קC��:R�i�cip0f���%���sr��nz𖃃�Z+@�,~R�K�����9W�:!�������$����'3���)�t�3���8x��ac��oߍ�w����_I�b������i|2:>��#u~稌5a�4G-b��+���꨷OWPVA� �J��Tɓ��4櫣��W��7�}4B�9�������T۶��&�Yg�u���u�q&����f��[�T��&H-�e-?����rM-��s�q�(�s`J;݅/�U\L&N��@��>
6�g��y��}5�4�7��%=O��إ�:ה{{˦1�q�fd��B��g�JXZ��.@��u(���w����uk9&Y��)���0�ȱ��G�Ȍ��^����߱t$�%"��~�lJ�E�0E	#L�u���v���L��?�`�K���{�%�~���Tï��1��q};M�0q�yg�u6;�b�7Z��PT�p�=S*�M����Z�qOHf�[�[��ؿϢ�@i/<S[��&b4ɝO����Tҡi����)��<���C(�uz���գhA�'���Lc+�0X�İ�c$�5�p����B8©�J۸9���R���
)7���ig8Sj��[Va`���;Id<�DV�2�D�f�7��IS�	�:ꍥD��L�p�2T����iѺ��eL�W�����'��K�F���v�\�-#`z8O8c��H)㡜.F�8`u&7)����`�M�Rs`���~�mm�L����Ξ�"q�DBU��q�Ȁ�v��aS�I?�F���dj��R��Z��7�X�,e%���j�:�$�ӱ����҇!iդ[ p��8TND����v:���"�X2SG��\d��s�L�C�x�Ȑ���gʚ�0�ΕQ>g����@���XXٔ��ci3"z��jt���o�i۴�@�?`��ӆ��Z�K�h�:�ǉ�p�z-���ܲe;��hϞ=�� ��+�޷o���v�ո߸٢ ��h�l��H֦J� �g�9j�+�)��v�>@6`��a�0cm�Czg��S\������Zλ�=
�t�X��*jD�\�Tu�?�F�OMM�)�X*��wu��� ��k�����\)v���Y{��_٪���t�P�;�
%E��&�l{��m�	L?�߻����5�e���k׮��?(%�r���W��Bqa?U2�*�C`ԢD]��NɈ$g�n�E�n��U>(mxU�{��$+����ڇzY��k�)�2���6����d�2��Š�og�A����X��w����aB�<B�PUՊ�ė����S�d�y;�ት�eϐ<�1�����YZ�6L�׎��-Jd��i�YN`'Jt�TC�a�~`��`z�.�ȇ2��/i*A��.̜�M{M��4�^��&�@ziZ<b:=��q�<�^�x��Wh���K(��;�������4����%���5Y���cN�B����}.j�)�t���+eXL��9��UC�IC�p0_���M� ����$B��L|C2���s6��ć"��E�H�9:2?)A���H|wbk�0�y�]��&��cD���kס���|5�$���=J�pRrIM`�ʦ ��_�xA,��\��Tb&v��x��z*)]��h�e\Vb#f
f�� �g-PkH�S��<u�g�T*@3q�G4s�a0����8C� T6a�h�z)���t.w��a�'��Jn�1�_5��謢� I��(�Fd:::,�p<��������(szBe��?b7��l[[K�:�mp��e�O���AEi��]+��@�!9~<��btR˲����tE�sF��Ԝ��=8��,� �3���Yn���E�L�vJ�/���J��(����=��t��a�/[c��T�eS��ϑΏ��3�Ͳ	<��t�ޔ�����8v�.3�p���'&*�仫�.W.{չ������l�.�R��6��o�(n� u�&K��;�xq/Ӥ0 ��
.W�^�l��	׼�Բe�S*K$h��f$J���M�6���/^�X�R�R%	=3��X�?��[Z�5/��⫯�
���K/��;�w���u����C�)�:I��
ʦ�36�R\���O>�aÆn����Ϥ�J�<7�Ţ����KN9唯���4vvJ�ȈԴr�Y��*��a�`���<g����%�L�T���ٺ_�(x0}���7)�j�y�|�uN
Tq�B��~�����y��d>q��IM��*D�x���J�ת�ׅI��%R���q/�i͞L���ש(���T1}��y�8�
��'�;����5/WU�&?H���r�U�<���'5�U20�~��(�^���l��+��
��ݱ�M���dF��Ep�Hn�� �Q��5��n!����:��o>!\3۔�9���33�я]H���3C�����:](��5õ'P��"���)����ɪ�?�6D��1�d��Ykâ4�$F�E�����Dsz�I��J+e��SQs�
�߅v;*���e���R�lq:}lt8�|�1< a"[�3�|�H]D��ry���F�(�<�*���8Q��)�/`���ɼ]N51�O"�A�+�W�g�V)�>�ܵ��3���R���&6,᷸�ԭc�A��D�=-��:�cc� cX�H�hCZ����&T�3�ӊ���P
��m0zH/BZ�1�<1o�EnЈ悪jG)�#��I�@zѠ/I�J"\�UJ�5�1�X6�hK���qz���ﳳR^���T���C����162.A�|�+��t�����Kg���v�G� (W����^���*�KSS:�i:�ji`D�~�"C�âb�)��I����0���|��Q1[�G4O��PZ��;eu�r(�dw)C;�\�^�7ZZ�E�pj:�i�O7'��#��T�fܧ��m``OLa����G;�[t�)^��ހ$��\���G�s�k�&��D9���q۶mk���A��:���٪T�8@̲��_:;;Hi!�Aϑ�L�%@�[o����3�7�uz�����,_��.=zI��?�}dߘZ��/��=�ܳu�V�'��N�����u�RւF:�u�<�9M�M0=�ʻw��[���o~�Ԁ�Y���<Z�r%���Jt���G�k�4 ��$--%��C=�� c�>�\o���5CD�ax��q�Ƨ�z�g����?}��uħ;kS����c�`���ã��L1��Q�?2���I�goH�ݢ�|��M}%Ҍ<>
MR튴!0gSv; @��'�_�b�ʹ���B!oa�.D݆}� �Q4������?��m}C&�xn�o�/�7��Q�ee�^��N½dc���������wvL����MDN�[�$ህ}����M�H�k�h��� ���0�43]V�U�z�����Pך�Q��/�u��]jy�b)����.���(����%��a\�ۘn�w��۰��j㟐��������s�s;�.�����B$g��H�Ҕ��p��.]Ԛ�;�ό��M &��z�������a�2���n"�j�!�� ����M���z��$R�*���6:��C����ʞ���$R�G'�5��D��gB�6ѕp����I�"5ǉ{�j��8��7���"��<T�sz�"B=BX�h�o�T���6�m�v�qN"��Q=�\���)`a�<22�h�ϒ��#����z&r{P���G9�C�3ɍA��+��
M�)��:�n�W���|h2hgG�X����'j��!����x׆$�0p�9'�vŅ�Ymg��9h↲���[���M��s�L
J�+�cS��Mr/Q�q~�wH_B���'C��G��-r�KLMɲ�XPZ,�S���ɧ��W�C�By�]<qhh�Ǔ�G�d�)%U/�(7-��DI�/6L[O >�3�
ۃ(?4��}HE�4�U&�'K�-��ô2�4�G�h�tw��Vai�8���#�bx����c �Qȶ���k���;����_ư?�p�؋�bٲ>G�N� FЋ��	ؔ�d������ۋ�944���oٲex� þ��~�E�]�I{{��5�|��t-_���W����?}�G�ɱ���V�Z��s��+��x~>�We/ |�aÆ/|�� �Z���<��C �xǴr��t�d�S����}��� ���կ���Z����:�;:0���6��m�����w�K=:!w���p�cB�;8(�k�?��Y�x�����oa6p��kRZ i �n�Emٲet��4H�;���w�{��b�)hpF�af%��81��ںttU��	=sݴK��.�p��٥�1qZ��a��故q�[��$��阷y,V���A\�Qk#�n莉KZ�hu�հ�ʎEB��)mH���ׄ��?��'Q=j�n���8Ytػ��D�1q�$��������P���ye���τGՋ!�m��7�dP���׾�~�����L�%~�i�Ք�[t��"v�v����r�C�2�"�n:��v��W�5 ����vA��͉+k�#��͍$�ҩ��oV�Y��)be��|
!|6��:�?��8z�œ).��<�5iS��aAh��9���'�f��j��T�ҩə�j�><:��E3ق8Q�&��J����S��dm�<wLF���a�8���3������@�R���5�������ܬk��6R�;f�6�`�kGE��0�7����ߥ굕M̒fR6��\�j�=�4gS����;OC�33q�㙙9v�! #b'��ި�U�\�\�+���|?39)�7�FSZ�c��pQ����
!�S�"�,��B���\dF��!����zi��+E��Q�s���c���!�-2�099n�ئS�׊��19JmnoFQ9*zL����}�;{0UX�bQ��Ş"��ֆ`��$!Kgg;�466�J�3�!{�zʽ	ݼu����~��v�"�=�@�ݒlT���< ����%h}�s)��ڴ����}-.�W�h�:�£ϕY���0��n����}Op�IC'4�ת�7h̔g�t�1V�a��裏>�c�.��Z�n}x8�Gq�駟��۳m�.L��5�Z[��4%�D��s��+�0bߪ��ŘF�b��9�����	�Փ����͐��ɜT�N�r�=?���y��t*9qH˦\�_�^}QVnh!�SqFGG�0�ή.���4��{�a��)B�%MI�lD��Fmھ}���@.+���L�&BQڤ�����g����[n��^{��8�C�:/K��/������'�!!�.�ʺ��8�%Ig�_$�p���_����?�s����c_c�n�x̂�5E9�x�������\rIWW�6�OY��CuC�`=|6�~�&����������]F�H��>2��N�PP��C΂<�yFo!+��qk�%i����(�L���iC+���Q������D�x�g�������b�Ր�r�Zv��ut%�jzsqh�DIcI�vP��B�9�)|�T6�T$�Q��)ٯ� J{Rꆞ飼H�O�Э6 o��1$L6$ ��BG�(36��O�-ز�8	�I3��ثCr��ߨ4Ό�h����.��ʯ�xQ´�8ʇҪ[{�$�������"�b1�r񗹿mM)3 b�����;�D�2A�R6��3	aT����s��L>w�T9U+{��� ��֭;J�<C<x��������*pGe���Q"�U�2TWW�n��WQ�0T*uV�ؗ5(i��hR1�j ��g��,�=ř�Ej|e�l3$hM(+4�lH��0�A`rT}������u�6������W�Ξ={�������y�Rw���UĐ�4��ҽG�A��qd\�x���N�Dr�;
�!ƀa���A4(�_e�߆)Y��)F��=L�2�
o�(Gjx�
�!V`u%9��PF��W��f2SJ=1T*	ӹ�dJ�֜��U8���c�j�!�#?u��~����cQȊ+N;��ŋc�v��K[����ͮ��F6f	�[���� �~������K/��A^1����t�u�]'�!/b���~Ѣn�hzK}���ˁ[�������hC�A\d7���T�q�� <A����?l$駳D�����j7NZ�\�t���FF�'��n��;�k�֭���x�k*9W���ꫯ~�+j�Dfǎx"nj�B����瞿��~���a_���u�n�6����t۶m���7����}�k�v0֐1Y?Q$N���ڼy�/���;��T���d�g�C���1�3�<���|g�M�FFF�� ��s*�65�-�
k׮���c�bn	���LBo���Kg*6'�������SN���Mi�j|l��*{�`Z�D��s�SO=��~�(�<�km�V� z�嗵�{�fd&A��[Ĭ�A�ͧ�g.����o���|�Ru�>fO�HӞz��2������`������{/�;�X�b����۔��0{Y[�曦Lc����.�Rh��7��#2� �5�r	�L��0u|	�+l��#S+joN	B�g��uX�e�D;$ϔ��D&2ET����6uznL�S!e�^��۾���M�D+p^7��Z��&��ĻQ�!#��H�$<�X��ճkd�7��1�Ŝ7��F�$�]�%��,��u/ѿ#p��{��]��v��	��޲d��S���8�:xݙt����x�mĪ���Op��'�|9��W"��K�c��b̄Q4w�u�g?qq��!�(/��x&�	�Ӝ�Q'��Di6,�	���<]*K�a��6��;N�[[W�3�S`3m�Nϴt B�#<ӌLN��_�y#ۅt�n*HJ���MTӹlK��⥃]3LN�ׄՊ��բ��..�x��H�'Tg
�(���3T{�%Iō�3I��n9d�H��zL
/���@BĪ��6��&�sD���:�*�3�^�� s�Ƣ�E�m�|r2f���|��ꃂ�5�
)�)��a���y�`�hV	P���нL�M4��,�ZY/F��	DWi`q�
_��ǝ�!�L% ��ٹb�g�R���Q�`�IM5��o2��9L4[��&Xx.�U�r ��iUr����7������@9m-��[n���K�ׯ�*�۬Zi*4͖g����ӟ��?��?-]�W�a��JCӼD:c$$��K�)V8FZy��
�/~���/���I+�e�;w\s�5�0���Ė�$N�l;9).���$=�0{��{�����Mw)�{�����l8�	�G�9mZ��%	K�fX����,V�#�&�\C�J�_�� ��8�n)��Y�p�������M�K�'��a�/���@�a�!$ō$�L:w��J��㩧�9�s^z饸ZY�O�������0���?��w���SO}_6-�*��'g�h��H;���0ܓO>���v6Ȃ��`fV<�V�b��]�v�}�ٷ�z������:W�H*�fA}�����O���+۷����	f?��,��4���\!��񥍸��T������ss���L&���T,Dn�ͥ󅬟v����q} ���N�s�jn�tQ�ʮB�0<4�"+�71!���܁�}��ט�������wߍc��+X,(����h���0�	���dtF�2��@�����d����m~��h�I��#�6�A�P�B.�A�/���^b"^o3���c�ͩr8b��2٦s���dލh ;�C���8���kHh�kh6gL�R�P�8�+��0�����P.�����ɦ�2ɇ�����*�s6����wg,�Fo,�x��}����%m�9e$�'s#�	��E�uO2�`�QLH�J�����6e�3l]V�~B��+����BƤ<��a����(�%�bPS��i�+�e7n|�'^ye���^{ͺu����}���V9����&�On-��>Q��4xԱYvݝ�n�)��j�|qtE���K�i2�[(�qd��[*�+�V��J��a2*m)�� �vPg}���w޶�C��?B`L�4z_��!�`�ۄ*��x�d��k:��0�<����G�^�����[�����A.�rYt��{[���'�"j��FE��z�ǀ�b�����G+�?�3�0�ݻw��Y���sC�($������6L�J�;3�qv�ĖZ�|)�<'E%d}��xw���TX�f����J�fS
vC
N��g�r���f�L�j����I��?�ӮsƵэ��Y0ȃ�kF<O�CL����P3�}�������r �`�,���yD�0���Z�|9���{�7д����  U���|S�n����s����r\��:� ͼ�=��_}���R�����Or��&�:����~��<����ԧN=�T����`�&6��������}�ZZ5������_}���Zu��5�"����8N�j�T{�&�3)8�]�{��\X�@�tQ#Y�k��A�o��z�5���^\}��XA��$P���>�nm�Xgw�nQ��ACC`C�CZ.^���3�^v�e��P��"�и3��Nc�����/�;�իWk~BKss��42)����������SǱ�X��p8��Xnl�;vl۶��k�=�w�5B��X��������/@�9\��=�%ir8c�pX������X�c�9�>c��@�۰^xwr�`�:Xʋ.��2�ε�k� อ�J� _ٲe��~����ܒ�K�ڋ1�&'�x"@!^sȦ�A#.ߡt偺��q1KtəG�����)=HL����9�<�MK)AlFI�[Z�o��6�*|��7�mq=.޼y3�������x�E���px�SO=���c~0N(<b�&�=��3[�nݸ�k�r����k� ��) ��^`])�R����֟�r!� ��N�d��3�t�i��0_h�׵b�I�L��L����j����Lƭ��֭��P�b�,2���4Y�@Y��Rd�ˌi��C���4v�r�/W��-�J�I��Mb g!��H�Kt��l:��c�� ܓ�|��J���w8մ*�y��Y�N
�舵�5+|����M0�X�/VϽܟ�t2iw���o��6�Dl��r����7��}�i���;!R �\w>��5?Q��f�Ƚ�{Ɏ�~�Ĺ}��*gRi��� ��S�ggk��P��%��7�W��'�k�O���k��r�F�Ne!1�H+�%�Hf��n�Յ-2��+B�u"��4���LroA�}����D	���Oj2g���z�s���Z�$�
I_����N'�v�B�4.��ޔ��2�p)BRQ�K�Ķ���͋wch�� g|_9���w`�>:e��m���{�,nX�)i-��ab�� Q^�<r��T^��w�G!��_�PĊ��9a�=��i�R �T��t�<-+;�	����V^0��[��h�(MCM��xf�3���{�ҥ�R~['�F�[��vVo(�bMMEaџ��0�f.�F_�u���?�<T����LyF8��n�� ����(g��y��|�y饗b�%ݾ6;6>�f����3 �=08��������T��2<�/h�N�NNL�Ď�V*�lNR�����ި�Z��9�+�eD����@������kB��aR��[t"��)��Ja.�%����0�5�=ݽ/������6ɥ�.J��ʔ�5�2l��1����/��;���zJ�вeKx���~���Y~�8��$F��	1�mK��b�8��������c\f�{�iγ�>�����_�����cZ�816V,��.����, Ĝ ��X0?Ry��u
%��3���W�.����k�Rq��c�&����ǧ�~�Ӭ��޽{1����'X��Bi�	qgdf�Pرs�U��c3�=����Iw�M�ڹ'���r�$�e�&�+�y�����/n|��\�����";w��\����__���C���A�����]1��\r	P�x��xǨ0QX�C=+�mB
[��k)���!���0�&ϝiY��DN3��!��Z�iب���x��4�c����������l�L^?�Ë<&)Ӆ��#�L���%@�é��+���� �P�(4+X�l6c�[t���Uӣ�t���mh�iѤ�鿞a��AI?A�&�8Z�V���$o���#�L��<�i%z6�{�9��i�O⩓�y��!�U�t��^1��CҶ��PF8�L�����={�^u�U>��Ȉ�G�a��H�|s���6��أ�~��_���˗.]b1n{9�(�~�#���%�²nn|�|����m��
o:����L���]��ח�*�y|�%�՝�I��<ڦ4�=�k�j�
�G?������Z[##�ҙԟ�8N#����iu�X�ic��N�B(.<���k�m&��ؔ�Z�?1��4?TZ<N���3j��rRIW�,&�3*q�-7.�+�d��3 �m`1=��T��ba�i*lQ���&Z<�Z�3"�ה�3�]wy\KKCS$B���L����9�������5�N�2��@a���<���D@O�Ey�7%���e9��k|ȰG�7���Dы��$w�Kk��}��E��e�����I���g�7�[)���-=@1�<s��߿z�j���Q��{���χ.�袋 ������/�3�)j!����]w�%w��GIFy:>ɸa�R� [�pư�w�q�/���d��-A&+��#�<����$O�o���1k�F�|.^�RsǓ[_��bq���D�m�2ݥ���������_H���Mz��qە+V��_�����U�W��VC�j֪S��8�&�@�Ai	<�?��Yg}��c�|�Wp"��8��_��_ \��(�-��bї-[�G ��������X�]�w=��'�tR{{��७;���������մb��a'��g�u`�3�<�_6LOM-���Da�i�d˄�[p��Ӊ�S��V۷o�m�2�u���t�nrt|| ��|�J�]%|~�����~PO�� ����t!Za�1�'�xBC�����b���FL�s�=711E�Gc��<�̈�@r�x2$���-]������!q�����O>�] gl#�ÀbX��N;�Moz�9��d���a�j��֬Y�jP�"��IY��d�hɚ���
M�E�d�'}?�K�m�I{rL���{���1���0�!�W��1e��
h��W�Lb��3@���r�AP�}B��I31�Z�-w�ߵk�t�֭,�ԟ�kמy�}}�0
X��1����O'��Z��_8Z�P�(Hi&����}y���O��5�)f-rH�v�I����Yr�1�~>$?Q�`�c_��uxh�;��ν��{�Autt��1��q4��o�>��-(��w��?�0D
PZҕh��F�m��l�L����Eا�bs�\��$��,vM�؜��E����R�ؚ�X9���TH��"렳�D�Z�dC�1M��/�a�k��Od̹���c�σS�YV���#ES�[�&���.G��fM:�C}ː��}��v��5T�)C��� %ҔYޡVM�O\Sh�?=)5��k��|(''4)ӫ�u�CCC<K�ykm	��s�:��9�����B�1��b&F�̴#��pF�F��U�T:nP�3��#�i:��Z�e�k�ѹ�M��GG�,?\�jb�E����z.�)�7���M�iqM�/ދ%��(��{���l8��a�75�9e;K�?�S�\��jq*F�dI�ҧ	�����������ݸq����O�A�u UR2������Yސ�Gq���iO����+[��8&?TU��дa��?����j,bȥ�M4b�\7|�[�rjZL�c��4*�
E�D&�ycL�crA9���ԕ^�q����dѕ��Q�p�\h7��>�a�(O3��=M	��n��k���`/�a����Y�nF�ϯ��
��Be�Fj�H��a��=�H�ٜ4h��x�O=�f8 s�x�b,����W?��O��e��e�=��c4�RZk�{˖-z�E$в�����ﾻ4��4�d������3�8�R��o~s��cؘ=h��6N�C_z�%����}����3 E�����|�P�ϗ��z{{FG����͛7cT�҈@��ر�	`�3��)V/�����8����-��i蟽���i��Ѭ�c�����p^C��1�扉����/�����ןz�_���;�q��Җ����=��O������9��F$���ߎ��M�X�@��pM�j�L���rҲ�,U�����*�+�X�j�����A ��He� yq^����0�d�8�s���ZMl�xy��x>�I�<AC�
)�U�Z��{���uD��y睏?�86�	������q� �A~���Q�r1X��ܴ��]K����0Z�gK�;���
A?��7ܰz�A��w gҟMe��d1T��>��z��&����v�Y���My��L:JƦ3����7����`axGu��>�����Y�c)q��N/&���_���Nx��ߞ���O��NTr9��ːE���-�#�㺪�J�V�e�KK+�jm.��¬�y���,.�&���f���9 &�4!==�b��8�h��C���o5��L`50%�wm�Mճ-0�Q0�3�m��]����U��5��=_^�oRq�g:�+#)=���KW��G�@�8�Q�J�Sn���Օ�i��_��!e�*���|�I�|!ɪ��Y�dר�(g�HB!�0��-#��{�)�R64�;{�$C[OZvf�9!h�3�Q�[���_�
ċc^�O��@�(�(�"�̨R������4L=��e!&
�h5��,`:'��=E�\�`E*mM�900��َ�a��5s�(�Y����z�ÓG70�;�&۷��=q�a�U_b5��^|�E|qϞ=���7��+�9N:�$�� ��z�h)MZ�3�<�w�K�I6�Nō��Z����榦l�\���!���1���}�:���s��Z5�x4���� �\�3̐J����_��rjj����|���=V7e�)���ʛ�l�YҥAi�����v�l���q�ڦM�����=�w�Y��Χ��ɿ~�{������c�[�b	%`�7���`Xַ��g�'�/3�1-�+����<����W.��ҿ���[�|�uc#mذk�5e�564\�p�\nٲ����>�v�ᇑUD��(��g?;���p  ;V�\q����>� 6��<�0��[�W�r��o(�cdxhTp�)Ǎ
�;}شsp���G}��S�4/��;���xL�J�����c�i�������	ڷ�3��ٵ{�u�]��/�rK�W�n`z��W\q�Tl.F�����3��:�cp����$������EO��'���ꫯL��UƵ�^��;����X
+'B"ڋL�d2��*E�&��-S������^En��ٲ ��m$�1�]�G��^�U+��i=��ʵ��zԬ��z+x�o2�%tLT�a�MG������ó�>�����:ؽ���m9�2Z��P��o�馛��8�|�;?�����S�Ǉ�K־�)�l�6]�D�v]]xD�]t�=�\u�U�]�l��GW�XAՌɣ�p�yz9"Weh��,4�p����"⤷�.��؜[,�������;��ppN�����}�C�>�t<����fX_,mb!��[����`���'�]�p���F����AV��d+2��nXp�`�5
N��
�2I���'�&~ȯ��r� �:��Q�����}�t����艹_��WZ��;�3�6|�z��U��J0��E!tr��x���$���X���,���:mH���D��u�EFd��=�V�W���Ik�t�� �21M�cڸ�jb�@���d�l��DSN�p|D��oO5�&��NDN��2�rިP9o�`����	�nM��Ǩ��B9�pL�)�R%�Z�E���� DF��y����gu}C#�L��#CK6�k=1�W<���xs�\S�n��o�7��s��=M[�)����0]�F:]�pmc�Vt�r��'��F����lw�<��c?���FG�,��wh \�v�Z�ҿ���:��}.��K.�"u�Ν�=^y�����tժU_���H��:\���{�$ݗ*��m����C��a��V��N����f�v��l���F�
˖.�d�xdz7џ��\399�F P�0(I�R7MK=S����M��Zbe%OG����'b'��b�dSO>����<�?3WƉ��������@��744�w��������ܳ{����"�no���iv�taü��tʱ͉X� ��>�N�2acٲe`ݺ��䗿��ƍ5�$�#I�=���(ۃ�@�>��s� ��6�H�E�7����fz���}��Z�?�
l���R���'&;��L[Lp!��R�ZX���5�}�Ε+�c�q[��jNT\�g��� ��\h�u�̔�{�
�H��Y//k���� Z�(�6���SF���w��L;4 .���5�x�?����r�T�E�Y���-45�IW�X��O}�k_���Cae�5k0�A���SLUW7\��t:�&T�'H�>���Y�!�t4�]^���U��1@Y%�zZ8e�S�4�ؒf��QsLl�~�a8Z��k�����L����3ӂ��m�����x��`��J-�bw�9�������e�Ō�[�u�]w�y'�^��O|'VV��
0��x�DŢ�#v�8�|.�����k � Ķ���W��U�����"�労��Qۘ�Э��.��Ib��oHv�eT�ф(���˨n�Y&�8��g>�v��R�h��\�|)L>��e��g���^�����Y��L��(�"f�7ԭ��^5�2ykohF�PFHXL6�~P�u�q�Oe2��FѡE�
/|Ъ6���t�����T�Op({&�+m
��d7�m�QǓ&�,kL>�XiB��b��2@ü�F�3�Jl떖恡Q��ِ��>R̥� Z-�)İI��Im�k�i;)A�Xr������Y�R�Bv3�ǒt�>G�Y��� �`[F���]�&	f�a�%�,�afĴ Θ��\�����p��}�x�j�SU���5�V4X��'��҉X0F"������DiB� n�O��pCuPg�`(ths[i�U#�>nB��J�ysGG۾}��\�$�C��&Ql����nh��JeFF&Hͥ��۰�Xb�Zc��骁9�sN;�3, ���g�=�\HNG����?�^��c�������(�J[�n���6i�$;$�.�Z+��w^K�g�UHr��g@�ڨA>.^��Д���͠��x%k�F��Q������H��K%�rul�-\ƳI;�9c��:E<�xq�/�q��/�*�Ft�M.�nK���#�0������O?{`�V�(����Z dyï�CH���n�X�H	t�-�pK����,�����k�����uI۱�i�c�q���`T��'�|�Ŋ{��p��-[���|G
���:�ƃϙzL�7GmH&�a$8
#Ò��}�J-���ԑ����Р�i��R��ØR�P7�t3��\������~�#Q{�
O������"�$��t�M�E,+L�d�]�̖��Ag���x�6��g����n�ZM�z-��l�4,�P��z{{�X<��֭S�7��8�8���Բe�m=<<���uB1��C�q����l��GH��z��h���*�56ݰ���s�:�)��T�z��eG�5��\C���6�9'9)y�Ϙi��I�b�F�����6N�0��L�6�T�[�
!#}u�bnz�r�W���Aƿb- �y	�$qFu���|��#�<�!��#�<r�=���W����>��O~R��ɺ)ҭ�L}�q�
v_�����o~�E)��x(��[o���SN9�#�:���.0DkU��m�[8b��E��an앺2O?�4�)+�`������[[�t�ך�b��?�\,]|��_���1`���T���S��K2s^ӊp�qꋈ�V)�55�1fމ{TƀϢ�53U�733j�1���Iy����u���L1k�BM��5�x�����w�\���=ʲW�2ĥ�2~��0ѱD~��᤭��ˤ��9�޹�b�)+��FMNx*_ȋ	�X�ن� :;'��0�wܔ��.���� ?�W���{��þE=���4�s����KyN(#���5�N�+W$E��|�\�T�*,(q��3"˂V)k��槫�]
�K%������EiUYm��tSwώ;ڻZ��"�j5OwX�c�"��*_ϔ�r!���4�N���p�v%��U�+Z�-��j+�I��. ��$����N�J�JWW0�#��ur�|�D�L�IB���#�#^��BJ�x(��=��T���{rr������c��Ł���.
�)�a7w��9��!j$n��c�����Os3��ym�X��Z4;;�H D%�ă� ,�F�+�fd$�t���)�a�s:�x��Pc���a�ى�~�P�NN1�+r3���}����_��\���w�-�� ��Z=w,��o߶[�VgZ*W ���:�,��*���XV̓���a0S�#uPK[qO�����%�:ݖm�b�QÁ���Y�d���M��*��E���`N{1u`?3��0�r�XlQkD������g��l�����$��8+P��|nbB�i�;Ӎ��Rh��X����7�`L���d]��o~3 �#��_~YFQ=������Z�P�N����֋u��kw�.����a��t�s���C`0t������$W4�&�KsSӪի��fv���^y�?��O8n��{�gߢ^`�l:�?�&&���+���gI�R7�j�zMD[[�''�_޴yltB�H����`Bj�6�D�2����m�n�[ޚ�櫲���Ro����w/�wI�[y �q(�a����H������
4"&�H��I�3�#����\�Rl*y�_j.B0�ڽkq��+.��G?�l	M	�`/&,�m�C\kr ��'���������K�o��w��|��Ĩ빳�����~��z;�f��FwO���vlN(�@�ؘX�p���C�`W�i���(�W%0�=I��G:&���aG���aF'��H�f�AR������0\� ����M*���0y���]A�8]S�2�Ʈ!u�N�M{4z�m�Ҧ��h��z�)b�p�C~��o|��G�/_i�ͮ];%W�*�C�(��鉩�i�I57����S��;\*�����Tb��/�g�\��/������<���%�t^�����?���_�{͚5dh�,u���Җ��xӪUk K1+�|Q�5EN1����/(�AE�/�Ŀ���V`ϫ0J�$,i�z�������W����CACr�q�O=��\�������n&�7�#Pq6׌�;���w�}�]{v�V{��G^���Ȫ��$�!(�E���@��� .� 4��:X@_K�S^Z�LN>��i��[���K��ĵ��`�n�\*�O�B�i�MqGKR[��&a`,����HJy��g:w1�!�=8���JI�b���Zh�W[�a�7�U	9%�-R�=�l:{R�|� �������OB��}���o}�����:���r����d��O`���w1ǔ�x�3{�W_Ë�j���X	�<CḂs4N����z�!4��x%�100@j1\�iӦ�:(��@ �2qs��ŋ�twdH��d``�L{�}r��&�Z5�/�usҁ��z�ۭ+��tDT�����>GC30�{{ce�/)	m���/[��^1�2��PI���4�iB5|(���]���t��э�<�)9c�ނ�ga�Q�R������d2z�0V6��� C�s##c�!K(�*��c�p�j�E�{�{yk���DN�_�F[�&luhgC	�s����y�q�q��r�-c��]�4+]7��'���%K��r�1�ҥ��]��O<Qh��/���1E�>�h{kn�D���}��%E����tV�.���Lִ�&CK�	F�w��FGFx"v����-.�P�s%��]>��Ւ���6=g턳_��|�ԅg��k � ��x�	�J����j�U��&K�.�q�������r�c9��O�=>;�b�f�E������k�T���Uy6��=����/�&�Ӓv�7��/��n�{��{�{�|d�f�X����)������'��«�K����tF+ z�
���pc��31�`젃Vª|��0�瓯����>K�*� 5��ݧ����ր�8&I��4�=�3N;�n�I�	�����(���6���WW���F<}����*�`�[��և?�ap��0m�d]����<�Ҕ�U��X/H�h��<�Ѧ��2�y�g1�yI�D� >��j��t��`+4ŀ&?��m�ɺ:l�50�h,�L�_���0잾�<��c��g�B�ԽX��T3���w�����/��ێ=�h�Mƕ����V�$�:�	�D��`J���Q&V���BZe�5T'v�g>� ��}�#g�y�FbI˨T�о��'��z�믿���l�rS�2sFi�{6o��]�i�pڴ��� wa .��\�ha�׽�N &{vZ�X�� (�C9 ���Qځ�5����裏>������?B<������o���/�������6��E^��x�������a킰Bw�u�r��3q�!O�-��J���O\?��L*�@�*u�v��5qβ����6C+J&���7�Bچn�EƮ�cjy���򆿮Zu ������}��-[�|��P�'�x�c(?x ����C]-���ޥ��	<9��׹�:R��jU�Wp ǳ��;��px$=N��\=ì�FyN;(�0��[JK�������[�l�)��NU
Pu���!A�C9v+��3I^(f���l��$!+�<����1�ȩ��377�4��B�%���R��4�BVO{��шZ%�e�O���[	�*��a����8�+g�{����龥3�a��:K>���s�o=����8BbJ֩1��j@6c~��ʧ� 1?6fM�*�љ�"e� 1)�Y�z���U�k׮W_}�HL��.]��(�vIO^��0TM��d����.�軗\r�/�<9��C���o^s�5?�������5�%�G�e��b�k�o�3��SpC3�>�՝{���L�^zvf�
Ϧ�[�����5ӓ�[8�Y+Ϫ]�v���;Љ&������cלz꩘&Hy�QՕN�Q�	�υU��0|~�Gz��J��gj������@i�������mmő�l�0o��n�)�1 ݱ�i8q0|�%ۉ{�`��j�{��>�9��C/����3�Pt8�H Ƌ0����<8(3����V	��k����/~���ΎN�F��:��?��xD�5�+��Q��[ߺ��^�w��������|c[�v-� �|1'\O�0�$_�Fx^b�!v�ȹ[������"-j&c*��Bظ��=�:	�z'���D��c\Y�)	�آ(m�H5��1��P�X�e����SI�k�����=7���351�I wn"��j��a�O�8ߴ%�h#��L6�����7x �ӎ'��p�(�s�X����;/^��+Ç��Q���!OJ�[���q��Rd60�}����?����쨣����0��
�D8�j��='h�;w���{�]у���?������sλ���B!G�dj=ga&�����ez��^�����E�������ptT|�CCg�}����>G�?�~I�)	���Q1�ǜ�@������U+�ђ�$7������f������$A��)�g�����_��\%D[��y1g	�5��6��l���T��n�`�М�D���I*m�-�t<���!�s��]�2��*�;�W\dC�=88����¢u���ٻw��yi��a�)��'����r�1���y�Ø����t6C|@��_�]�P��q)�"��J�.dwu��|�2��P��C=4::N|��K/A,�����(�-d�	'��t��0-��8�e�X�TOt:#%4dV���grr����/����U<�̴�!�Gz��N��:T��� J&X�]o%&�����&/-0|"��U�a�R��7@��1x:�SLJfy'��Δ):b��_�8�����E���{��H2:ɩ�!�U���d�s�h(<G3~BC�k6mڴf��Ob;����z��g����H�̱5=���Ƿ::���j�������C�*�;n�������:.M���7n܈�y�;�q���Mw�܉)�Q��)5�#������Uf@�}�h�0�L�K>�R,6��M�H ����X�j~�^MQ�3	�A��n9�a9'.8��U��cK�.�򗿌��C�ju�A*In>F���5��I�z�˸L�Ν�j��C���=I�.q�BΆ���g�ҍ�q�7఼����ooo}��W���ʻ�������Pf��SNq㊊�4Թl��Ho�r�A�t҉�r{*�U=���i�t�r���Q�^��D;�-��ҥK���YO���mਙ�%�H=���n�-�JC�������]�(�ܨ�SB�BLj����26���>�P���JrR�
���������'�x��c�I� &��,\�5t�F�آ{��y�X\b_��b"����,	�6�AI� !1ag܆�4��ţD{J��m>17jM�}�9�GK�fk'#C�j�7�5�8������ɣ�F&�߆4q:���Mw�
�1�hdj���ډ2J�h���?������a�}��􂫽;M���M8��w��<���'�Ğ$ �@���>C�SS���"7煤�w�����q����n:��p�XF��#� �� d�u��e3�p���������^����G�X�~�&�%2��D��k/K.�]_�{�	Xh4��v��ؒ��aV�h_��m�e�9��1�A�s��@�3���}�S��%�cѮ)�H%�
'��OL��T�:qR��N�4(Lsi/x��F?���Lp�����4��ǁ]�<��m-�]��'e��shj�}�+��x&��^`C<L}�-��� kpqww7.���/,ӣ�"0�#��a6�c�+ųGi;̄�ĳ�GOS���Д�S3�3x�g�Q+��rnn�����JJ��r����<��O�׿}��6l����������޽��$,��jW]y�G	�:�3�8��:��q�i�&_��3�6t�=�����B�`�&oo/d�M��_�w�����z�,#S�{SS��e�2y�OD���8Z�I���7�P�&���j2�4l��sO>�$��J�@������X���d�P>��tP�'JA�PH7��)mm�����i���8>vw-��N:�E@P�lQp�!�0��Ͷl�2R�Aj ������P*�>����T����w}����@<��Cvkco��O~�\�
Ĩ8�"G�$�F�4̖=lx�2���Ró��e�	�JR��UI�[���e	��j�D0�c��oǃ��<=�L�~ƭ�Ç���uժ5o�����6�iC���Mug�7n����|���o�}�zz��q���p����������~P��B����;��8�T�K�����1� [@� �Jc�b�nHd�o߾j�*���K{_ZZ�������ɰ�d��M�%��,늘��ϧi��f�{�GjL3 ]�&~�$A��})%��T] ����=�͹rYv5� KIk{�EV0���o^�z5��݉��*1�U�=��Ïb7�[<n4̲��>�G,�"C�V��[�!,����m�-���j�	&��	�l�;�C�9��6�~��o���3�d5��4@n��ۂ��ú&��fPX��J��B���$z��<�I��xkh��s�9}<�Y�ӓt.$�2]�)CZngϚk�G�l6+m���P(a���뮻�����*ݶm+$�QG�7���ŋ>��c�c���t�����~��ga�?��҃k������	M�H-��]\�b%}��<��|���J==�a��l۶����n�j���z:��#>�|�K_�13��1�n�i�I`�ߠ����u�_���(��9b�=����F��Z�u��\���W˟Lxlg����ΔrR��O�%`c��w�b��o4�$^�'B��O?@-�z��S�E�X����3���'S���j�:��]��ٞ��f�<��<���O,6[Ӱ���:C*HLj�%��C��Hp�G&�O�H���W�/.`ȣ���iӖo~��!�x�l٢yH1��EW��U�#rҐe%0�9I�l�+���u�<�ՠ�ȀqO6T-Cs�K�Xq	-U��������zhl|��^vfz����}��݅ga��,jf���������<�93��Z���4�d��T��Vk#����� �K
 e�\��}�{��p�#�8�3�9� 0B��c��FD!<��P%p�3�Q>dŀ���*/2T�<3f��bs��4�glC:���LO希Q7!GH��oց��fŅ��+f�hpp{	wf��iU6�c�n�[�Cf1)gݺu�_�I�����j�x�w�qx��^|�E��WO��Ћ�du�
b��|fP�1́��W�r���<�܋Xz<���h�O=��JQbtM��g�1�
�-����"�YYɈޚd�bgR�ӳ��\h|���AL�a����W���+k�x���i&�*<1@��wr�0�
�$������+�E�`<*w�D]y�x/lu���K�D�o���Y��.�Ca�m޼�4/��B�z꩷���	n�W�4��W���{�seߓ�8��h��Lŷ���>���駟���T��[<0h�Dԩ���� �������5}2�=�H T!H˥�D�pAQ�U���
�WDT������O)���d2����){��Z����L�����af��������ޥ����!�I�JG�
������)y�y���O�o���Wp%�ѹ�{衇R 66���477Wk?uL���˕ٟ|I��ҳK�Kan՝w�ə����J\v�q��,744�3�Y5��o�2�ؠ�)�Y���Ej)AV���M(�+'�x�ҥ�.zgS{hS80�Ю���c:m�xx1aZ�Z���S2�c���;l��F�;z�\������1)1N��1���'^����09� �3a�X�I�pЇ&�0�
a,�ͪ� ���y��(۽{�o�[*���&�c .WUU�~��������)�����i +��裿������M��!i���aE���f�j�5J�:3yL���������/yٲ�J��t���-y���?�8��g{}�q9
�j�P�7n��T��3�8RI��J�B���@����\ĢJI�W2
��@�`ݺC�G�����%>,.�OJ �*Z�#W#�)-+�!}��Ba?a�w���O�X��|=?�|���
��ם�O&E�a@*�I�E�C=*���
�!3����,p��k����C��Q���H���5kȻ��Λ7o����c/9ƭ�M*�L�Kf�[gc<���v�1��N��a֋��Z�(_:�Hh�%9L}�=|qW���������/�큋��}C���Ѧ��r�:Z�ބ]��
5v���s�=���\r�a�-���������đ�=�? ١�l_��$8��vxͷ�~7ill�Y}��'�<��C�K�n;�7W��L���u��E&����Z�ijŨk��8�S�MW3- �p*�r�0�h�>Z�6JX���#�6`X�nr�ПǴt&�����G��,2�Sୁ� ���a����;����A� �H�{�W�LF�2xf�s��P���L�3��;מּ�o��6����#���ú:;4#�FK~0;�zaqIZ#M9����v�����'�3œ�K�׬]�ы/�H}�T�A�U�!Z�d�*�#`�@�@��D���i?_[]���o�/"4��\2�1 ���~e]*L������w�x�q�$|�Z700V�D]���7�q��g���#�%E;���3�]w�u�s۷m�Gm˖-�B�&M�b嵈�8���G?��	'��h�
��	l����`�Z%�������b�Ms�� C����$HW��,�(s@)s��h�1w�F���e�.�c؄�Oa9�]�U�S�����>g�>��믿΢cBsL N7�P>���)S }����K�Q�^k)�aMMWs���D�u�ݻ�`G�}��Lcg�4�BZFQ_8n!'6%�jh��,uK&Q�J4�
&9���x�-pcN!�U�)CZ�7=����1�=-�rLh�꼸��ƭ�W�;f�w�]�u�ٷ�L9Th�׬���<=2�;;���k׮��c�`��^���	�7��%�^$�U�~���O=���C�k�Ο?w��C`^|Ʌx��g�y��ϑ#GiVCPS3��0b�6Bw��iL�$u`8�%%e<N���f%�a���v�7���B��݀��SPUU!�ʒ=���^2�C���Mx`R�]�8j��w��\> �}��a���.*I�)Y,�m���I�%wٴqˆ�6Y�s=t=��0�c��͘��9<;Gw2חw�vIO��>ԔPј��]q�S����ӫb��9���q����M2�%���1^YK	 �AiX
@p�2HF֚I
Z���0�X׋cj<1,{&���^d��޽-,����tC\y�8����@�]�����O���LNh����rl�&5bc!4T�o���PD���z��"Ε*4Q�Bޣ�X��������'9�)��U�">C�6���
ֈ�t������A�M�6�=���\s�q��@����!�
��AI���8社t4u����󩧞��,�7#�����r�?����=����;�~��l5C�%^A�xR��6���,- �:���	���&�ivE����ube��v���1F��(�u*�S(!�A�6:x�~��Qr2�ԪÒ�֘�W<{r�sH���'�~�QlV�DB�⋐��
�ƌ���������O��X�[G}ب0.�ߍ�iWُ?�k
��� .�ꪫ�3�]VUW�I�kL%S�f�R1:�@*ƀ���m ���om�ӄ�c�ӦM�&�*�ꗿd����WY�~��?��Z�|��_�]>v���
V&����������ꫯ>��s���BK�E:�Jg�j���2ܥ��S�M*���ɓ��D���f�:ꨣ0	�W�t�JV e��W��&N���ư~��N8��k�]�r�TˎIY�ó���zCI�5D�%�"=L�����T0���E���iG`��:�2"U ��\��p��������i�(�);J�����v�"J�K�p)��Rl�Y��N�2��U�<��~466��+r�����K꺮��q�'�x"�pq����������44����0���Dx�J:��b���2ꁎ�ߊ�D?�)aQ�c�b2F�:h|;4��0�b$���&v��v����Di�ȸ�)G�壶K��q��m-C��BӖ4���9����ժ$udB�cx�/qO��"e&E�Um2Z���݂�Y����];�j'�tҗ���V|�p�����zJXM�/�>��x���X�6��w��� و��t�e�s0X�M��O�'��Iv	����s�:�,l����f��H���jdQpL�,�\eq@����͠g�`0t��R�w�,d�<M����!�Ѷm۶n�JT�d�@fx]k�[u"�:x0���o!Z��&3�M}�$R�1���RwZ�T%�i��'���~ h���'d��<Q�F��r2�E-�}�V-��ǖ��_(�yJ�@_��`wK������h3�m�Js\�l=�x(6�r�zL��Acc9�?�����Z�5�xl���z,C'tb�������[�➖��O	!e�	�h��,�!��4�衃3�-��.p���8�e)��(oimK���`6��Jl��;����[�{�9|�	=M�:d͑Щ����.)-�$�ܩ~A<�F���O�] Co�馟��g��z�+JK�D{�B�0GS�`�І6���/��7^��j��;�)�.=���?�����R���>^f6D�#��;/}�3)ӹ�a_--����ɧxb�'�5j8Y;�W�q�B����C��&�FAeA��s?#%�7	��(� ��?-�+�� ��t���C+y��� Q�/�XUUM�[��#$b���S�E����կ~Ub�[ؒw[�x�e˨��:a��u���֍M�:q�D��j�vء���}�YEY9�i<�aOCJ�0K4R�fpV���T�17�ʃB_��{���_�u��T��=�
��?E*��x�G~������Z�k֬�Z���>� Ks�W/�&��i��wvw��>���}�sP) �r�$�~����:rϞ��gx*���1c��r�~���k�.<�POk�a}I�s�ȹs�'�x��w�ykZZ\B ���$O�t�D=H�뮻��O&%g���M�gP�C�8r�ΝMMM���0��	�}�n�/��Ϝ����5X�K�.e�O�����CK�]NH�{zj���.q=��K/����!��Ű/����� ,�c\��)5��B"X���f1b�2��WU��)p��!�ͣ0���ݻ%5�
�"Nl��`jx��F��Dⷶv�@ϓno0�$FX��8�yn!"Ŵi O���Y�;4DĎN��?o�9���к���y��2 ���7�cN,Rf����e�4և�5��ߎ*���Wq��>*�
s��%M[B;*���\���ѱ�p�ϟ�;�[��o��0�����{�
��(-��FurD�瞷�}���|�8)�fǖ�U�Ɔ��`���M5����C>w8V��#pj`M�P�T~��S״���aU>�tègwh����]�0C�Lt�̓�,;���>��p��5���~h��ŧ�*VGIj�?[\�ڴi�!ֶ�iӧ`r4�7��x<0��?� b��[�`Ts�}O��S꘴H	����K���y��rq��<4Ծ�� ���.�o��K�vN�K��!	XW��⴯]�X
���čP�'r}a����Z?Jސ�D5S� T��Α�[L6b:64Ӓ%K0���^�ě7o~��^y�L1�y��Rj������c����!-�!�i"0��y��7�����Q�m�{Ə��Cͯ$�+eH��F97�W�7`��m�[mݶ��>�hC�}A�g���y=�.��ޝt�1���,�x1��榦���V�������u`1k��H�O>�L�=�X� �L�f�<���UL����s�&�z�0��G���:�/)1���H%;�
�+A?�;�������䦇Oe7�2E��ݩk]h`5Ϫc�q���zz��� �p1^����dSg�0N&�p	��8��ĖF��I^O�v�ԩSC���j�B������I�3C+����z�f!mo���u�֕i���棎>��;� 8kjj>|؎;��b�pVZR:g��P��0* r�o]�h̫��{0wP�0���(�v�G�>�(���Xaԡ�e^���z�o��u�����~i垀-4}�t��\��j���ihh�qO^=�XJ��D)+Lxǡ���e����=aRZa��`ca ���
�K/�7o�_�7��+�@��0�m-�X�mۥ��L��?XDvX�C���U{��'O8�ѣG:�M��������a�elQݟՍ�Y�!�b6�Z�����a757Տ���b'��I��m ��z�-��^
o�������@�1I�F�`vp���@���,A`��ȑ�T!������6n��#L�E<餓�7���m��r���Q#G���޸O>�"���Ѯ�$/I^��*+K�Yێ���0��qjX?���㬺Z2�h��"��qT�ħ�����i�lQ�!���h�k �	oQy� �@��M��@*ŵc⌴�쟸?mb+��ޝ���3����C$4m��3�B��	�;�%#�u���'w�BX�g�}�ؖ-[N>��}�k�n�<5Q�zd󊿩��X�e��Hg�ԉ����q�����Q\�Ŷ+����NfE?C�ĺcY����//Z����݅$Xċ�Wy*M��Z�cx`�.�3�9�k�7kG���F�4R�+n�"Vo�������������_�iDjL���W_=s�tu�a���`��Tet i�Y�N����L�u��'~N$mZ�;�K7t*��Qʤ�D�4��k��#����!�f��x�e��1#G���e�����,7UWT��3�L�gA(�{���g�yfӦMM�����\cd���J��Ξ�⁤�O|ɼ%�H	�ƚnL#%��U�̎�j � ��h���nQq*t<�_/dE�Q�(ɇz�D��1k箝g�}6���,����I+t½���ښ�'�N�� �5E �'
�l�t���:�-pT�����ցF�����/̞=��z��98� �סf֯�����I>?a�x��El���9�n8�Yл��MX���D��a��!��jl	�m�Ƞa��:�(�Va� 瓕����+VzL9-0�n�Cl+NR��(�\QdH����M���$/`�԰a5x3��h7�L����
���<yb{{'c4�w�Nh�qP���QG�M�����{����AXb���;�3��ꪮ����JJ�~��;^}�U,Ǩѣ���M���o�<��>�x,]�l{BFچ��cs�18�Xz�cL�/�����BwE��V���8q"�_��F�%�r�̙3M����� 5 �z��h���X
S���J*+��u�.���iӦQL`�A,3_�F;�:��{���p�1CqJ�F(���~�}fI��1^�1u��rx���q10+� v5N:��{����(����@
A����/X� 7��6Ζ}E�"���,��_x��_��_�-�nX���U@�����:��ք�����z*f���MM-�R*++0Qo��&C�t�	Sn"j��g�E�`������I��JM�d�}J��`eu�t�5Z;+t+�� �3�c1`�L&��o$��^�=�"/4����0��g�粫)�]Ψn6'��0pJK����p��G���TWӠIY]�����vZ���v7�]T0�`�-q坌����`�[v��d�Y�L+�G!�~�z�3��Ī(sh	���8��]C�ĚA�k��(=��)`�GO�4y�SN9� ���#�����ak9�'�V��w��_,\`+c �I�U^�n�ԩ7�Xq�+���f�{�B�{{��aFo�c����j�Y�f�{g�M�����.���)bhkxd�N�D*>����\�_1p3��Bwh�3��:C��w�"[|�0]ȿ���n�c����tG{wu��	�����ۍ�:d��\6��l9���8$$2��S�;����$C���y�"�{ܱ��?�	ϗ�|*�t�M�7����Ȁ�g�r@� l?M<goQ�$ı&�x%����С�a#x�b�L[/Ҳ4
U�G}�id�%w�W>���~"�Q8r�(� z_�ﮝ;�4�$Ԧ�G�E~BC6³���+�ż)A'h����u#R��r�;*N�Y�d���Z��?eʔ\>��n�:\?fT��w��ð���+*+1{�U�a�KҞf�� �W�z���	pt�Q&�Oc;r*IR_gGǻ����U�?�<���O?}����N`s���z����ۍ���q*�O����N8�[n�5ku��P5�}��G��+��tk�,~G�Oiwbu�m:�,;3�\���7�[�ӄ9�j� Z���N6E��{q?����*�c�v :�=��#���a�^�.�t:I�)-��"�3I�HZ)m6��a��vx~eɒ%�/w�u[K�Bi)�`16,͒#� ��z�~���>�7���M7) �����O9�d��0�Gx�p��`-�ܹs.�q@ف����O?e'�I�H�z櫲i)�m�0/��R�f����}��?�q͚58���,�����	_�����WU��c�p�c�8�{�6k�L����@�U*T�x�!��..Q۬��o�����T�>�S��Q�^�'O�
��X�|y��q���_����o��b�!��۷o�w����`����K���raEB����k~/����r�!�����L&��8f
����(���`0̑¹khh H�����R3�J6l؂�h
�4��h�f��)pE65�BAbx�k����Ƙ�-[v��b/���`}��M���d�R>��'�~��0R�X$>@�?��qC�}`�'��f�:�� ���U�ԅm���[�
�!'���h�?�]��H�m��f�~FZ��M��B7�`p�3�L�r��s�E�N��/�x�t{����%�J�ƌ�Xk; ���[-��EE�jhՆ;=�����2ϳipn�v��Z:>�a�h��s�QGA O�~��K����]UU�Y��sc�Pqp��}��Է��u��g�x�e�Cp�����R�Ӗ9���8PT萙�+�m<c�d��C�	֑e�wt>��Vu�=gv~��Qc�O'�-̍}�%8�T�j�{L��;��ؾj��}���ؐ��qƅ_&��t7��]w��&������Y�Ү���
AlA>i��z��DrC����Ɖ5��_zC|F������ͣ�H%��׳}�6���S&�
�e�e�xno�0��+lP-�A��
	�����Pt��������������{iu�1��=A�V~�QnUWQ)2�ӧb�GE@/1���ٻ�b&;O>t��
c1��n�4��u�cjQva?t~�֪�~�ኲr�$@(+��
0��;��3�<zB�-��n��jI��)}��ןy�۷k�f>[�;S÷����5��+�/�9��'}�Qr\�����b�5�WJ��8󬳾��oΙ3���{���A���`r�=S���r[�ɐ4�$� *c�{+9u�Js~�B=�?B���%�����&_[�U����8]5�i9��R�+ɜd�8Q�l�Mh+	����q�v$�Tk
_`l?܊
�#p+� �?ϟ?��bU���������SXK+����#���/~1u��}�����m�+W�tܠ@�K�܊�|��/f.<,W�<`��^{�W���U���v�tR
E[)�׸�����H�rW3=[\w@C��]t��Κ>}�#f�6���ꪓN:V;����o?�����_6o���NC�m
�����1����D���ڈ=��n���.�I�������Xh���������;nٸi��+.��++V� 56��ɝw�s�=EZ�Z^R>�ͱ�d붭P'xt1�@�]�zu�� ao��%�e�]v�m��iu&M�x񡘐[o�c ��e�|B4ٰa�GFo�
����vܓ�M�;:"ۣ�������Z�0�r�����)�N��S�$cmKp���QÀ��x6���۱c�?`hMM���jgB���&��I���c��ݡ��u�}���\�"��ө4iS�'�,����E�E���9I-]���;��/��a�+k�e��޾n�4a�uCb�/���;＃��5R���w�1�|�k_�9R�T�/o�[BI+���5�/X d�A����j�~��ݘ_��Ӧ�:�Q����L�-E+S�)	��.�<w�k��b�O!(�u�4R$R3&�>[__w�%�@# ������
��*vV���x�l�߆w�&I�[[�2^MMu1���L�2~��_��9���$Th /O+��t5P38���^jĈa���Q��[%��|z>��Ϻ��X�����}�8Dۏ�L�U�Y���H�v/���E�� �9��TT�������O H�ɨv,����_���K�1_|#��Ί�l���&�"��T��FbO-���`O�?�Ӿ)@��t�1;V���{�8�0�-z:a"~��JL�/���e5Yx��{ҥ��2M���,s�i��He67���e�^q�m��\�=)}¡���U�5n��9&]�izLxdN���t��ۓ�~�Tq��*�a�yְg�8�$3e�ˉ�$�Q�KQ,���(����'���K�?v6��R���7w��ٳ���+a�WT�f��H�YO����6y�i����ᆕ�ӟ~������1����E�ܭ�#G�"3�0����X�V�	}�
J�����������9s ���޸����7gz5	M8��6���د��H�3�F���I�ț��Y�u8{��2���}�L�W��JW��>�"��ț���c�1�	蚒�S.e�鏤{�P�L��O|ϪX�����݄�XD\��K/�}�� @�#����Q�"��K��͛7�����#���?���8i�������}���9��<���M�<�S�
,֭[�׿���S>O*�y��1!H������
bzGXր�̙��lʔ)��[1qO���u�5X��'֏s�y���/��G�a�M����A��@��q�I[��^��"hRҋ�%�{�H"u[4cN�p�!r,0�g�}6i�Ĳ��gl�;����@ �4y,).Q��h��|��?�����L�ԕ�_q���� ɿ����0.�l�gyC��FZIˮ��i�������n�B�@�9y�!�������G�i�
d\�e1�4�1���|f4�Z��{�Y�F���C�/�۶mî�9c��ŋ!i(�1��?�>�U�\Ĕ�^���>�D��ѹ"b��F!{F��k9����d�ӑ,Jd�����T�Ir��ב��;�c�+1
�:<,��^��JI�|ꩧ^y��e�kz�ĉ������:�BC�As70�e|)�k�Biu�Ex�ϵ0+��mf%vN�l��Bm�*��O�n�V�{����X��!�@ϖ�?��'�Eǈy_��$�@�}YN����� ����3):�������Ǌ�rmN�_��fI)�ϙ6m1�ĉ�١g��j�Gm���-�L�ɩs!W������ ��8s��-�r�����\C�mћ��\�@eeiOw�g_�ɇ��y�x�L;�s`�Y�αY���YC ���9Rt_쀿��J�Z�7q`j����5E \/*V'%w��!E�Q��Ut��e�����rE����q�*��K�����~Zi�d��*O#�RG�؈�v�0�����o~��ol߾��ڵk)h lb8����ٍ�������J:�*G*���M�+K�L�Z�Nѳ3+0�-�	!��&�G$n�x��/lݼex�0�9�frg�}�M7}wΜC��ʬ^�������YH%x7lkL�ԩS�֍��׮:��3��]�v�+#i���VU5cf�5u�n�-ɟ8Q��x�ݻwK�e_Mm�ܹsΎ;�8���+pf(�B�iE�È0�6�-樢�p�����X�#j1m��=�<��a� �4�5����$�Юf޴l"�fx��������sNRV�[�w����#0ԿҁF�&�%)�@��R�lݺ[K��kbup�׿�u �vI�SW��~�zN8v�7�x饗B9��ת��Չ"h�'����o�VYU�AyE�U�p+�	q�6m�t�M7���`j�jA1�R�������[O=��	&�0��`*Emɍ��-X�:a�8,��#��19x�1c�3��--���'�|�)�����_Z
X%
��%�///����p4Ӕn�Lv�7̢,R#�enC�W��2	���G�B Wց��V�X��__e٧�b����tQ�FUS�&�v�b�u�0����:���ŝ�Z�I����2���^�~]���Mݟ�QL~ FIDD-Y��ؑ9X�-[����"������&�C�\��/r��O�?�80(�O�E0�|�7̝;k��7J≪�0�--�d��De�獓�� A�5T�,�c�U���A�3��J���qx"p�!����۴�p��5K�.֌숷�m�p��c�M^}��w�}#��>c[!R�q��	�%�ў�ٴT,��WӵEW�HV�LB�՚V�����^|�n�,0�$3�U�c���2��a5��X���..�W���g�N��V�Y��2�YpB��@l��zN���B�������Hx	��%���=5�qe�������	Y��JX�j�NM�,��b�\G;��<�هE��w n��u�.3�9�1d2=�����7߼����0�}����v���/�~��tI%Z�c�8"��f?�us���P�NTT������J�@f�;��G����qN�84����{�ߧ�ʲvqcm޼yɒ%$��V�醋=��D�F�}���O�`3KL��>�	����of̘
9�����	�"�dmm@?w�y'�=�?�pv`{A�1�Ji��Ps�R��&��={�.��ތ���/�8��Z{�)L)�E��ȋ�2��c,I;#�1r���tlG�L�����~��k����hCe����S @��4EX��"�e�&t�-7��կ~����<�����P�-e9�X*A{.��5��	4G�N	ҵ��b=��#��̛'ŀ--����%�5_�Q	E?�D�Ոg��P��:�ʪ������\4^d�Ү�̺U�MyN/D��I^2�:��(��KF�g�X�J�)U�����
���1���$�(�6�t�p�)�N2�\m����ip�5ˤ��5 4Xٛo�����m���,�x�k� ndv��W�ܹ[;�{����1�M���Qb��� NT8��$Swt`�U�j4���d� �z�j��e˖=����G��J����h��Hߔ��������`���]��v 8þ�£2��z�ub���ݤ�$AL���������M25��]G%M�G;��.E��]rH��n;�|UUWqb555�T�/�������=
�Ly�H�0u���d
��.�=U���B�)�|��92�J��s���--�(��*���\��K/1	��i�����"J�P^�7�4�'�
��\:��˶�6j}@76x�>���|�r�TGiq::z0Zf��Zh��v���m�0��Y8B�;��q&�g��yl�B�K�����_�A���بC/��Б4,���]&�(]����SO͟?'&LW�����Q��J�<R�G�/a�`+��Kn-5,19Q���>�����՚Rt�8�K���,��͎�ߵ:���yǄ2->�*�b��j�д����Ժ��g���}�I���I�S��r��&�L�;M�l6G�D
F���@�����i3I�9��J/�Xk�!�4�}�4��cz�$��a�DB�S���[�z/B1jj�G-��+�>Ȟr�i�i�z���3!<ņ�Hə.ĝy���Ɯ��AigFr�a��?=��|��gE������x��1�3f̀�Ȉ�8���/��B���R=���a/%�}-�t��3��,�E�L��n �D�x~���H�Vv�������g3cNa��|�c��;D���%����D��F/H��U��@�9l�꤉��M�h��K�˼�����b��B"��䄹��l���u���;i���}��k#{���M'�;�T�������۷�I��UH8\��Lskˀ��)�(������d"�:����T2ᦺz�<��U	�������b�,�t�>���)��D�??�N��TPV&B��CJ��}����S��D���O�������㩮��ܴe3�����_��1T(l�E��7��uc��=g��Ys O��8��S���Z[;������J2��gK�$�����ַnR�9���ۻ��p[�^�Y!�P�5Hj ��Wq��2�)mm���;;ۃ B'k�	�tVUUU$��L.���Sh��5�eޏ'��T�7̟S?d�>͖`O�r�x�Heh�1�Ǿ�t�`6�Q[_�������C7#F���7n����۷����\�'lxO�B�i��Y�	U
ܣ�ʩ}�-��{�o�VqZ����h���?�S���/w���?�?mذ	�mƌY�U���o��NQiEk{7��`&8b�S^I����K�'����f�~�m #�w�D��}����y#G�nl���p���@N��{Wg�ȑc�� �qqkj�B������I�?Q^e�wI��($JyM����u�nشa�̙EN��B=��	�]��+޸f�&����/��;��-=����Κ�a��L�!�;;2��BT�T��S��F�X�'�6m\(�����x�[۰���"�J�Ϙ1���Oc���|�A:�f� �����U�Ǌ8��S�([��<�٭���l��E)!vI�r4Dce�/<��N�6��GhlG�Nk�r �J��IXO� X���1�B��[�n�@�jj:����Ő :�^�v�Q3
5e䷻����F{p�f��6���\~X�"��� wPA�Og	ӥ�R��)��ĉ����\P�"~+%S�p�|�Mc�~�~��)���1<�M3r���/I��7�Ox}�g�ϒ����N��Q䘴�@���X>��x�YWĄ2��?5X�^PRIz�̖�t����70X�V0��6 ���+/�eP�!FN�t�����ZV�w���(msp�uh9�1/�j}��.�b�����8J�s%�?_�����TETr���d`8ӄ��r2����5�4�����c��.�~x�v�V��h#�q�@�}�(�-�A���`��<W��c�C���IѺ@I
���̆�^KK����٬P�<������LC���B;����H|p!�
�ǹ�
����J`��X�N�EWq,e��Ac�9d{..I�3F��
AyMUO�U�<M�)W*T���Ҋ��B!Ju*�s}���T��[��	1���|����w�bа� ��6�N�-�0�9N���!�o)����j�F�m��^�3� X�lϞfL�������m'Y�����Laj ��
��]�<$����O��PC����x0�DuNER�abcn>$T�~萘5k�W\q��˷��/��s�9���M!��Bx[��_�	��ap(��5��?��O�>����Go��vF#�IuҫL�D/#�*h~�d��_�p�5�\�Do�:��K��0�-�� �:�~:��m���$��\�M�W=��-iGx��lGWi|Ie�R� ���M��!Q�>fZE��(Z�,&��uLm)OKt	5�p<	cǎ��So\D��PE���ċ㻻w����b�?����u 2Z�a��~�gB��r�qR
��)�aY�Z�����՘7�,LNWX�x^��AZ�<X*�L |E	�]ƅ���xYQeeQWWF2�R[��bKTUU�|_��kQ�0z_�Ҁ�0���q@�"�j޼yYC�J!�#����-�z���}�Y��^{
��zɒ%ж��9���q���x5�8�P���L=�C�x��z�-z�Y��?Я�^2�	��j�B�l3�(�p<+�w]�n�g�/�~>���%���X�/�Ǖ�ݽ?��qn�J�w��1���q����qd�<i��O� }+1��{(d��
�4551Q����X��q��=�ƍ��T&
��\����R,��3Wk�|�L��sp[TD.�a��P}Cq���>i����^:��S��ի�L�>}` K��:���'I��j �����n��ƹsgd���1�
�dR�o��V�汐�d�֭x��?���N���eu�c���]�|F��xXP�pC���=C����զ3��Z g�xg���b��و�0f,��UD�I��).�)�o�Smq^�1m`r��o���A�
s騡l�#g�4vx1J@9ϟ�a鯲qX���m�4Ʒc��gUܿ�Ŋ�BCMg=�	�Vˍ�x�;�n�-��[��Q:�u�����*�}�)��I�W �������*�;�����lذ�Y�r�Q�,�!E�������~_^|]�g9d�C�ϋ�;sN���/M�I����<�������'j�n��_,��q"�#�aR��~&�P�/лC	Nw�x\S�0�]�g h��/��dI?W� �˥\��.z� A HL���M��a�Ұ�S�+��GH�'�h����82v�تOf"K�����R�����#Of�O�|�W~��PKs��8������a�p�z�8�{��u�)աӤ������j'��NZ6a�?��������)�������~ڔ,�3g%��E� 2(�X��S���m����H�b�����,�g�g�5�=�!�
�q��	�(Ii���۶���cǎM*e.�u�9��8�i?A�pu`^�j����:D�Ĭ�"������C�t}��Jb���7̜9��x�����T6?__\��ȟ���-�-����GN,l�����nnn�:��_�㩪���ʲrhVG�C��q�4���J�OB�Tl��@��\v��!	�Dxf{z����a�k���0�  N�6 T89�I�Ȟp�;;� �r�:$ 
q� J�
1-���@A5�$Bخ]�V�)��ZL��O%�ᶶv`P��@+��E�$�*�
�DQ#��AJa��H�OF6��*y�`:�7��5��{�r�)��=�u�y�_���LN�Lú���>��]=]Օ©QZ^:y���[7���ǁ��)�I���y��+���ܹs?��#F���ට1� &l9�jg�tCCmd߱&o���͗%=�ۇ�ucGckABg0���ذ����#���g$�Ճ�?��ϐQ��.\��'�,^|(�'bǎ���lV2���w��իW���츉�CXb�q֯_���/?��þ��a21���s��'s)G����c�$����N�@��=΁�0��јc��NxJQjSN�k��艧���T@Xez�M�N���[���X�~�w�QT7V=�]��U�8��3�90)�`m� ��x��|�X|Ђ���}j?^��D;�Z_QTg!�gJ�;����r�� y� P(�=��]I�鯨�f�jJ��կ~�jժm۶1i�r�^xᅗ_~y2-��d���`,(^{�S^��`�X�3��"�<r:�?K��6�y��	\���A�D|@�[j�$l���X�E�WzbXB���A��(�5A(y���v�fL�s�9zIXM����@| �`�ᯐPУx7��Ao)�d�e-�⏙��#����h:
���H��1���IXF�O\2ZJDH�4���Hkw��e�]��}��'�x"^tP���?H����	�  ��IDAT� �9��t�qgc一h�h8��Ji����Γ�}}j銿����HJ��`����f�W�8���;B\'�ݲe�EvL6����Kyz��a��H��K�����`l�!��ފl�wbӧ�\ӳ���֑CM��6��]]��L �d��d�Ri]�2Ԕ8�g�����}F��@�!`�Ѹ�i[0TC-~���W	����w�}��8�$ �ǷN;������f�[�n�ͩ�\tn-0��32rd�g���۫����4��C���1����cާ��*yVp?�����"�>�l�����T�*��7,�`�� ����h��~4Nas�> UOz���0���<���zZUU���}��$b�^oYW���t�o��_���KI��Cg��;wv�����z��g�� @������>7c�;��(r'j���~�$�(//�&f�$&yϞ�'�x"���U�A2�2�����gJK��wg;��H������X/L`[[�/�ˤ/xBH��Ν;q�+;�0����Սf�ް�ڞ�~5�D�.^����Z��i�0�(��?�qE��br�0�#�#�l�p����
Aʀ��_�����S�-[6b��BBc1Æ��l�y�fX��0ܱ�����s�b���J���]�|��w޵e˖ɓ'��҇;v�z{յ�^����a~��q$1��w׮]l/�9��a>��C���n�mΜ���-#G�d�*�90�3o��p%�@d���RI3 MIB%�]�w �j�ጬ��Ɔ!q�c�z���C��&rr�~>��Xq(��w�udX��͊"�<�B�A��T:�*rx6y�`��oX�Y���x1U�x=w�Q�Lv0r��-��L�=S8h \���K��� 2����6JNh/c�v��%c� }KJ����k���+N�%�����+W�<��s������-�g��<s����31�X-�s ��B�`�2��G>�9�C���MR�8�����=*���g���g�mP��A��޽�������^Qi�%��R�i�!��(h"Am3��t�jn�s)c+�1cF}�A��Gr���k�&?�ȣ��[�����}��%%eG>�&�����Bi:��%b^3p��IO�p�b3�w ����7���/T�n̗ˉfD��h�H7����}`BPHuU�H��#�L[[[Uq5ׄ	�zz�8���|[�(M٤�����?c������1c�P5VU�^w����$�U/�>�j1_��'��1�Xk,l{{W\�H�X��[K�J[7J���2��i�Ҟ��\}�p	J���w6��>�L���C��T�=v{���Z���'��]D�h��7����
�ŝm/�T`z��1��a9T��7��裏�_P�sUX�K.��;�����5�C
ǁLf�ĉ����HpP+ut�\x�X�_|��%��q�pY�~r�����o0"��������~���'�{��9��2�Y
�8lxf������X>�~X���t������Pai'&��,��h�m��d�,�4�;�>U∯]�&����젶-�&/���|�Ǐ=�����뀓��3�`���⡗^z	�ߴ�v��Ky�gN�X�ejhh�a�:.��ȟ��|��_�h�`q�47��/���߁B��9���G+�����b�/���-�o��o#F԰; �ƍ%�w5�6hko�4y�E]�\u�wR�vu��#�@�����رc��X\雾�,l��p͟?�g��z5��j__F�3���)ej�K�@3g�X���9s����
�l���,�iӦ͞={ժU�}���E5Ă�p�h��Z1	 ����=ŬS&�Տ�[�n��{7:&��yrs����S��۶m�~�ӟ.[vBoo?���={I�<��uq �Bc υ�}��'L� ���gXЬU�����-G��D�w*g�=�!p�y�XwK�k>�I��0��=���r�39m���b�h6�ɪ�8��O��V�Co��A��>%��	���ap�n-C8�N�N0��tV�_��c����ԍ����ܸ�Ǎ��x�Y��AĄG�u���ʿ�	�%�T���x��?̲6v�f���9��s�Y�`AQq��7�,�d�)����7�K�ag�X����|fC>\n[<k���-�����r>=CϞ���kh������Z��ZO	a>s m���nw*%�y�O��1GOU��Yr���-�L4V�iO�:�B�������i'��ק�>4" dy4��C7�c����4���X�C�hΐ�G���ԦZ���M�_ۄ������՗�4г}�>�6�� ���"��D�u�I�f�y-�
�=H91��K)�TC"a�����nySM������ݱ���2O����@���LTݦ>r�r�<��l����d
\Nl2�����K��g�I�Tmg�X+�e'0=K�b/�(�$5����#��$���޽0��@�7L�Y>��D8E*&�utt�R]q)1Z�y��� O<���wߝ�ڽ��z]-��9s�7�@�m��������.%)��y���#ƿcǎ����;jΜ9PcӧO�H��'M��Q���	¿��o���
p�����T�*?�lr �>N����,;��++�3���W���~�X��潶Ǩ�[Y�Z6`�L $ ����g��؂�%�o�F�|:P��5x6vIq	��`e��]�\s͢E��3��~�b��~z�=̚c�`�`s�i�H�n�|!��[o�|�͗_~9�^3w�������#W�d.X��/|S�H��>[�ys�5ƀ?����q7�t�;�S^&�F�%%��̉��ɓ�N��mCH�T$8d����-//��+@XQ�؂V��`�\|��*R���kho@�vmZO0r` �c`Æ���!-=˵��C��b��P뇹�"��)�G`8���yT:6����Ӧ�3fL� 8�ϝr�)=�����`4�G��3�MT
̶��������ʕ+�"��0�`g��!+w��"���8��]��a�I\f1�݌�0X�~ִ�������T.6�o3�C���d���n�I��8�����&^�&)͍vXHǍ��1�V��M9�6y�f2E㬏<��/
�CINTh?�xB�ql�9KX�?e�:�t<����c�'�@g�8�?H♛�8�0���U�#��~��lj�!c���W_}��+\Mom�Pǋ������aK4��'�q�&Z�e#�΁ ��Nuf�Y���s�}��r�����$�z�����>9	eFey������Mbc|nġ���M�ޡ���6㉞�a�U�ˉ���x8�#)Y$�T�8��=8(aVMp�'����<��f���3�J*)l��r�G)	?�ˆ���F�iŪ���	~0%!X��.���0Z���,���ڗ��|�i��<$eb�+`Mʁ>���Q�s-���vj.��\l���}��Ͼ�nƭ06�C�l0��FX�I9C>LE�b��y0Ԛ)%��~��iU�ƚ�a�鵢��:�(U���*���k�GP���Б���Y��(ff`h��JL�P<	y�L�{�F���2�Zs��D��U�W ��4��o�@��3���>�(n�U|ɜ6J^�*:�㎃�ݴi�֭[���$fo��;��F��̀+�{[0��[�H�z��!�˅��Gt@XEy]>��#< &L 8kll���6|8�U<�{�{����*܍�ƪ��e���K�=�Z�_L��i�>C�H�JT�B1<ԉ��@#M��)k���J��Pc֏���1q�DF�=��I�&a	�}��ήNL?`]��7r��M�:���#�ZZ&��E��@����� �F��?��jk�b�ǌs�E�3jϞ��H�zʔ)@ ]���	���������ɃMF�9���~[Gk>�}�+_�Lfy?E���4rM�%ʫ��Dz9M���G�rwO�����:��c|%��d�Zx�2 /��l�|b���V�&q�A�������ӛ��%S5�F�e4����"R��$Q����3��L6�@Ж\�ϐ�%�<2 P���n����ޮTZ�1�g�(i��h�.%d���ի�3V������BJ�&$Æ������1�B�2�)�}E�C[�:!�z�Lr7�=��R�$x� Ԛ��K�_R��[��B��w����c��ө3�5*9�eV�Q���Ӂ��9`��ۆ���bq1����,��Xx��0�����OC �����%p��0��7\�i�@/Z<�/�9��G[M�n� �R�����M������Y�̆�ڼq��\ d�yA����KnV���"\k`��ٷ���~>�:v>��&)�S��ws���m��h3�M{j:0BfX�n�=��&}Ӈ:�Cv	gJ&�c��B<09���v5gOݲe����I)GŔ[Ӿ����/�N��{O�œ�y\Z�NG�9h���ivBEE%Q���� ��� ['̜-�f�z���rqy�\YvIU�1�C��p[����(!^�o�ҹ9J��V$c�z�J���@Ds*�(ҳ*�M��"0�\@���Aa;�J��	ã��^C�nq�mt��q�/a�c�
�n`��7�V��̓�rL;K�O���3��|5&�����l�M��J���b�5�m%�˅�j�ĉ}��^;��LN�v���,�T�Y�֓7ԣ����x�̫���0ݽ�/�$LxnE�{�I:9<���xL]�d��1@��`��֭{���31��n��6%�}�嗳��Z�@g��u��yW��3��Ӕs�,`'gs�������vst8T\��z^R�����c�2u�g��N���sQX���|�^`�5�\EQ����f�e�]_*<�#R��^�`��=��)�m�6�B{0co��&=#��H�|�J�hZx˖-[v�e��� @r�9j?�#0f��k�.<��l��zbh�Β%K ��C5�&Y��'��N۾c;ne����[J���͛�	��I��������+V|�jio��l�t4�@��;�L��8���D<��Y \\T\�0�����S,^ ��>ۄ�Ǣ�;�cGý�ދ�b�S�O4	l��ͨ�V��{5ʜ�L��t&�1|�y��u�];v���R>Py+���,"��J�ik�Ƴ���o�Y��O>��݆�}��i��!lb��ot��7_|�Ŏ�Y�Ul6L)$�s�
b����U+:({��dK���QM��-#��C/��&h� RS8TT�1FL�a�)y������Ycٵ�'�1�9j���*NM��)m[�d����6�ʰ�CN�͊�s�p!���1�����
�?	�ŁnO?Ӹ����'i�@��+�"Y�d� �I �ZԔ���!�^�ӟ�D]�y�H�1m:6�UW]��ܒ!���Rv������&G��"NF���#�%����{��j��|Fh=d\J���q{�E��^�z�'r�<ĀC�f��Ե�LS��o޷��S+��O���/42�rʊK�$�?lo﨩֜�AI�o��������G{��P�6l�ɋ�5�<���|` �\lk��<�hNt�@&�����0f����B��4��R�b�#0��20�D��Vh�S�q%[Z�������ݻ�vQIQw��iVTUүC5��d����KDR~0��:ea��7n�$?��9n3$��b�
WyX�ha".������ab������S��"m�ȘK�����%ƌ��d�0*�:�V�*�S)�]���*�C,����A�0��~M��b��r�z�Ӕ�9C,��oF��ٻ���ǎ1vy�XF��V�3���==�:�6�w�����,{]�%C	�9Z�!�8�O?���\�3j��<߰e��]�k3ٺ1���� ,��-X6l1b8��y������!��Ǌ�]ef�Q
/��/�N;)�����j�+-*%�bDLh�%�W;_\ rqYXp�JJ�� ~�K� N��(N:���˻"Y�Ki.O��"������"�H�g2����Clݶ����9j��1�b�k��Câ��M?h!6u4-=r)�`���G���W�^��?��Ņ����'L���.��466�3�8�?��?*++zzzY
��c$P�u[{ne�P5�Ql�!�ZZ�������o}��k�ř����C����hlD��������Y��� b>���	�'u�Q�:P	/4�ã�ɢ%筷����lR	��ўN�q��ٳ�P�)S'5��h�)b/M.khh�e*%�2��o��~�٠���5�5���:[j��q(�!�A>��=��� �H�w�^R�1w�A�3gb��?�|�T>"At-z��@����u��0τ��������"���c��)���,m�KOrL����U����+Ià���Q��w4h���<T�:�E��M�k*C�'�_ê �3����m��_ۨH�Ύ�X��*�x�\�䄨��F+�CŸh�R�I�Lq�KD�y����.���cj<�0��Q��o�i�Y�⚚V'Vo˃Gc�b7��)�nN��RXId�@t�>�УO?���ȑ��a;}��_����/+����^���@���+�g�d��ǅ���C;f'�(u�4�D0w�a�7��a�t�����Ή@m�^��$���-t'86G�X6�>���0���Ri��I�͘�Q���|��5�VJ5�?�n�J;��ԐD��^QAO5oM.n�&����ijIe��R��1I%��T( �������Zf`�LS�0 �<��ZGfYfz�))"���+8o��"d���A�a�@��J�	�����!�$�V�k_p�^Hr�)�@2Ef �j뵙[�XOEu�9��lJz��PțF���b14ŧ��-����w�Nx�q70 �i�h#N%������������
��3�K����i?�����<�
�Ҝɼv�W6Ȉ/
7��!��ݰ�V���� k��C�,z��j���ήi�k<�
���%�.*�,h)� ��du��{�ԆO�۷�ll����sF3]�p,�BC�Ŵc$��dբ��L>�a@赴t��ښ={��{���Dɡr�w�} ����-��G}4��#�����+0(�p��b��,#Ȭ�� b���>��uD!\D1�$�R�X��z��dԨQ��TU�uv���}3���	z�Y��� 0�o}�[���7��qF�(�]�@�,-��E]t�m��=��q���؀�����5�\�j�*�gʦȌ����h�(�=�w�-������m��}�v�����#�8`��۴�.+��i#/���w��X\\ZZ�����	O">I�9��C����9���x�@@�tKm�G&�3�<Ow��[��~ #0o�펎N�$���f�
y3s�ν��+�͛�i'��&Nd��=TH��ulii���=��H��|MJȥK�Z�T�*��27L��ŋ-Zt��?��s���:F��q�]-�"N�6�c�9��S=�P:�!\a~����*�zB[���Y��k�Yze�<�+�m?��|�L�ț�0k;9��~'�L�Ǵ�sSM�z�j���O�ɔ*%��rb��tN���kX�QX��4=Bl��3D	��*oh,�Xy�kF�i�
U�l���Wj_�m���ٿ�3��X�g� ��ӛ�ͩRy��[��Sz�X�@��9���Ĭ~iC~Q"p��|��g�=����ƩS�R�\}��7�|3׮����{��Q��������C����C� i�y;�u����[�'���I��݂?b����8�C�����`������=)��?~<E�����4I�c� �E@�R
��h�[�BU���`� �����0���B��?t���ZiN��j1`�|S>M(��F� ���AoWQ�YQ�3�o=E���Gn�J&`�fS����J��&����z� �8#2Dr��z�	��/eb%|^��M�z!�=�s�U�rEE]D9|�Ѯ�>^��]�d��J9N��ũ|w}.F���2Vp$�W&�2�)��cX�(�8�L�˧`2�X _0eV�*_+K��8����;"�D�f�y�r��%+�:�Yy>�#��j#��I��x4c*#
c�g�&ut�i���pI2!N��>�U�F�\�'��!��4�Akkט1����%���	�r�,=^���~�;LM)��ʠ�p�©S'ClRX������:R!ΰͻ���݊��1F�]f|rr�8Y������8QaE?uj[[�:�㨫
���0`�֞�P�8�O4��ܵ��#���ў�!������M7���oVCCDH�RX]2\�%K�\��;��N޸I
	�J���&�M����⋯��*��=aZa��Qs�e�a}y����w%-rF��v7������N�v뭷._�<],]n�'��|-H��使O�Ϻ;{��_���:�(�tV�Ym���y�Q��m��g���:�N8�	���bզMҾ��j�-�3�b-��C�Q�wimm�=��ƶU�}�F@PP6r�I4úQj��}��;fݺ�6n��MI�2p��&Lp%r-�Xoo�t������>�V�Ң�ɷ�j�-0��
8�á��2�qu�1�Q��Wl΍jm�ʧHt���2Т�D���,��m�����������9&%���V(Ӯ�oMߡoX*
&�?0�9V�ǣl�Ͼ�\�a_�6\͸��<�#P0�j,*rM�и��k`��Ѱ�).--!��C/քʉo�k��n �b����-}�lĒ�S�7o{��Gv�ؙ�����{�{�)������7��5W�b��0�vR������d�mˉ�<�B��ԐՌ����J�����;[K@�.����Tۯ=ʁ�Eۏ���u�Udd��t�� &۶c/c��J0q1*աG�O�g�� ��T��J����>3�CIO�ygW;0)|�=��`:Qj)3���2���1kP)}K�}�0Uq�;͗����\>jѕ3��9�)g���1��iC�eɄ�H�_QIێj�rM���_�>�%�b�~.F��.�N��Xu�nq��;jv�W���0ę5�2�$�Es�h@�P22_�\Pܬd���tjCFژ�D���?�qSSFH�$��u���6�M�/]�!�}�t����W.h�?&�6�+H�q�m�0Z���ǂ3�T9�������O��a�t٪�;v��?΀�;�}�խ[�:Z�M����k�WZR���GFYM���7o��6r��-[�p�MF;����(++�k@_B6���V�@�S�B/��U�w��n���3|��둋�%L��^��EDÒ�姸'��I��3M�]u�������U��uF��u�7��A@T��5
�B �d@���F����W��ڵw�?o!���O��+`&��%��3gΤlٹs' )�UW]1w��{�筷��S�i
��B�a��@fs��Q��4�%A?v��]R9��'N֟���e˖=��3���*FH��������\p饗b��o6/ŞI����5/�Ƣ	�lW)Ѵ��|��ѹ��Y��I~r�0$G�䘖Nq���Xv4W;$1w�,ls�1qƎ�JP图~��*9��g3M��v���Jh��+CW�A$Re��͉���.�(vL�&_Sl��f͚ŝH�.`
ӏ��A;�H�ۨLWP&�3��mq�UiFeJ�(�t[��X���h�(HU�;tP��&��>40)�qXc���kת+�����*��n	�lҋ�$L� E�$�6�A��g��=�҂��M{I��M�gQ,wQ����z��t����XV]hLY@2��R���(��'�!B�n�v���-����x���2,�p�����n�k0a��`׎�슷io�~��g{�1��	C�x�_������>��5ܳ$�d���?5]�p��(����M΁�=���0�s~�ڭ�X��2f7���,,����/Đ����φ̝u�u�H:��$�����7n�~�z5�ѳ��A�����x&C0��*"���Éw���$�=T^� ���Y�@��`�`�������)c,���n94����t9��`}����L,1��_�t�t��W���x6��Z�c��%�=.���^M!(9<�Kn-f����6�U��Âf*-����\��b} �O�(�_�-I����M4˯:�{�����R�����e��`���4bdFhz�1H��W0Ҡyݴz� P���#a4-4�� S^�2e��+3+3#2#���Y�����='nD�yd�#�����-�|��=с�%]*�Y���B8�$yE$�O<��|�{��'(�P���;w���#��5���7f�%�o�o �:�礑1i�3 �(��KrKR9�SX�Q�B���$�^x�*#�;�
����r�~�@��*���?Щ�|����Txn��7�����{�,��W���g~ZF�;�s��5�ea��h8�u����/�p�κ��n���<�������Z�����ݸqㅗ���⋔�y�.Kl�����`���ȷww���Ov{�K�F ]:Ut�r�c�p[�ĝቀO�Qc�\	�d�-tOpĦ"��!%����x����?��������[}�����ٟ����7n���w��/�>���	��?�/��O���D{a�%�R�� �����;�|�~��~�3���F�����6X�x�5]���O��O��/��իW�A��6,�>͉��-j/izXh,��_���}�=�d	������+/'��ow�*�W�Vu/$��;	ٜ>�"�a��%M��|i=|�4��c썚f/	���z=I�=+��
j��O��>��59���"˰�D2�6~�{�un��В��"MMAP`Q��w�X����	��V��riN �ćz�8Z~h�jU"��T}�ŉY�{�"�2D2!kyq�eN96:����
呷BJ--Dcf��r�r�C���3��V�U[鶵>$0�V]O�������_U��=����[K_^]=e޾)@׆��S�S���/�]8]�J�[X~�a�x��	PTGJ
����,�h���`Yk�����[o��t{�܅�/~��݃A9L�_���[�<Ju�b@�ɽjbV*�^��6k9&����[ߨ(��>��^7$��G�w�+~0�Y�ҙ�G�|z�Ok��f�R�d�� ��oܺ�39;����#^� *ˌ�gc]��NܐmQy[��3g��7e ^�"�I%k!0"	����g)f^��d���)mIU��{x�Ԯr<hXI�@�Y19���s��>h2��To�,K�.2Rwv�hc�7����.�"���*��<l8FH�#���m��[��s�0���Hn9���޽{dr�8kT��@���� �ss�kk���Z�Ԕ.gV33)�QfH�r;r��c�)���5���^�"��� �GnH$����C��+�^D���d�i*�Թ�~��;}�4�����O��O���鷾�-}_�@ڥ��E:��3�}�;���г���hl�n"����c��g~�g66�S�`��`�aY:/3�G��y�ܹ_���ǃ������ݾ}��%��<X�a�ӄ�`6�r�ܚp�qP�8"��p.���d��a�~����u �פH���i4:�KFO-���АV'� �믿��o��/�|�M8#~����Ar^�F��VW�Cz``w]ja�1<z� �������M�+l9��	-��)���u��K���������O�����?t�O}�_|!ϛ ����Q�`n���\�~:D��������.]"}f၆.��c�Y7땕��zb�5�^}�	��[NƆQ����'*��ժO�c�����f8 0r �n]od�� ��`��}H�? F��'�!���t��G2C�K�
���m�l8Ȅ�%L��Fs�CS��+"8h�ɐ��+s�|�{�;W��+�D��&���ŽFN���T�vmA@��k���O�x��ޚwT�r����y� �G	>ڎ��ausp@�}�1�����j�����ӳS�3�t<�, ��<,O4��aq<�H�����F��\Sm��x����H2U��L��p���%B%a�_<�ۿ��?��熣����eզn����-��G8�*�J�g@u�+㳐�v�����"�Iõ�lgU�6xF<y?�s��L�s��s�>ƅvؔ�FYc�$eP5An�f�w��'��s�ɛ2���ʕ+��0�2�u;��ٺh�ɲ����T5�7:�%ۗ���QT�ro�c�E����	�Y���֣��򐬹h���%�>	�~�qr�rNN������v�
�]d�rm���
ߌ*��Z&b�%?��t��R�%z�>��y֟� S9�4"4�#O�?$�ݡ��EL�/S�D1<`�I�iH�����w7��]ԉ� �	���Y�H��⏔�S��u$x��Ku�Md�'�|�I�	ҏV�PFȦ�4B�'�D�˳&/*�?�Q���	>��
���lZ��@hT���<e�+o����ׯ�Y���������EI �p@#gH�&����}��>�75��7o^}��ի��<ٱJՄJ%�Q])
l4$:�b��'VVO��Wo"Q�@r`����8��^W���,�ָ�G�'��qjz���kU��N��y#�#��&������mP3������k���>[]��:kIe�� �k#A\s�������ݲ���2�O�Z¾�@�2��:�=ŉBw��1P2����7�XZ& '��*u�|�M�q��L�q��a�ʇ�x���!46]S�����a���#�U�=�?��X�~�49�f��2oh�
�+z`đ�
g$5G�V(#���Bfga5����u��奃A�)��C�;�!�CW^\<�Im1�77SF��R����<�3P:X���i�LL4<�$ؐ��sGBB���2?Nq��"�C�ƫ8J%���:��K��N��8#�5|�����㽞-PXZ���*�B�p�T���扂����EJ��@C��$1	�"��I����Йa��S���&܄]Kץnݺ����������G}� 0B�A����\~���Hn�x�(</���t!f9,<��d�:�jЀ�x7�y̯�,
���騁|Z}艈�I�����?gf�)�2)�(���J��٩���ېri��Pˆ���V,Z��� �6=\Kx"bO�lD��^��˯yh'�M�G ��ռ�=��'�ݒ����=���s�A[02z-�T���AF]���mZ�I���+�a���޽;=5a�&){�2�9�:}��wߕ�ϓ��e1To��V��Ω��f2���^�X2��%�&#�I��t~<�s'H�a.O��|4��p��kcq�np�i�����K�.�WM�&ҖZ3`80>3��{� OR�6���<ѽ�F��8� M���/P����(t:���p�+¾`JX��P�Zx�s:�;c}��ޢ*��&�p��E*������>�e��v�vJ��V�-��q�[��0�7	k�V�+���J"zd�}"�l�H�E\/7g���{�X2�Ξ=��b�h:������>~D}_����"98Nm��q\�����[*�E���Y�6#������������3ZD/UTi��D����!���7�^|�E����hT2u�aJP(�q�&�2�;ӃL��ƀ8fn�厱��CN�\�Y��f�����T#Э�?PK8tko5��%A�	An��iP[R���$��5S���'�YJ�s�w���V�����߃!�����̀�Z_���Du�\4�><}zUП@�ŋѯ:=�;��"����������eqbA���r܄Z��;��<�U�;�����n�}��î����p�%Q!��0��-�7O�ڕph�4l�Z6�t�F��HDXi3�Y�[mu���42�#�}�H%��!�g�̭�4��'��i]�2�����h�����y�4U�hӒ�����<�i�"V�{�ufl����f$���Xy��~N4��q�.~�G� I�
��Gf�ٴ	��de���:�z^���aQ�B����s�f� ��S;0�E[���@�إt� c@[ЧG����d�G�� 
۲�v��[�-��rJ=�r_�Nݭ�U�ƀ/����04ul>��n�
��QHފ��/��\z^?�\c��W�*o�%a��:��#�9u*x�B���P�3z*��JUp*$1�/v���lǳ�
Ϻ�"s?k����Y�r�Yn��z|��>�)��Yԕv���߯�!�M$��Z�U9��u�:��ߓ���ےʝ��<�xb~fV�t����|��մ�=Jrܸ�f��'��������p4��u����w���������NE��0��H���`4ظ�bO����7�?H=��	�=~�H�Ϝ9U]n��R�}���`�˼א�c푩�\�̧�����:M����d?��S���`8��E@�y�⌑X!���y���r������d�'^�������~J�yp�>(���v�m'gN�Rg�Vvz���M�\:y��'ֵ�Ľ��%D���j��1���\ݝ&08 1У̘�Á�BW�;q� ����!�X�et���]�p��R����!���˗��8��D>F!u]�s�ySR���}r-WVNX�'&�}��/\?�&B �7o�$�Ff4`KO}��m F����?�fK�K��lM�w�\�g���5����D*���x���;��\�կs�э�O�f�8?�����6���x�ĂD�TN�;�;wF+���t�����~A�~�����ܠͿ78X>�:95S������6>||��%jeƃt�ᾑo�k�ZH]�7GR�{��>!�:]vggϜ��}+jO�����o��GU%����,y79=5=;����ٳ�<.s�)�vbi�{�{���;�������'��ِNI,3�^_ rBt{s�s��;'Nh�tYm��ݽN�x����Y��5���'5 � �ȃGϜK,q	o�L/-�|���$�Ē$����ý��WA6zp-G�A��`4��#p����4�T�2��S�w�����h��wVO�&�morp0�x�����-.v':�;{��S�*��d�LO��ᱵ�T㼷���ڽ�*�I�����'�&�w6G��ҩ���n]��f��Hp9������3��)'�Ґ4��)ԛ2#�t�{nꧩ꩕��v�nz&����Q9H��R��vv�vv(v�~�L��7���FY^�E555�,��#d�'��V&�*pC�`�V8�V܊��y&��3D�k4��Ť�z�d8��kG��1!"�>¬�'%x���]&IS �@��8�)D�#v`s���V^	�	p��V��B�M���-w�ٱ7���S:�T��\�p�̫��T����<�,-.Sk��ω	�s�<�v�����:+�6Tm�Ğ��o����\�d��:yO�'� �p�ތ(?��A��h���	�aU��Ђ����y��w�ЇTՌ̖��N�0�Y������_z���x�3��10��%�e�ٵ?��ݕ �ݥ�t�\u�����{�Wي��f�������#�36,��4K�y�5�Nϸ�$T��vE��*�<��֢��qM�<����{�t��Կ�����}�If�Q�˕���f�"������f��w�o�p�/^��?$Y�HA5^$��{�VC��Q�iBҩȒ�f��ީO�dԄN�y%4�S�� ݺuK&�����ꫯJ�b^ �����䞐�>����N`H�I�9v꼱u��(9pt�*�xԳ�SP����q1 �9��G���LfI�d���fp6�W�2"	��R���D�޽k�w���� Ƚx��ӧ�d�I�be�`�+�#A�G�#�$�%�S2/K!��:��$15"4I�'�R��k���� �Q�t�f5q! ĩ�4�/�Ձj��	B�㭁W,7zw�E��R!16*]K�Iee�T4�`��O��?(� ��O>�D�J�� wԝ;wt����k<p��/�fY�K�є
 ��j������n!�G>�5Kx�&�މ��q i��O��@��hQ3���J��L�`7i[ t�i!!]Go�N������K4���y���"�x	bZ�����P���:A�䀾	Ѯ��5>!��DL$-�[H�C��D~��t�Ǐ���ZS�A�$����CgK�"\NF#S����y��������P6|�ȆF>X�̭p�,�ǉnt@���ַcM����"L��J�П:D�e�v� {M�FB?B���$t<�?Q��%}:��1{�"sJ�8��SK��g��K��C����'ط�t�!,A6l�(��+:�f���p�΋��'>N�=fg��D~��SjϚ�Ƕ:Z�r;�6�~k��������[:�\�'f��B"����3��%,��b[�ViȐp�T��Η���VN�_����];�^t��SzJש[;��sK�Bt��fPuZ��n�k��܃��
:-�9�:M��(�i�CZ�Ƭ-Y�B{��-�K5��c/��OR�"�۷o�'��ˤh$o���o'bg3��{ｫW���N��]`q;o�^c����b��y+d�6ȼ=�Z��,����u�n����ov�<�k+�:Qz���ա�}�h�R�H��������V���),����_�-�#�����I�
�u�ĔT0�ɥ���f��<�6薿����y睑	j=~��~�lߛ'�������%B���p�@�I�h�E�� &4(Ϳ�2�{;9C���3�;(���W��@�R�����i����M�Ϝ��8i�G����""�\nKIgh�#� ����0"�{c㑾�����JD�>Q�ڳ[8N����"A 1�a}۳N�hq��z�J�Κ��t�Q;2Z;�� � ?�Τ�H+���2��qi���\<B�񠕷L[]a��m4�Ʀi�� K�
r��5Har�tA}��2̴��<Z����$��n����e����A�@�����R�C�j�@�ŗ�dlN��*T�M:V���!�OZ���B�EQ~̕#��p�R�5���� % �ˎe�S��:�&2�À&J�3���3�֖ۀ����Bc��V�.�ͣ?��8��t����/����c��m�!��\%Ҥ j�1K��J̋� �sz�ɓ��(����I\�"y�v��A��.���'Y�<�ӥa������Jyx݊��`����a�>Ky�1y�bQ��7s+c�^	��=�%�P`5�@��+6v��`�0��5Va5�M�1��2۠X��Bl�A�L�=�'k��r	q�v �	38d<)��D\!oq�W��Z��V:Q�<��Br;�g��Ѹ�9)T���9%M[y���8�Y�"i+�� �'k�؊VGΎ���M��×�M:�_����>C"�j�kVdݐ��ؤb�n���eGY���E�z�Îm}�y�ڡs�Ӵ�-��>��|��0��E-)7v'q��W^yMx�H�ΰRE�_,-�Z�7?b/]N.�)p&u���y=��9��3h,6R�o<���V�z5�#BD��t�减����mtX$�Ŭ�Z��9{����o"���N�P��'ɩr�=ڣ��:��L�Ν�0ʭ�;9���iv@�Y��K��$�Փ	8*ĒصZ댞6�/��{�	NXd����@%0AR�M���5,���!2��v�,	DB�R�)'�t�RT<���ΩS�;���;��$�mlDǆ&���v(B�5�$�:C��]:�	�A�.�iI,�ƪ��/'���=3>K��|*�����G%����	�h?�θ���_!�3���h�e{P����sFO'n��7�4P�xx:���U#��Ae���H�KIZuI/����@uA�@!�2��:X�% �ґtO�l
�iZ���û�7%G8l]]��A��R��V�� _��@���g�W,����A�b`�9JskVF1
���e��}�Z����m���1�M��&�N�.�[Jf�D.�(m���� ���k��6�C�L�b���>esIN4�^�Z��H���:����p��W����MO�-�����u�?P)y��*!�9�rW�兕.֞n"E��y�&�����F�z^���*Y;�c���
�����G���;�~{�=�ؐ�#Ò��[�#d2{���ɭhG����خ�D	�2��!E�t� �X�]��t� lWRJx����3��&B{!C��[z���%a9�9s�� =�$�Y�����,�S�4P2�'S��o�-�3�$y��W��պ��k#��hVV�u ���f^h���r�4Z6�}���%֬i�u����{񎃶��>�ٮ�s �O���q$��e��.�}�E�\Ϻ�xB@�w�y��p������j���.]�Lߔ�N�/b��F��m�Z#��d�5홏Gk{@��+�a�(���!�8�N��ٱ�vh�k���Y^!��f�d�Ûݐ��a]���U%T7+�˓S��r��g>�6+�Tbi��9r8c:���e��{�z���0-�#�ƽ���@�Bx��ص>ȣ�;���g����Y��L�4��Ɉ�:�8b������X���m���<x��ȑ��� ��O��������FJ��4c�k�LS b��q,I�㶾x����c�_)��'I�r��g`���ui����6�.�suk��H�J�R�q���ا�i���Oߤ�"A�}~�������kd�#c�'�D�Ŋ:$t�]�/�/a�{��r(��9��J����G#0�-U{:�z_�E�;�6 ^<5e��2+5	�\�yj�Q�x�p�,8vS+s))��-�9���s��E=��<�N#X5N�%��sAS\Z���׮]�=*�֥{�ux�X��m@C�t�oܸ�����{�[X�O�Ռ�x��e�H��ɓ� Zc!�h�I$���J�s\Z��D2�Yh\_Tj�5����,! {�ԩ�":Μ9%3ᑥ�޿7�k V�9���z���/�Y@���6�vU����-��^����z�Z�3����;wF�!�dDbA�ģL!�����{>�N���LU�9�H�M�b��F`� ���"X�������"x�i�,=��`"�?���¾���TH�01�h��c�$� ��h�(��H��$���9�r�4�LB��	�;N|�[��m��7��CQ�{���)ay�؛��ퟷuy �N+�f�jqb������h�y<'�N�S2���zo �:��ĤW�����)0�)oZ��~�Ad�r�UN�X9o�05u��.L�����;��C������̶b������������AwTW���էORLovn����3:3_�Ύd錩�.E`�'�/�@u��8˙>�P��Ա��<ϊN�b����<�]��������"14�9+*�2㊁w�#�#E��G�7�I�����Z��Ȼ��a���s�=��+�:g�t�ѽ`��`�)	��PȂ��7�m���Wլ��[����6"�)l2������-��7���M�&�(Ns�Bh��4Z]���G�Hfx�r"oD�D]$��ږ��{T�d�<a���LN�K�޸q�_��.�su������I��O��O����ߩ�����kkkCo�˽�d�
1���Н���VR*Dn�$r�&�}�6gO|��B�k�=k{�ga��@X��e��5�T���	��bg_�x�ɓ���x�{Q�QX⚶nK2��W<�9#	��#'Ԧ
U?�1Ƈ�FeY6�M&�g��Zf�!��|���a�3����C.�0pg{o��$تY\������"�R[~�xS�S��?Ch�lS�l�u�B8��&^ 8U`F�"<z���3gV��A��|�x��A��斴�S�g�~⑑��Q;�e���#A|�t�'�K_{
��Op���Z���kr-�;u�~�X���5)읚�6�1D�����:�%��\h�S�Nr@�\Y]]Ֆ�g/�ڵk����8��-����� �|� �o�5�X `&�o!Ͱf��R��^�g��u@��@�B$�e]�{M�%˂�\EH��`hY�1�YM���O셻��a�8P5wR;�{c7fqG�w`����Ǟ)_8�}���H",�.���tu[��'k�F������/n���B��
5��/*=%?�o�N��s�x߱N]��/�|U++�v���,sj'�I�7+OA�Z2��&�-{��fic١��1�5uZ}�90U��E+ꗷ*=���������c��w����i�І.y%f��dο��+����y��ڝ;w�^�������{_���oH9~�ߔ��ٔY&�5�EG)9�ҥK�����	�D<'���fg ����Y|����a�4��>����V3�d�gm�o������:�g�ʶ��w�)��
��lK'�u�?�yS'�`wogsK�K��|�X�|u���0�T��;6�x����_ZȲ�	�ʖ�P~�ͯݿ�>eO^[��į�t"<.4G5�-iCtS����refۥ��D��'�V@��3N.-�ˌ�f� �(�8��!�ovv ��3UV�������W�1�JLRrŨ�A�l�6W����u������_������@�����L�59kw�jXS&�5�������6��SZt� T`{��yט';�NB�
X�WT8"��B#R�U9�7��ӁZ�9�U��x}�r�u9N���X>" �v`$�^%3LC%�[���3�<0T�ɽ
�q��?������ʍ���=��$e8��e�s��t���M��seȷcdn��ٵ�T%�ð��	���x�)(	r��!#m�B������\XWWh
~O�d�A�H�4t��X��I#���x�p�˪�bixd+���dI���V�RǙ�3� d��۽���w��0=���� �Խ�4�&0�9�&�x����u�D��Q.�Y�%�Ў�d�w}�������<��
}�RB �ۡK[�Ɇt�����J_5	s]���g�k���~�-��ƾ!��[[��y�GY���#�IxbF�"�0T�8������]��Y4��@N%{#�,��VX�1-�$`ʳ.����]g`�<9)��S ��(O�����ƕK�'��'y�]����ѭn�����K/����X1��-mX�^.K�\*�0���$�xӂ�(~������^�O?��R�= O�X��cx��h�g�=o�U��b��y(���	6bH���B@��������I������_��L��/\<�/�ՏI���K�tۉy���;��h,cR�E{���)���[���E3��,D�Mt�#�v�W2XaWͅ�*|rz�vhnoV�Ӣ6Z;.��D���@�5��}�_�3g��H<@����,9"��f>1��L���8��ݎ0r��Q�3�?��M_{��ׅ�)���n^ ̶~2|%4#�<x&�`&q3�h#bU�����1,��A�I�b�����&C��»�`�qB�*�j�4b�P��i�t�o�f����)#X�HKII�t�����D����'��������������̋�o߆B���{�p�	4������s��ò�wD�&Pn��Dߑ5��Eî�'��c0��i��A��2�3Q{��M�M����:W�^������x���lC��qb+���=y����ok�uY��ٳ+���Z�y��Hb�1��#��\`)���m�ʪP�[�2��=��zd�O@<.��;�s�^a ��U ��=0�m�#��ΌJ�#�[\YY�V2B�U�1\���������-~�ȕġұ�G�?�"�����Hc"W�(u�zie�"d���.�5'��F^_����y�ÑD!r7�z"�����ml<�Zw
R ��c޻d���ʪa{�Kr@vX�'�;�ڲ�'q<��!vE�fH��������א �D3� �|�	�X�c�ؑ%G��,rD���tQN\D��@h<}��\%ӣ�<n	g,+vo��@WQUG �g�:_wx�sϸH�04W%���t��$�mal�p�Ԟ_z .���;����d����1L8�=c�xȽ�2�V�m<9ٰ���5��J��ک&!�
g�x?����.�
ߵ�߈�b�C�[z1l��E�
k�.�6�+k��(k���DZm���|���x�H��:Gf V�]e�m����u�������3�a�j�0V��l�x�V�B@��vpy�� ~X5q�C\��c�Q\\�N��H�@{߶n*b��%�k"���on���Ok�JR�YJO�92O�gE��a��E�n5�Z�h��w��?���٦0��j�g�SѾN��@�! n���0<`�)�%�<l)�hv!�
<},�u��@ɣ哋�g;y1����+˧�l>�ևc�6�Pnޅғ�Ah��A��r8	��$�20.1G�/5���s�:��|�r���0�S��;M��a$�S'��߽����=��t���`�ƕ��%+�,�?�u� A�S�--���1.%��LM�|s�>�}�b��_X������S����r"6,:���u�t�Y��)$����ӛo~��_FX�P���W�\ʢ��&	�h5Q�pK ��������Ķ�[�
����w��P��H��������<ʜϝ���׿�����ϟ��x�J@5jl ��///~��-r�q����Y�12����Y�VN�Woذ����!�O��y%id�/������B�$���}�����$�}Y)N�n�� �3<����q ���1�]__��G@�E�����5J'�ؘ@�C���@[&#���ԊG�	���w֖#�Pc�1 ��tY=wGUX	���� uk]�&���F���8loݺ���H�)P�p��l���;
����^�������������txM$#d�A��k$�@3�T�Oͭk��(%��n����h��\a����cJDQ�6 ��f�K��i���2'��KI���w�<ߕs̢�tL��� :0��gw�����I��n��*?�m���,�Z��������x��|�&?k�*�������-,�����x&n�J��l�=/9��{Q�9�de=-P�h� |x��e���s�w���a���0��T����êɢI��E*݇"�Wx��Il��z�x6-�m�ՠe�hN?��̳�+o7t�~���&��%ғ�e�/�.�����W��+���oI:��Ty;GvM�j�M��J����J�#X�a:��'���We6�z�„(雺��F3*��������>F�B�[STN~�ɳ�Z<,�
'�m�+f��S��"-Vgzfr0�o;A��,��Ͳ�j�R����lY-K2�}%_\��q$X�1�a�+W?M]���'��3��ɵ3�#cW��������O :U+�{��朗mxR)L�1M�k}��׾�����%\K���/��4����_b���#�(HQd�6k�u=Q����O�$ �Q���vv�v�1G"ĉ�s�+@�[,�+�(���TxI�13���P���w��fbh"S�N�r�
��?Lʀ�!&xU5m�joNGa&	�������<=%�dw����e"폢z|K�;��d�i����ƥ.ߞ�FOI���H�����BDN�޽�߮��ɭ�]����͕�W/���T� ���ƕ����a�G�h����0Ф�����ہ"�o��)]$�C#m,���n�;�L�"V\�m�mh=N�x.�J_�x���'pv��i��:�U����{@��7�v�f���-(�ѣME�$ ���>5ךsJ%��p�����РN�Qzg�d�Q-�\���"!�L��裏���Ѷ!��@�G}D!�իWeIk�a���ա�ʠ,�0m�d��l >��ӄ�>�l(-�*Ԥ���>��K�.ML|oSv�L"1���)Od+�@�sh�6�2F� b
���zS�ϫ������3�X��f��ֳG�ED��o���U&�]&��Y�]����H����?�w�[��̆��.!P�0�^
T� .�~NE�B���
?M��#�mlU({�ÞSWƎ��8z�70�3�#�Qa�30	�]��S�Qa.���>�E+�-ҲK��+ˆ�1�PT�\�5X������fƽ�D���Yк�'�
���)�fI�nj�;�{��am�V7�	��+���g�ջU�N��ĳ������-)�?�v� �����r�ã���0��Ų�u�_�-lU��kw��>c�8��:�8v���Q��c����d�3����dK��xU� �#65����z��Wn�����'oX�B�Y��]��so�����˓KKkw����o���'�Ρ� ��.�Nn�'�$�Y��`?���IK��6�2I���L�t���ɣ'�C��%�/_<w��������@�E2�Ʃ�22W
���`|�fx��K��H���N��q���\#%�xDJ�?n���"�
骄w��Z�g͹1�^'����qZ>uYz#��w�br��E\o�!��ԭ.3�B!���a)��#����կt]��KQ\�v�i{t�3i���<���96뤑wS��[�P�<)tNKP=��ƣH��l ��:N��P�e��#2��,h�ڗ�K�A����
�U<0�Ni�$pP��H7�4t�'�Efؔ7����,~�<���"����V���s�M� �+<�d���S���t8��6܈N�0$��z�d�56Ǚ h��I���|-//=���0��4Io���?q0�8������;\��fr_����K�[�L��lQ";��H�FAno��͸�f���y��Jљ�`4����9*�p��
l	��RHKx:���`��i�ف33iKoo���N,��ulz�ס�$��m�{�Ē����fM�t�TN��}��Q0J���3����+��<�42�O 	*=�2l��X���^�Py����3����|����_�����aA9�,`����F
�U�[�Z \&���5p�&
;3<O��R��ߓ���z��}*A~|!|EB�#oK�r���5����b�c�� :�5�^y�n��H_H8^{O�p���������c����9�e�����-�$B�0%wv�ʋ�	���A�r ��01�4�١�,;�;��%lV#I?(yY8��B
�XT4m�ٺ��⡲V(� �a��c�6����4�,�x<�UnV�����4=����!a!	�p����Q|�R5���Ck����\�@�͏?�xrf!��_N���E	B��(ɩ3�T��p0����0C��t�k�VI{��ҵ����?��'5j+E�@���o/���F�?k�>�&�p�EDl�J�(!��'����p�]g
��K �F�ym�*�4�z�{�jA
�~���Ԕ�K�'�ԓ���m֪�G�i4<�Br�-G�t_���*�Sw%`�C�t���	��؍]��#�d@O�2K�2��U������E1KLKaIZB9�PP�S����q%Кy"�=����3���W�
Z?z�x���֮]�F-d��Ud���!
k�4#�F�OD3���XR`���/�g�&�2d|z��W_�EC��I�dt�uv7R���8&J6=�Q��ҕ�����5Ix��_Z����5]���:.���!�LW���$��Ć���9��~�bQs�� sOU	w��kM�hF�r�S����+2Dx���G�̋A�BlW��9��
XL:�k�{�{"*$�;S��Pr��A����╚X�4a~'�	�&M�^����'�[�n�$����6���6`�Ik�^X�����Ch�&�z�.�a��3gV��tZ�)c�?E�Q����
]U8�w;�VZv��ēZϮ�t�l�~��&�����l6��+`�h�	�6��,����wR�	��C� ;�0��V�vΕ^�xFN���&z<���3�(*�cOL�����q��k��]1d^r)6y4�S�c�����������c6D���K/�x���JrokA̡���c��|�O,�=^��R�C��3Sc�"i�R��,\M�h+�+��)h��Vh���o]9�hҸc��Iv��t�ch���r�=)�j����vX�a�#�$󴰢U�\x�G��q ۀ�=��ypYW�@��w��R��Ő�yaG��Uԙw"�ˊ82�5b��ϲ��ʤ��6w�&gvw�ol�{�W��?��[�Y]=���$ťa̙�B�q��&���rXy)o�H�"�?�o��؀k�-�87	j���%;[�L�A	HM��
[:Z'����t��I�oq���.�&�nȃ8�ۡ�*R���ˑ�PV��gޅ*8��N
�����ЉDi��t��fu}}��T��s`��YK:���\�t)��N��f�g)6�9�^� 0Q�X[ ��P�8�ޔ���c��"x(pD�Q�{���T! ��?�h��J��*#$��:a�_gΜ�߻��}K��+++��rNB���3���L�)%H����ku=/ǈђY�Y����� � f���b�[�y��s�V��ܝ���|��d�5I�į��;˔ƃg+s�Op!��l�����Q����L销,�"�e(@(�(Ķ2��V��I�~�w��橙�Th�i�����sK?�dCAI��͎��d�E0���C�`6 ht�j�[�/c��=�MH�]���ԗ5xAmc�N:R�ٱ�u}G���A�Fi{h���Q�E'-<���9r�4���{�y+O�� ZheAQ����ά�2�=���������>�i'�M�]�����]f��y$��H�4o�� ;
e�=	�� 1����*�N���ZyQ�&Y�{	�'��(����ʪ�GF��t���D�u<դrΑ@<��='.@���H䂁<ڪ=�9�!��u��p�en{�mi����H�����Bu�1�v���pc#q��(8{�����۫h䠴 d�L�5e�=�*/�eۖx��"�[�>KfA�_`�M��g�Χ	�NVy$.�}��̴?ɒ�Yq��NM�~3��o�^���E�m���N�1�RyU�g�1����ޠ#Y�_=ȏT�և����;n��Ę˦����a���Gbs��*h#�X�)SY������d�Q[Bfu�ј�{F�5�Ȭ�54w�+*��'�{����(GFD����Ν;��������[w�Zt/	%a��ĹU�G�����[��졼L;cS�������;&��PR��^{饗 @�U;ч��K�`�H
����{�f�p�S�U��i-6.(��鑢���@'�&q.�U���U�`���;YN:"�Nu[���$��6��r"?�N����:�!�u��SF�Gɘ�L�0"����Ш�8�U6�t3O�ݱ�\�%[�ŝ�.�$4E5��d)�-�����יm�aE�7�Ή� �\)Z��;�D�X�����էP���A+|���Қa��xj/
3�㮌�UW���A�������M*�7%w>|��`~~nc�W��i��(�_�c�G�#ixn4-�.�`���F��$}-�}��՘y�[��vv��I04p��urv�^;;��������\-�B}ٚ���G�6Z�b��.�%�x`x�9)X��(!-���#ѱ0�ةOH�����`*�榷�S*��63��x����E�1ͮSg�^O���s��;�X ���7�-q���Ҩ�yN�%��$�B��"��L@�0,--xI�EЊ��1t���s�l�vro��������i��f̤7L:�nf!���e�\{|6-�pu��Z���Fe��.BT�-z��3����=���qpF���Z�����u�l��xU<{���37��.R����y��b#�7�:�����,�����2M��DE �AG.����H��y�
�͜�Z�C�S���C�A.i��V<��'ȍp��,�^y.]�/mh����۬��h�Kro	P&b1���m��ê��?�h�0��;h����HSy/��N��l��h�3k=l�Q���!ZuX��	�K5�ǴvcK/���EC���,;�i6���|�u��ރ���>�������ۿ������&[�QEvr"PZ�D�t&�`\B<V�9tU���ѧRR<���K4������_��_��W���'���/��t?'��Lۥ�1������b��5]XX~t�����
Ւ'��ͣ�H�5ȼ>\_ r�h�elw�森�4��pD�?�݉CS����-�I��D9&)�+��QI��L�s�3�s\� 9�g��̍r
أ�8l�լxnHF��ɽ����#z��C*.����!v��MO!��+��G ,s����*tSM1;�JǤB#�x4,൵5"V��p����/,<6�3��7�{�B�iK��]#9��Y�V�`���ŋ��޽��O�>���5y$@+��C���@tM��6����sW����@�o�ʕ+���}�_d��4�$��}�Q<�����̓����M�^�saaF9�.�!��Qe����KK�������	����
Ġ�dkiz5]�%�l�L�#��=��� ���Ł��SV�����f3�81O�
��9�A�gV�T{��t��
�+��I��_ג��D��L}
Y�����ζr��x�tk�M��ɓz�TG�M�dK�'c�q�P�R�VN�ڎQ1l�]x��Vk�7� ߨ�� 8��*g���$��P���0��P� E$�["�?��u��d��G>8ᐮA��A�Y+s? g�(�j�x�:��j�&�yz����B_��P���g��+'�0�t��:G`� }��=o*�_Hu�u���/�����'�jttV�ɠ1�����0�v��>?��N�6F�W��~[�p_yͦ��6���k�@2wC���L���U��Ԫi,��_*��w�ʇ�m:<mjܢ��m?�1�V����:��=�7�
�!MF��s�U��*:�r�R6��>��v�����ݪ�ek�5�?�к�?��õO���_��_y��z���s�(�Vx��K�r�eތ��ޙ[�iW��ӥ�>�7�[�u�h�A�W�;w�K_��o��o��꫈�eL��nb��Y��כ�Y
{�_���d�Ŗ�O�!��F��ȩn'�Q����2\q$��K���a^Ո��GVי[�d���&�` 4 ŏ?�X¬�	,=!z�}����t���W�.�fbc�!^��Qk�3ط���ؙ�u^~�ebg�g��' ʆd$}�� -7e��m�Q��Qqj¯\����c��h��u�r<�����2ϐ�Z��f����f^$�K	v�� rҽ�`����b����G.��nW�9�+ �K�H���/ߺu��߅����w�a���j��S���}95�u��T,K����kahH�o�S���r�u2�|XL�AC;}��Z�ڡF�#���Z��Ӆ�� D�Q��s��<xd��iP�>��)�z0��[E�i��\��ʱ'ͬg������&>c����ܫ����C�g�H31��i��ɧ�9/U�z.�y���^��O��4�o/L�²4-��CE0&z=K���t]��
04�W�G���7E�޾}�ܔ��'9��cr��Lol4Ap�$��PQ��zeDkKK'᳐U��+�!��v#�`Ҡ��Q�BHJAh����xY�Ы�#��D�������P�D�t�� �̓�:��9��Æn��y'S0$Uy�WE&bh��+0�;���>�9�t5�2ky@�ړe���V�V�˼��SD���t.huBI�LQM�� ��ܫ0ހV�s�Z~���8u7��c���p����������[�N�M��ʙ�ҫ|2��ؔqhe1�������� @v�������	��ܞS�����F-�w��;�YUqne��l5?��*o{Py�7�t�]�z�k_�=!l��_Lsh���<�Z�#��I�̊�~9ўEi]!�^�g&N�θ�I������?|mo��Ͽ�/��~�~���ےh�'���=�UÍ{wv�Co�WԐ�C:�4�fWϜ�N�w�ǣ�:�٩鬬:� q��C���T9?y�u���n��ٟ��,RK���J�͝mG��Yw�N,�nB�>^'\R^�[?LʛbC�lo��R�2t�$(�8p%��r|������T?=���v'�'{� ����&��ÃA]V��ۻ�jѡ�0�����6��S+p�>~���s��(z���:d�`���)Ձ,+���U�ǣI��!��o�K�Nz�\h�\`)��e����ʲ�����h F5?T��S}^���}��kK'�D?�7���2�4��&k^М�"�k8�n�"��I�&�4�Gׇg��3N2(�?i��R~W�M{��ի�TD�]X��RaD�)�\�?���^z��a�O ��Fe��9]�	�E�6$ǉ�Ƨ���+W˴��k��x�:��n}��r~~fm�)���+��ݷ�r�u�*4q��z�]�}E�s��'t$5Z���U��Ae�JG�儠��u�c�̤���)���mo�� �g���\��fO���)����Y�wd޼yS� �j2!3�z�}�	R��K�.����g���=����?�X+��|M��7�?�;gN��r<~�hϠ3�OlqcBP�@�_2hqjjT,+�u���:����w�M���F�n���!�W��H�!Iϥ�V�ђ�4��\�CB@3������`;`4�gL��:v���-Y"�^��ǩ�pM�����&'&�fg����U�NB�3Ć�\�&;p"�X��� ۋL��š�w�َ�R��"[>�6�f���<(�)��L�'�p�M޽���p�p�$.v4H�Y2s�C���X�����ŉǉ��H�����s��-Tg%�N���˾,��h����������=��`�1S�at�!ҕ�l�����*���D�SB��lM�~��t�S��AC�5���j��[Jp*�`��y��}��K�ՠH=�-.\������N�ٮ�V��!��(�
�ºЯR�i��Fh��ZdM`1�6n�[ܹX� h}�^C�@ⷛ���z��2��;b~��vOɼ���xX�<�h!����u~�4�[g��Ъ����k�r�-�X��4��a����_���?}r���5�-�OS|����I~n!�kon��o�ܡt� �<���$p�R����!�0��$@�t�/)�ҹIo�B*=�TrA��*�w������i>��� p_�|`�hq�M�D���*�3�12t��TJix����y�,
5��������fqr�a�ǥ���8�[^�+��b1�8���q�N=���fז�ˋ����w��}�嗹E���z�q�!�mG���vyk��D^�V�Q���>؀ݴ��s8�pa���5"Dʺ�G̕;�|遽�r΢�����Mխ�B�a8"n�ӎY�7���߀�}��P��t�J]��p�v���H�K�J��M�R@e�o�s`�#�ZJ�ނ�O�l��h��Ȥ+�?����~���ek#ه4_�Pfyc(���^__�~��!��;΢�9%!rz:yڠ�/�t �������֞�K
`�2[�r�#��ω:DSt�}5
���F��uz6�3`+��Be��z��%z.���Bۤ�e�`�e˘���G��������v��IT���p>�E��C����J`(��UR�K�1�
����#V�2!����PR;=i�Oh\^y�坝=�捳�O�Qi�wf9	o"L����X)��Қ�F�7�U�ܚmuB�ysm3�[��6+Ά�
���Ӕ6�w}��\X�6�-N��7Z�k�Ί�Ɋ8�]�xee< 㬜�w»{ٖ���w�d�������ζU{iB�t��"҇�h;J;�gBx�GB;��,��U-���׺^6Qy�H���v��(�9L���_xȘK�}cHi��,'R5%&E��<N�Հ�=�c�T�j�̽kU�1C�Abk��S����jO�;�j�H�� ������bbk��*DD5{&Xy�њ%�O���+ml}�����2�LNTT��`���~���FJ�����@2��k�����^�g���q�l)虧jfU��{�0ż d{ �cZ~�&�S\8�A�y�����M9'�#=����M��W���$a$��\��We�8��}��t� +��q���ܕ��������
u�Z._�<�ݸqt�^�@l=>}Y?���J��v)��e���(�+@RR��.]�$]����[|���g���f5�o��ĩ����W�}�����*g3�hCE��YW>e�+���R �X�����:�8���"A����N���dU�u#TQ�	��?FSDť�����X[��p��F���zmmml͂�t��)
A��L�a^���mY�0y�sb	��4P�����t��ӓ�Rhr_
��+J�~e�X��2�'T�y��j풇�������fib�=��|b8LKk1w�r�-�Dt$����8�eY�>�#���O!ᥥ����7ҁMƴ��j(�'SM?�p��s6?���ҁA+��Y�1�
�M`N:Mw�&{	|6m��Ir7���WS<�.���#�,�;2�ٜ�8�_r5m=4(��V'�u��텅9;�#pҨi,��^�"���SO�������#�&�DTh�Дe�d[I�n˝��<W�쫰*95Xĥ�F���q
�x�h��n��� �4<�"g֞ÄXC�N�-��7�Vܥ��6����C| 	@��ȏ�#vN׋'�{vk����l���y@z^��\u�Д��9��a��:7�3���Z���@���;d���N��F��ۺ>���CRe-4�,0j�a�WE�ҚjBL������z��@(F�Φ�A��7qi���������Q��/|Aj�<�[�IFT��o�P��<Jm����S[6�lk�B&�����{�Vn�!�XH#�h�+���%����`��#*�x&���`%�͌�	����&�?�"|W��i�E�����C�\�@��>8Hq[̸�����@1CN�����W�s�֭[_����IY�z��_>y����k������Zb��)���v��	�
\�yea;�uB(�
+�Cm��)�Z��ɵ;���M���I&�� p ,�O3j&�miXaj�!��}�d{�������%S��a�~+#gb������k���6i�B�h`�e��-{i����(u4]/d� jd�Ũ�Z�Ǿ����6G�����-�0	8�zc��J�)¹E�jbxڰ�^zҙ{�r�`��{)�������Zb`6���-ݱ�KE�^S��;���޹s�k�¨c- ���hju��	��!<�C�gYYY����o%ٽ�[f�D �㱃(N߿y��q�i��g�ɓM*`8���1`�oݍ�M���In�&St�.�2��RY�ԔQ�#�pO��x,Jj�����s%G����?&q4)� b��k�$���"�0��٭�r
�! �7rhnV~�!� �kg����ل5�t;�&�u�Ü)�6T�V��p����Z�so�#)B[z�̣�<O4r��ʉR9���:^G�Bt����͔x?��Jd-Z�܍ۘƀ5�"O?�W��߶?�ΧE��4f��Qr�*ˏ���yO� Iu��U{���l���_�3U��>�@��ȉ?�^xȰL8��`���6E�\�zt�!�q�����+4�Ʃ�u�ʛ�wZ���jC��}�����~ �Y�v���m� �d�jb@�O���1��3�?S�yl��g馠I�)a2/�N�e�Ϊܔ&�0/���{���ﯜ>537-���������߇ݘ�L��7����`���dE��9-�\h��5���(m�e�ci!�6�v�_1�����x���gZ���kaA��T��`�Pc�Y�1�x��@��x�1h�v��;�K�������R�H��`���V�+�t��D��D4���Stz���}�t��t�s�=g�,��O�n���`;�ESb@ ���2�#<�;ѳ�%�.��Դ��6Ma�7�;!3\H��SΕO���*giDM��%Y举���������!I���G���(�7�"M�e(�h��GW�5laԈ��=���Х��AJ%K������?��"��2K����0o�xX����ҡ5<X��q@4r��ܹs�O�� �jD�9��Xʞq�	����^��
j� f�۷�uM�P���n�@���������($i�˿J�t�d>����qVV��oL_ӳH�K��R���Bi����|���w>��C���իZh���˗��j��,��J>+�aחaK������4��"�_x뭷nܸ���^���JG��˕C���S��f����E���z�,��z��d�֖jB�v��B���nk�f���#������ضZ�<�1\��ں<�F,��z^�����0V8E�B�}i6���^#�F��Rƃ�N]�xG�݇*?w��}?V呯�k;B��G�
@3t���EZ;�B�4Sj�i���¸bi�=��q6l��}�De�A����cR�LIE+z�V�m(��G#`el	EǛb��&
N��y?��C��I=�-G`�ΧX8PDx���<gh��a���|d�����X�6H����OG�(�%���l_������9>�,<�[奕�A�tֱ,MTiykkk���	+��|Y�C�
��U;2��C�����NBĲ&���O�+�<7���Z�?4�Jl�d�����ߵk���M%N��a���y�P�% ���xD�n@&����(u�؂ȞD�@K�O\#�wN����ڜ
�C�I]��a�c��X㌽�%���Ng��%/�r���􅹅�,i��fѤ,��ș�^��D��͔�d�zop*������w��ā�%R(hZ 
)�Y$H�v"G��r�m:MQ�~N9dx#���>H6|<mlY�ϸ�F��&w�����+¦O���?�6)�����B��!��p.k �wt�d}O$'QO� ����-e.jI���
���c���l�&��m*|c�ި)(�}�3�y �@���:6���LUҖ���x������i ~j0XF ¢�F���Z/r y�{:q�=SM�>�z���i���g%�s0�a��K�'H��X]]�eR'&�i݊N$�w���o��_���z��?�x����_�7~�wW@�*�85?�s�@��=��M�
�Nؑ�;w�hgά|����/Y��N:��4�{��/����������un߾�DaMER *��$�7�nJ�6�[�\$�Q���Uok6��q}ml< �E�o�q�/�(��x2�,�W!��L!ɼ����V�����a�;����93x4p2��k��V�����5�cK�F��c��-���?!���Pz�qXA��B���I�����	?G|��2Ɔ�˄X��fa��J�!���1��{�B��C!g��Ybc���{��u+"Y�bv�j�HD��4�j�	��<�����5�#���t�6:������>Y���䵋gW�K:-��̉���-�,&pXL����4V�U@*�Y�&��溵��}��xb����%�A�F$���q��fu����}5��Y�տ*'��e�������c��ԟN7�G��Fߘ_<1�O*��w���VV���� JG�\S{2���s�{J/W�ySp��9.xS�p�������`�����6O[�k$z�:M�P����T�kU�85w�焢�F-Bv��I%���,�JP ��,-�XL�S���γn�I����F�B�+٭gѣEz��hH��<���3�R���_L���{��6���5���>ZA<�LiO7��0�bxIjX�
�X��m{N��Kk]�qV�� #�V(�3�6f��y饗�VoAD/�Ӹ� �(��?��:�a�J�\�ƻ�/'J`�����oQ[�[�*�5@߁%DH������P�SDX����tRK���ܐ�o�D'�c�r��E,�d��~�t� M�9�,�Sn��2�O?�<��:��祉�] ;��>,�n*˝�������եK���Y��'�t>��݆ NQ�-}d̈�������_��_ۧ��ēǏjuJ��ܼyS����?��O�ꀬ I�e� }���3��)[�U㘐Ȍs�oxe�������?-Zڀ|��'Y]�&��|��_��W~�����a�|rϳ}�=�&��"��*o��>��I�M8�ӄf޲�����bߖ���ؾ�H5��y
-�N�D���1���y�K�:�+8z85r�/�#'���0$F��Kv]�ٌ1rpוξVz�[�bq=W9����j5�[u��g,Ӡ�>	��s �V�/�~4���$��Vd-��ЫD#��-��q��c	���Go3��g5t������B$�H����-Ǖt��\���C+����3韉��ʭБ$�c�ӊE�*����V�1�K?�i�֪c�ꌸa����0�tV��,-=8k���v4��~СG|�7;�7 $b�uӎ�p��R��ģe-��c����c�y���<�ql<��GH�у�|MS����r�?����W+���+���l
�Y
Q�'��p�j�ΞI����K�\�|�������;�*�JuR����s�َ=���J/p�2�k��a�� a��c�� KnB�o�? ��r0Y�Խ���,�3�� �=�3���C�C�h�G�� M�gOt,)JÐn#��.T�F[O����ׯ����LQ�~�,�*��K�O��r�
�$kR9�+E�������|p�hH�`篼��҄�'VG7L�Y�`�8�
�`4��:�4��8�+�bŕ��,>T}S[���D���?I{,���ESJ��,ޱ��[Ki�t5��#ƣ-�gk��aE,[+��2���"e�U�,�p��v����(�\�,:N��D��`
I�/C��ԭ��ֈ�ki��	�a5�8H�)�'-�.u��Y�pt�UCvs�QȄ+,^��bio����4`Z!�L���X$�^ʽݮ�=s=d��43���[�~��?��#�%��N"��ot`������//_�x���d�����6O�f��:�:v�b��!X����'ٺ����o�
��k�4�����NӀ���o����?�#?�e2�9�H��9��77S�-����241	d0N>��E���#�y뛚�^M8ȞU�Ͻ�يS��y�|�+F��(
W{������j$Zw�u�|��G���kߛ�CKAnG)�q�bk�5 h���m
���PBY�|�%7��T��Uͼ�^���
pjBS�e�&i'<��+�6�j��l�{"�,<�^��޻xp	Xמ;�7���MS�|U��-s�I�$�U+�j��W��6
c�z��=y[��OV6�(p�'�p$\>����I�7��s���=h5{h�ըž�9�^�����k'��)���f�r+�-f����!�����������@Nm7�őJ�,l�ڨU$"�}��Pލ��[��T���pl<�6$�3���>���M�<�x���e�ם^�*���=y�2���n��&	��t���ղͣ2)l,�L���*%��Ý��=����gkw�L1s�h����|Q8��f?��c}��+���������|��l��z����֓���߹��ະڮ����Az_��y�{i�#��{��8��D`�ܸqCC=w�<"W:�Y}�����P �Ff��	}?z����������atęDEX:6Y=ݟ��������(���$m%�%��҃���Kr@<^`Gt���5�@�7�&�	�[�Kl���V�������_t�K�.��t�# ]{��V�DGJ6�<���9��C\5�2	vVV�J�S�θ:;���{�T���Ț)BR�5�={�w�͌�7mk`(�F*\�՜���e릨^�@-���͛������3P�#-C����^y�Eɩ�~�����*H�C�%�D���'��'h͒�8V�!>�����7�i�D�㘁Q��<dh漠��Y r�*�����z:���	�Yψ	�hD��W�pGw�b����;�co���y�y��m�g���W��$��,��e�˾��=ƀ�|7��;�����;_=@6t�iȒY�͝IY�*֞YKV�˷E��_�'#��@'"���"�x�s��=�.�ᶵ� L�r�\]���v�1!��1��p*',��k�)����Ç��^	\��PC6��D���K�&�$ӎ:|닛���n����h[k���fg� ^CH���[�O��`�v���b�������VK2f�o�_A(����X8[�{8��VO��66��������[;���FE�9S	j�y#Be�F��	� Pe:�Z3 �rq�Ӂ&('L�A���7D�%H�憏kx�V�6�UB�t�	|�i:oI��'&����@sL��yg����g1i�U�<9�eې�o#�Q_ҝ<38��ߠ;1�<E�h� H9
dfJ˝
�¤��f�>"��~隇�2�1��o1�u�y��O��+�D 3�=������iㆴ:��-�/��駍����Q�S⪐WSessړջﾋ��XN�_����U�	2G:���[�c���	E����iث�����F�"�m5S��kŦ�F�.�M3}�2W��F�^�Y�����UŲ ��.+�&YLjOb`�.���v�?s��c�۰�;E��=2[�h>S:2^��G���VV��*c��p_2`���UR��Ed*�tw��
�u?|�$폓 ����W�^��b�Ο}����/`(�� Ʃ��m�ʼ^KD���X#M��,1?-N~w�Sf_�b���Z���J���!A|m~^Fv�x��2KX��N��J���n8��W�զ�<���	�d%.a��=y2���ؖ���#�U�\�g�"l77;���]�~xVd���2�4��7nܐ���KF�Au��P�>���<t�z�jZPɀ \�pO$��6��.I����p����;ٽF��Pj�S��i�`���k׮]�p�(�S�Aj�X�Ʀ7B'���5�f���t=b���(�d����ӥݢY�������F��̇�y�`�ٛA�&d�H�w��aa����{
����@hS�����m�(���4�z�7���y$��H���%���:���V7�2M��RcK�PҌ�[�����E�����@{�Z"S]�<8�
8�='��[a=�ZF��a�{/��ʕ+'N���'L��o��C�E�&��O���ϓ
&l
�
�����^��m �ƣ/�gϞ\^^�O�:}�MԴ\E������^`�%v	��:fV��W���_5}��E�`|�t���;w����/,�xx��?Ii����Uص>��i�4N�
F�N�^��铒v��ͭ-4p�+�+�h�Iҕ�F2���=�#���el�d�	����fuh>�
$"(���it۵F[�c������Wq��o���J^h���g��Ue������1͆
	��k*���J��;���yB�(�?�߲�����c�5��gt�$)"�4���'��yx_��!).�4ܟ�ˢ�<��[#�F����]���I�#e�W�D�I���R�=�뻥Ե�[b��P}��+i�=Z�́a�FD�i/NӇ4n0~5/hb���?��)Ud�c�Q�X8��"���_X\IM�P��=/TtME Qo~x\�zY#��=ґ���k*���b�?s���3`Av�5���'�Pu�h���t��Y=�`��/��)�(�Y��n��a'����A7vG����k�I8޹{�_���($"d�l�ђ����fZֹ�f��l�������/u�������QU��3���R��$	�h&]�%�&m��7�m?6� ����f�bR���j�����DD3}���Mb��O:�7w���"I�DF �é�;K��-�i�:����v��~�2��æ�:�����+�&���`ˈӎ���\SY킔��H_�~�zZ�<CXdh\��c\k��!!��(��^ڋ�8��դ�&2l\\���+�&��K ��|�;S�-{7R�F�i�W���܁3	�O����Ի�CM���ٳih�M��Q8a�����dyt��G
ϫ�-]�� Ŭ+5Qz�Фv��ձ���A����(�<ZBeFE��j�K��!]���΢���t|f<d�^��wC"َ�b`i����Ool�h��G"���O:'��!o���??����C��Qj�O-�m;�>���D8�=��s���J�0������kn7�p%�Q�c�x��{��1���q�S4�A��l��Im`H�kz��������������G�c��W['X����u��s��*���[S�D�%n �_c�Ŏ^idN�Y��K�*8���,_̦��~�uʄҠš��}�:��55�"�XtH�y��@R���G^~j*��b��k��ۻ��$�#����Smc�:��)�B|�W�L���Z�"v�� `�f��%˘�$s�.N�k�u�	YLWO\Y���:�N�� {;;��BM��#eM�������M����j�/?v��F�Q,¨,�z䧇@qG\-@�C��l*b����lI�x],�+@]_�;?��d>�����{4�=�}�0�h���A|+|C�����6�,�����؄���~[c�/�t��`1����s��׿�Э�T�i�n&KB��j/w�R	3��dEN�*h:��V�^?���4����J�������PT��.���O�I�5�1����'i�-�!���Jc�-%�vo��ds'@��e���6�qQҍ��fF�O<ӵ���� �9eXQ���'V��W���F�-��w��8�a8�PT���Rh�� �Q샆�������b�Q���S��{Z���N Yt�'�1�M�P0�8����t�� �NG^�Ӹ���.�IdJ_�"�4Fo�_�&�\3���/)����8̃Z3^�<ֽ�����C�y�;x�[���R8�<h�<f�҇BQ��P��[7�n{b�����r*I#C�MX�q���-uYL�$}Znݺ�:Ѿ�$@��s��G�<�g���a�`a����R�2��_~Y�ݺuO�H_���?�5!$�F��V��Ow������&��@�����Ly��	M?0Է�XoG���^ͭ� �9.1���!&���
|�;��럐�j�V:e,������m�_�{CO�|��&�,�ӧO���$���Ӆ�;�Wz����bnN�l���X������By��B�.]���,}]��ʕk w� ��2�t[=��VђL{�w���OM��'�,�Y�'H,���&���Q��"'h�3b<A��q��B ��f���%�&-Os��U)d�H�IB� �ʚ0�K�0!�M�{��rgAx[[^á3�l��Y���f��ⳳ�8�6�-r1��:L��H<�="�aSՈ�y���Pf��"y�Ǘ13�)�ye�vD�J��'�U�j�46�d{�1��V�������xq��caAz.L���V�g���W�����I�Q}���z�����'OV�NW�B��>����� ֚����!���#mP�e��ʤ�?KiXi#��INlm�P����U1fǶ7a�/c�� �e����D������l���b-p�d9�+�A��k:��a��ڷ	���;�y�d�~�f�C�"Ǫj�AS�9�PL4]}�����ܲ*Va���@z�mni�}v�fh�v�l�rWۛ�A|�2*�vM?i�$\JZ>�rr���`�g�l�"��3�s�é���������D�a%�:6�R��zn���"�%F��y���4��@E�܌�T�%l���UX^g�!8H�B�A�7ul��Vl�K�q/i���'��믟�pA�zX�<'UnY�޴�C���@	�ɔ�A�SJK�Щן�.(Et��u΀~�����t��IWM\G�LE��u��g5�j�]���YH�1����;��'/#�t�s��!�nܸ���m �g�,�E��040I6^e��x7Q~�ºQ�H�pƮS���z��H�ge<'�?����ѣ�/���̙3�L�.���(S�^�yW����6�qK�����C0�a�w�W}B3M��5^P�D�\�tQ�X\\����̘q���Nz�M"�&Y���(���ؕ3��Ġ	���E��h
�X撘 �0�$�B3�%SW$ b�ߴ	���zBN�ػw7]���GFpC�#�`_@-��4S��q{��%�c/U1o! ����Ғ����WI���<VuH�2 � :�R�F�.�zJ#Ksqg����e����X��v�`�����������:!�:��jn���D��F�x��ؚ�bL�m+�P��C/B �?��ۂ���9�F1�����@�{��ӄ8G���C).R�M�ΛAlL�Hb66����10u/���z�Ef�,h;rX��]TF��,GeLT�F�kb"�1��٬�h�2E!��wmw����uj����Õ'�>4���&GǓ�P;8ؕ})�r�� ��S6r��d_�AՀ Y����`��M�ȩ�E��J�o��v^{��y$�s^� �H�;����#t4�+h�׮�,֖����o���c�(Mc3�*j�X��L�h�8����%B�����y\��Fc{ϲ�/񟅓P��RX/v-�Y�����V�-Z���^	2t�C�~ `,lonm#�������� �sff�ѣ�al�㺲89�etϺ�,�4���`k�T����#nt��/�
)�.'K �!D�������n�s�?�ؓ
#R��j�!|x�|/rȑk�����7Ѓ�����ql��O���ʾ=�����~�ρ���1z�>�|�2�������MR�4����lS]I��8�]����
��$uw�����H����t���m�{�Ď�*���H��������"����31��T��l�-p#AF�Xjak66h�����c 1Y;_�k<��:�#��@[�@�k�\ztf-����R.� �~����nVhyT���HPo���@r���7C�����ks16�C��<1�3�y�p6�H/G�Lw�
@d�I�lF��:jM��~FN��Lo�����=|2;�&+z��~�������ώFuq4��U�_z���ΐ��� N���������SB�Q.|ۢc�J����w$��Oy��B~^�����1G8X�(?o��1�&��+�����\�X�nd�n��x>�I�Xb���`H�H��5���ޓZ�?� cg33���ư�&��! ;�H�Q��WԊL�Il���B8$1��5.�A�n�	�DgR�+-oobcc�	��E�b~zҨ��>>e��)"�Uf�RU#׭v�.�-�"򵲵&i]��Ӻ�NC�"s���)&&�Lz��c"Ȓz�B(\f<��qO����i�#�#̰�݇1/��r?����Z���S�d���7�oU��|��� �C�&����,~�"��'1��ϵ� Yp�������r%�q�h�&��h/�?G���jb��/oP14@Y$u�=~�n�w�q�6���ګ===�����_��4��������)�Y�Ӵ��e��dd�u4��o��m�2Ѹ�؜���\!�dc#%wsd�D��zf�d�t#��`8@r��,���ACr�I�Lb�,��SZY�0Dh�����Xd����n�$�O��������l6q���+�����׮]��OB6^��y�+v�b&ur��}�.T�2��-<^���0�����`o��%����5�C��I��u�RI��EnaG(����Ũͬv�r~~zy90k<z�G#���W�0�N�Y�GbP�u$I��w��Ǔ���@oĄ;��Lz?��t��ݴ"��	�t�Ç�N�>���(s���P���Y�D0Tڝ,o�}�xq�!�u���^�/��=~�L3%�����JI=��w��*_�xQӢ
���:�����	�����Ý@�OXB���J����5�8n1'
c���}�����a��!j�Y������z��Ա���*G�$��t%B+��'O�03�&�H�)0<߹��Gvr���ϳ@�$@>�%x��%��==r��).jM4����[�۰�0�1Jc��0]�[���i��tq;"s��	"�05^���z��y=��tli���4���ńwwv6�خ�Z�ųH�����`�� �b�S�����j�G�:GS?���|�H@�U�y�2\SZ4����!�Hg�E6�*�\��ci04:Ws�]
�j�����a�7�J��S�'��a<��@�1VY�ӊ� �y೭w��&�!AOZ�6F�HB�����4��5�(���*6�Zݫd�V��mtM�j��B�Ȫ�u���I�a��ޕ�x�����ĉ��&s:J)��5�&���ŇX�o��>M;��iHi#U��H����m��q��2|Y�F�B�(�l ��فV-#Q�;����x�s���X��8��es0M�֜4���uD��?#n{5	F\H��o�~I���?o�����<5�	���lY��R	���܅�rb*TXY��|�!����%VZ/��p�l�ZZ����$�� 1�t�#��1@1��d���h'ŁCA�@ǃL�)��U���Y��L}�����ݚ��\�t%'�ЊM<`J��	i�Rx.��Nl��x������wa;F"� 2.m8��؏\h��6���d;U1�Q����?z���ޓ�歁���{�������+�4lж��P-,��[��Da�����c�ܵdz��U���_��W�N���ASA9Ui�5���N�,�^��g��ņT�9A��\�f��Z���&�tss�H$���j���pѹ�G��1�麒W&e��S�j� ����l_�7������?� NY�
�"!i7p��i+����B +.�,�'}��ի��i�h����������Q�E`rЩ9v��
����EX�����m��8��'����J�/��z<˴���˗u��;s�$F1�U'6�I��� JE�ͷn���ĜmD��Fy,n�r�v��q�ɾ�q�i@k��Kv9`5�+x�6�_���������ϒ�߷F����녰Ë/>��Ѳ��M���19Q�*Χ�^����b�R���F_QM�ٳg���<��<w�̃��aB��1�eaqK��c�04V�53.�l� ��Tۜ]��Vu� �=�<l�c5�a���$V ��f�0D��0_�*�Dc��4��Z�Js�J�/�:{C'�v���JcFM���"�IP�N���&���r�l�m�����#I f������&�mL���&+�����ၖ�G&���#���׾��K�mW��#������P]j�?��3|�xtLt��x������[�ni�h�7n����}H��t<�G�b���x��s��U&I����V���'�L��~J3t�g���$�jǱ0�#f�i��{V��+��[���Ķ=PT��:�rh�S{��繷ȇ�LU�X灉J� �Q&�=��qͅbL<I�RC�# ������<hE+�d�����fА�>�j/�GUQ����P�;1=��xebn����n�����vo������;S3�cS��'OV~
$j�eV�-��Vp׭����g����N	�4�`�:z�\;$[�Ζ�E����	�����֮�րA���ԒL�����h�֟�vЕi6�V�p84s�+� ��͡��2��0w�X�T�U��*M�76�k�Ao�[�%��=Y���k?��|O�l�l�D��.޽����U�>�Ɲ��t�ԝI���t>0���_�]�~]2�XY	ۺL��ً�]��W�<s8�C%��HI�=|�������GÑ��i�7��Ӫf!՝���B���������ɩcǏ���J�\���4."��>?th�t:�V�k[j$_�V<5S[߅�C�S/"��cm�Z�g�z��޽{R�Z�ҺQ!s�S�0�G�糓�����?��h�/�zIC�R���an��(}�>9t��S�/��ڵ�z�n�7��5�1�\R0�>�%@��q����n����i�x*
84-zS�j���?@��t���ǫ����Z��:����n�~��sK�Fc�������矗&x��4Z��顈x0��AO��6����x��s"��\�����F���׶���s����oJ����p~~���S�t �<b�����Z,,l���勏��{*�ϒ�S���h�%��	y�7����~���~��_~�*:up���z��<�p�.9/�V��{E��k��g��,�%-�������c��-]О����ٙyi��ـNvv�nW�'i�;�zS������ ����ie���������xjbH�j���������~��)S�ԅ�٠=�Dbb4,�����[��691U�ɸ�t]=rd~rb�>;=�Y����ؙ�Ƈ��3Ʒ��s��i�^�[�����8���f�V7ˤ591=5�e4�4��ǟ���;B�:�\O�~؜��N�+_�}���!��ł&�vm6z����+��ٱ�?����Z\�ZJ%]��N��$�v�"6��_Z	 ���A�'�6�Eϳ
a��軲F��V!q��K0�����Z ;M������͏?u?�!
O� +r��wKp�T]Bl�at<N� l��e�.�`t��ǲTe1��ãI#tX��alǂgKo� ��bL�s��l������,C�Ui�{j0��<���b� D���ABEM@�{�����	se����GZ+����I(*��L"��>�=c�[=Ǆ� �;��Sp�W�YY`Z�k�;��$�S7��R������5/a,k�MN��Kg5�9������@V�� ��#�=p�[o��c���fl'�/@]!�p�V��'�^��_D�x���w���?���)vY$^ǋ���f<~g�9�>�r&杚����|��y� ���$�RP	H�e��ڭ�Y�D�c@H��3��`�
��A�._�a�F��$Ƞ�'�"��Vt��}�����k����?����҇�`
��1H��K�� ���[$u!���6CaoHl�y!�#9"�977���������^*�z�:���(����鞮�z�@,Բ��5�χ�*�'�KZ���u�	y�Ii4*`P��9�I�-��t�n�0M|Y��W���nz)�����2�}�����w�(gK�S@ �w���ssS�	��-R[��z$���O�������R��fU��M�	�-��M?���駟�сqԌ��)��G�`I�����)�E���3gNܹ��Ӂ��
�Տ�����9&��Ɛ�����45*iS-.ܧ��!�@CEYR`AF�&_7�;�īQ�;`�v�>������6N.σ�/��(O�m$m�K=�%P['A�v�y�&��X������a�	�j_��S�y��a��	azrK�H�6�O����hDvv_����D���j�2��B`�G&O���'n޼ۛ��7���ʼ�Y"���Aȑ*ra�lf���a�!CE��|u�gv���K/���51!ؚЮ@�r�X�u�%=4Z�}�/� �T�%������L��O#=���B9��O�A��m��j_�K�.A�+��#�TSJ�3�E�CY/߭m��Ъ�VJ�Bk��<E�1&q7������OMOЯ6��$Q����DRx�h��xǉ;CD�
L.�������桅�G}��_���YS��更K���z[AQ{kv����_;i4��E�h�b[�!ș#V>c��V�!"� �<X�U�^���E,lLc�l���ox�W�=OIL8s �ީN쵅Xh�Z7��<BD8�w&�]z�R�F�!���Q8Ł��7�54Y�k�}i���:Z��E#��%����05���ʹQt���	��"mHj�����aP�8��ڵ�B���4qҔ8�}�=�^X�xGǠ
9�ۻ�\��ӝ��`A����˭JN�~zr��jP?�đj<}+g�H �6
G4A��|F��,V����6%��Uq)���6,��܄g�3���
�ic{�n�1[hM�G�{&-d�2��Ԡ �gz�NZV��N��JPw�q��ą��$�I�� `lD�$XHT�d�y ��J$Q��ۂE�P����N���O%0?&�ږ�O7�Bb� @��I*aGEl�����u>OC 7i��=й��m��5lA1	w}��dc�3ޝ]����Bl���*�z]�l�i��R�q���5O"6x�L��9�;ĳF�9���S[[�!�;�o��C���@$&-�;�СY�Xf~>�Zʆ�"��GK;�=t+��I����D�H���#ҬB�,�E����++ƃ��Z"�fQkz��Y@	��K��X|'�-�Y�b�+T:D�����E��S�臚A���/
��cK7NN�>iYY���Y�t#��Ҥ��N�:u��Pə3'ww�j=����mV>a�Ų��Ο��d�I��ܺu����'nh8�e�\F�Y���� ��(��/�>dc %���bi��B�Qr�J(c��З��)�ee�J�������5W?���F�J>�wlKY�P���,���o�ϡ������^}��P6�d��Z�-��W?��
p� �&�@М�u��m��7��'O�.)p��G����;s^�׮&C�A�.��RrП����R��^6*��:Z$�������cx4MMNyJ+�eUN�Btf{g[��
�ǒʦ��n��˝`fi�-Mn(u$�<�'s�|�wn"�<;�i9	g�B���GTz�f��=�Ȁ9�xu�o�qlӞ7�4f����Af�I� +�U��3�%m!J>9CtH2��<�Q���Fi�bZ�C#��?y�A�<R������F��5m�4���w��xL�I��p����`cGf���������tY��W��L��"�,�r�x\]#� �Yi����=�D?�R��0�j�8�z{5?q�܁%K"E_�(/��+�+}�a�Ʊ�WN��٘$����z[�Ưi������̅L	�?����s��h.4�Bɚ�+��L;fqb�d;� ��.����Ѹ��1���a�@�i!�Au�����Jh��)-;��Kc&H�a�?���U�6�Z�'�qӠ�C'6�B6���t`� ��:o��LX9�'z�ʊ�5 d%na�9e	Y�.x��%C�Xӄ$B�09��foݺ�[Y�u�����A�!G>���Rg��K�m�ܼ%��p�C)�^O:>�*J�hT�+<jF<]QL���!D�@�%fӳSZ��@<xHGԋ�����%]�D|X̾�{�^fKC�)�7�Oh,_-�6�d�*���7��9}���j�O�:�� 1�?��[����<�,�Zgp@�i`�#;�6��=��"�l�憤��{156}EE{���$��B���}�`/�ׂ��7�}��~��W^��V�ѣ�ӧO���)49o%�����@����)Ds�.IE���8m�^x���Y˨���s���X�#�Q�g�n�!Z����	Y�|~~�,�����H���\_���f�$bH,�o*Fc�	���M ����������3NS�|�v��Nh^��0^<5da���������r��w%K�ǒ�g�Q�*j��������$!j�*��h�Y�o۬�Ѱ�x�	 }��g�k<|���N�g;H������,���>����N��73�ol���e��#�a	��e��5�n�a/hEp7�ՠB5L^�*b�@nޜȃ�� 7�l�	=m=�&)�c.����C���E��m�$l�^�H�<�R�26��j��g)�G���H�pH�iZF:k_L)qL�$V�ey�Enm��@)	���%n����)i�'��%16Ǟa�uNaVC|���q#��a��<�e"Y�ö�?swT�JxY����9�yd�R��pɮ���b����0��qF�b�Eh��C�Ŏ ��M�6�S�	꤮�����K����S�K��M��=�^$���o�J6W'������f�������?�"�L�
ss��yƄ�:�|��ơ�g8m��,�ϭom����ڋ�^�l�����op/�n�33�Di���9��^�	Q��l%Y�ȝ��؈��&�,z.Ij��v�"���E�w�X�Y�m�Y��c�_��w=�����*C�8�$۫A�wb_a�2IB0-5������+������
|��H/e���bA���ܹS�� �p&M�&��q�u���/��צ'&;E�6:w��Fe��up���*ke_���A93�ऺ,�#]Zzli|R����_�ɌE��Y��Ci��I��Ç5cC���ZGU��-�[�9/���n��/66v&&zs&P�oƄ/5l��.��N�)fP�Py�?����c�b�f�Z5��>�TW^�tiii�g?���#eI��+��k�5��d뻕q/�����W_�Y�I��8��bq�e���&Y�� �x㍯~����	W����{�]��G����Z
�o�^��ݨ������^S�����o�Vz�&O!�"g����1~y6��A�_h��ڌt�X�œ�1 ��{@�4ݟ���y�4z^n۶�PN�� �"'SH�l�DJ���gi��%���Ѡ6Db/^$��+Q�z��c%��<��v�VM�a�ȨQ���4�;�%2ltO�4�#�������m���#-���-8�;2�\�w�!��ٔL'tbU%��gO���zh?m�g�f��|,Mۢәq7�]����B*H��P'zǓ'Ob��ZcP/B��FrE傔'�G�D&�u���}�:�5����M��n�����*����������V+����ꦟƝ+�sBn36�a�{�l��P�L)���!v�mp���J5OnH0���h���oR=s5�DF	��(6NMc��j�&1F_&u\�!˸�#���(��I�m������8��T�?ޗ��a��.	�đ���}]6�{m ��{�|#���5B�>����]��4�?�@z9�V�q:�Xj�d� �Ϧ���z�a�V�D�o�\� ܚV����R�Da\�������E�C|�
����_�ԑ����BY�S�=�km�=~"�S��q�0�:�:�� g����r�"��(�k�e��#˃�;� 5_0���Q*-���:�؅D�(���2����ftf&�Xij\6���y�[nu����P' q�V:g�-�-�����1�}a@!^�Z?Զ��В�D.t��k�~���̶������ҝ���������M������?��� �M��q��
I�|��_|�E����(�~�>��C��p�s� A�d�V��΀�4.\�����������N��������O>ѳ�R��+W�h��-�.[�B���h��-�D�j�ZX<��z:�����2�_ H��\^Y#P����� ���{��A��?�������W���6
}que���3�?�фi�5��n�����M���q������c��u�MX9��r��`�/~��M}�����ֳ����s9S������6�1]71&RRM�5m������p��z�6��}�Xh���i�	�$�<��Zx��:�T��I:�B���]�u��rL�'x�Tɀ��녋�LP��(�L�Y�I���I3��'�G:6�
]kU���j&� �ap�,D����ӡE׌�+J"�9��t�����N�F0֠[�p�aq8I��gVW�h����ҝI(ζ�GP.�2���`�P�cp0A�]��bZ�#2s�ae���l
йغ�>��dY�b��<�/l����n|�@�/E�3Q�"o�8>SD
;r I�R��5�i$LvF^��v��t��"�{�Q98M��%��U#^��X�ãq��X�O�Țǳ��5d���VV��vU4 ?�;��]��b�Ό���H+���&��b2�J�e��/�@|�16q��L�z���u[�'����i�[�o��+t_�<v�i4�f�#\)��l��`�@���ʪNAۇf���U��`>��~k>�ix�[��?�'G��<�na���"�X�����,���D���ر����a�,I5f�lm���gN��tl�G��θZ���M�����.k����y��%�B��n7��ٻ��,Ov�VZ�v�ڊQŶ��C�=�GW��xߨ�V���&�4�`;�y3q��y�}�l��ܠ�8�a�[�#o����b�ӛ�Q?dbX���h������»�WOC���-zb��ةǎ]^�>����c7o���}���=�&k��x��������N3O�6�SH( D�n��e7��Փ-D򓴠t��>����J����ٳҎY,�e�Ɩ���m���dП���y���ۿ=|�0��v���P��\2���>��d�[F��R�2��5�L覬4����o��I.��h������y�4T��uV=|�;�UŨ��?�я�F���{��	��H3}~�>�-�����sV�z�[�(tq}�@/���׀�
�L9[�v�\l;Ӭ��=zH������PN��;u�4�$�5*86��瞃�_�:r�����9J��<y��͏ˍ��2�f"�!�"�@$���A��2N��۩BНg��VBYd/�X!й��������"�6A������U����6cҕ�2!1 �� �j'�:����޽�X��΅�N�*��=���R,�,��@��^�т�e��|��d�#�������bM'�hLB��uo雺�����H�e+�ɡv2%K5�%S���&�h!��DG֧��J�|i@=�1�h�1�|������	�y�8}���"��̒,2l;UG?�/���c`��ظ�&)0�7n�"���%��P��;D�����ȧ��e��U^��r�ʋQZ:y��hc<��{@�5����?����N�t�-������7�n[# �����aJ���#0<���g8I���F�i�p;��&:Y?���G�TCO��"���r i��"�"�K��65ѕ��Z�����O~�c%�u��V;25����+��&�#}��Hb�� U�7o��b�*���#}�?J��bݨ�ݒ�k��A�Hƭo�T������_z饍� ڭ�ϑ�*m'۔�H,:5���z8��	b�����JpP��~����"�%����FA�D~	�-P���ւ�jdjm���&M�,ZoS�1+���i���j >4\ �S�S�jt��:6�;� 딿��O?�TCT����K����C��s�-�^F��"YL�ͺn(pƢ��%�,-.�����������ʇ~�%'�<������N�&�w�;��vcs��@$�!,��n�;5��nݺ%�5e��Hl�Z�,�eo���oY��w�_O�,�����;�\�������8<%G��������Zt�XM�[��c;#z�>XZҷΜ=Kb;|���T�0��H�x�$�Z�0��V�Y�s	Eų�.�=l9�Դ�����������׮^=q�$"�O�mn� T���$f���7�Դ�Y�@?���1�(�Ɂ�C˘v�G�lv{?��jf�9��x�� l������:u_����`�(�E��y���Ç��׷����zA�=jkx�6J"4��G�eiF���c�-4���bj>xe�X.����V���چ<1���v����xL1��9P$���	_	)�xt(���"�%��?�߃7��q�e��&1�9-��ʼqP'6cO�D���GK�yXY��F��p���*F�0 �7�b+'�N㨺�'����*���)��o�F_Q����?q4����w�aW����(
��>��>+�A����n[QU1Xى�˃�^��&2h�<ʵ~���*��{�6�̿a��ƣiI,�,#�q\�&#�����A��dT�4~����06�k�Y���u-$�oKl��ɻE���;0�Q,�Lb{�,F?}��h[6�{�m������wé�O�Id2�,��9���j^U�?[��Mcd��� �i��DO��M�������Br��q�ĩ�:z⒎�+_y#pd���Ts����v���������x�ԩ���L��d����WU��$[��;��7U��IC7�I�I����cL��b"&������d=Y�K�'=��tv+VB�.^�S�̓'O�ҝ�Νc�������9R�bG\��M�S8ɾ�⎾r��� �l#��BG/�Zȩ�XX��e�5��#�$B���W�[g�ٙ=�w���BĖ�8k�X]\��IbxȎJ999mߝ�"5��N������$vO7R��p�s�p�eC� IL���B.��X_�(��Bo{m������0f\��*��4@O#=�Mp��ܜ�0
K��=X�5m��:�(_Zz��3W������;�v�$��oH[��3gm3N�G.F>ֈ��m��u�O�A��. !O���&��u�L�<���E�+��R`�^�.��ي> 8@��΅��z�"Ʊ�>�x�B�ڭ[��:�_(�h�t�9���.�����#�C��\Z��p��vM�!#|\�`� چ�p�?�k6���0���d�TbL�ZJw}ط�9��,�)����䎅���s���jgk[Ǡױ35,�hcs*�oL�}��RV�D4�iKE�����Xd��<�������v������W���h�2C���a���<5��v�醵h�'	�_iVG�Н2�
9C�S��/ Op8�2`+��*m"ڹ�ɱ��amKmߴ�pUlMF�.d�8��Z����_|70fZ��k��'8���&�+5`Y�81��Ջw�'HxͿ7�q���\:���ۄ�Yn�����[��TY��n�W�M�ϥ��,�&O�d<u�w�E�nz�g�'�?̀�����F�N�NbO�Q�ƥѼ;�${d1U�";֝L���ک�g�X�$%D�`ѭlk���t�H�F��<�jP��{>�tee�D� a�&��%��� �5%��	X�L@IV'�
�4�y�#�O('��$Ĕ�7�qB���}���Aõ�T����!GLh]e�J\�z���+4$�|�c�Hl�<�"C���8�G��s�n	�Y�ʡ���/L���u,ܷ�9�f�
��q�$���Nr�٠$6�ղWkێ��̈́mMn� �>�F�5peƪC�La1�]k�C�*��N��q��rVs�n�~��k���)ը.]���s�5["6�X�'&��F�B�I]�|���{nX7S��?9�yӉ��V5�#9l�ƿ�n��$F7e�7"[�?�* ���H\�pb=���6�eL�mEڛ����ƌ�Ej��8f�z7me��8��o���ulR�P��!���)s������\+�F�uho�'�r�{�p	�d��{��N�M�v�i�(��?�CHq�����I�}�����N4�'29�	���[j�.D��֦� 1�Y_�������
벺�I(���$Y�g��!\�=e,:1�,�.�)t2��^�B�[�tT&(�\@��{f1�MgY�֙F���1��
���x�zȖ e��cs[��=/�,Yc{�ȥK��So} �}��^o46��i���*�U7$��I�\��M	C�9S�O]�73�P�I�d!��;��I�Z�:�o�q�V[F�RY�J�2YW��|���̛&A3�Evo���뉟�F�Wx��Մ_��]$����U�֫����F�.��@w|��'zI��G��xi�ϯ~h�vGU�'���ZI���.�s�9��DA���V�SYڮ�J��T����_�+�[� �tóg��Dե� .�?�:"_�u<���ƅ�[�]�.���2�;��+K� �,�j�5��ξp�23��s��t��c2ޱl�h(��r[�����՞nu�:��R��3�+�Xs�:5=mv�[M�>�yv��.\_У�"mu[�O���x��ѽ���[幋�>s|�Бc'��R���s�vX��c
���T�!�4$����R�bn~WoG��� ���@��R+�#�&1���vJ-��@9x;�vA��qUtG{�k��u�$a_���fp}�Xa���bp����H"_��bxb:�<����}@�6�ZCkrZ5꥛?���{����~p��y�[C��S��ιv՗U���p���2�7��l�w`�%�K�ys̀,��§���GZU����99�>�t��k>�����ƛ�rL��"�eb�'j��}��a���8w�����ӐTџ�Ѩ�2~MF�X���S��p���7"u�9MyL�K�5E$�toA�hN���Qd�v��ӈ�8>E�,Jbw�mnn��P�Pζ���NHKp����y�{�LO��<���c�A��D�lfÇ
1aYz�W)�r���/n~�X�)�(����q��Cw�z���6�zԀ����WD$m���7 ;,.m9zɠ!u{S"�H�����V�7���žL���֯�ewd�=$�d9K(� �.1���*�N9>ҘP\�L�7I��t��� ë�*�1_k|��4��j�&� �Uh��f7�6!p���Q�C0<b;��b�[�#��ج�<X�}B��@3�v��_Q�W(F9����S��u=�����B��/_��Y%(�c^�:w���z�_����Nh�c��LJ��W^�K�@� �ŋ����}�j�(c������[�2l쐣��g�ȧBE^�vMcFkf.\8ojT'J�ʄU�|}2��L0��[�e����)e#�ۄ)�}\�x$$��?jT�U�n�[���g� �\���@Е�8��҉�!���։�#W���z
Ow�����u�ݿ.5p���~�[U;#B�uK[��E���cW�Y����+�to�Q�L.�~�Q(_'��LQ!��8f(i� p�?��J�<:8l�1H���[��9;�������#1��,h^�W{7M�Y�I��V1A�Ԑ_�5.i��A:��pg �#�H J-K���/�tn�>��<����ߺ-5V##5@a�v���6��9�@Ilq	�_�U�9s�y�9M$�[�9�[�����agWI��?��,~�|�<W5Q����Os��}�4�F�`Q
Y}�j�v���fD���ͭ��I��VE���QI�R�|����#�d1b�Do��<���#�0�/��	C6E���B�p�`Z�9���ޗ��R�1	��\VE�3�nB`�zr61���8�^��n�$FQ�8l4py#2��x�r�J�b;E��~�,/�/,X�fݣ�\q53bI���b�^㿴1��z���rnnjs3p�Й�l�$� �Ǒ J�&����$=7���X�*�;[;���(q�fxSt]&�����PԙL�;���iF��!U88_���Db �!��G�N��2�����΄�Y���k�c�����<MN�ܬ����tc���}��k$��X�T��*��K3T
��D�Od8�yXnlo���XO��N^��n���z��,�BI��ҥK�D"r���n\���>��9e�{�'p��5���������/����vp�
�@��ɕ_��������z\���c��͛���75r�.��d/��!-�u���o��o|��Gx�����C��ԑI,D��[::t��B���|�͉	���I�.�$Ṱ����������N�����Z1]���թ�-��)��ȡ�٥D�k�AET��{z$��'(Hggox̡�V�Ȧ֔��S�'m��Y#�WE^=�������p��*�gCxBS������ο�O�b���X�]
h�����|fɓ��5�M��T���+��C� ����G�3���9ڙ�R]����^7t�M;+jp
�r�|0�=Y+#��g�L<u`'���#�	J�ļk$�`���!�x>�p�>@���X^ǜ��L��-I(W��<1�4X����<�{+c3�,2L�&R�C�޾Z�"��;�g��O�D����h��J�2W ��:%���ف�<n$����Ёߵ:�t��o���O��T�oRE�������O˪}�;�F}���1+�]zh�Q����t�"�v%�� �p�	�#��%��]��I(�j4 v��N�����8��kĪ���:�1��=p1��
�G�#p'�n��̤��[<(�DL���	�*rSy�䩙���f8�B%-��2B�A�*��UB����g��Jb�J]��axP�I͗�G�ہGR�+O��P��&F߲Nu��<
�L��\D�c'�G���ؙ��w޹�ɯ>!�����(�q� �Р�PxT�Ia��Qr���v;�Z��h`����c��&B*��埍mDE�aס��C��[P&KKKz}~�N(�>q����{� ��k�zk�qHx�ܹs����� L�8�_qt�Ǐ_�|�c�H� u'z�^y啅��[�n������Ώ�c�]��s�=G�������'���%#�x�F(pC��`J�k�A3ip*d��3:4��OO�(�Z�1��~њ�55H��4	�|�^�ر���v]H�N�����ܻ���CW�oώv�?���kYB���D�]����x�u�g;?��@���^{c���ߐ�SS����׵n��H�-���C����M(���tCmձ���7
����k����lmm������I �57oh,��`[[�nY	y2��tp��,�!�9�U?�Y$<�b>�G;Dy$:q����c���4�]v$3�؜���Pc3֊���Tm�{4<iX�@GQ͑4U�#�4va*dr��'�G~�1"�Dcɗ�D�_g���R)M(YE�f>����C��8�=!㠃���e���j�fϨ��d����(�#_�,p�{愫�؅�,0�����F�� #\�Q�5����<�Fv�nJ=0FiY��S�J�Ц��L~�xY��&��%��ېV\+`f�l/b�6�|���!/��N����@38�F�;��2�h0��$�z�>�%KK�Q�d�|��/yUf�Þ�'�I��@!��ٗ�=�=�T���7�X�]�>�3�J��4�_�>����qǵxY���2j� �_UYnZ���Z��t��<��\�ql?R�:sr��FDW�$�Z�` ,e�*
)��94
e
-Kf��B��p@���z:⬬&�ժM&^��:����˖���)U��3c��H�Ha&�3-��,8��X۴�����(���LEiy~�'�b��m���u�t�tr�xw�z�WlO�Y��5g,�S�d 0��A^�ϯ^G�[�wuuS��uj��Ǚ�gH/ñ��B�j�>|�9��:p�S�~�����''4��CEa�-��z"~A+_X�[�ӐFCE�Jv���E?8Ȯ�����~���+J��G7�{���O`D�]j �v횾��K/]�pA���=Y#�(N��?��h�mgɐ+W���BW��D��Nk8��=�N��9�z���LO�o}�?�ai)+��2G����]�yet��6�!�ӈB<}(9K))�(j���4$�_g�>��h���[��W����&o���M!|=���ۚ@��	$��$�[`q�����l*��hw8 0�Ϸ�����Z�̅��>�<�e#��q�2;ULBhG:� 틎Ь�,���m����Rlf�c��0�q7�_��r�1e�lD�(����6�mt�TYu{u�Cu�����4�&	u u�*
�}�zr-�F{���]T6;�F��r��6:���l@�`2s�W�ѲA����=��R��������|X6
\�¡��CK�l�e��]�(�#{������L�4��kP�:o��5�Wiq���A��F������s1�-&�m���Ĩ�0��^�듕`��LΠ,�>+:��W�JZ5m�<"\L�� ��0z4���Oq!�b�?ĀlGr���1���^t�X��E+�~��U�}me�c�D��ᑉB (����p�EX^SK�F?	�_�AHoY���#�?������{�=�p�4hi|�.����\�T���ؿ5�����G'�s[5��V�R+iSQ�4ƍ��ݓF^��h[���3h�m�tդ6��=I��
!B�M�׵����S��z��Z� ޅ��^�LˬL����ֱU� �q������Plaep��֌���&�v�a$$�ȓ��5��{4�f#Kzd�Oઍ^}$k�@� �m`���L�V?[����ga��w'Q�(ɮw!�˶�0�����QB��Y'H:�igW���҃�7o�V��R�y,��裏���&'�|sJ%*��a`�tޚ�M��g� 	3��������0r���Ν��/~�x)#�xH��ٟ����A����}w��w�ŵ�	�Gc~��g%᫺mq�"��o"]��
�/Z�*��e4���&';i�)+��/G�9L������:~��|�/��"mR�-a�ӧO�B`b%����{���?1�=w.4�	����_��m�kӌ���)Hb��:�:}�N�l�ڼ��ja�<vҤ���C"1�(�����@%M E��)˺��6I�O��dL��[GvX6���,5~nn�ɓP��7={�,n T+�7é��<��w�������5�A�P0`,/�c ���[�LL�}๧ t	�v�C�.�f)����.U�n��vB�:0�U���fXS���]F�0.#��Utq��vCi��t]�a�ү��=��8id0�uq]���2����y�y�J�q���o~ T4QQ�}�Ou����B�$6Tm|���l�>Gr�p�1��oY�f����㛪!i��#���hg�Gq?L��-�;ϩ$������T�w��~��-��+lԏ�����CgC�J�"���C/��̲��RT�VZO��'��A��F\�F�3�������>%f�#i�S8J�Q�-��#QZT;5dE�G't��l�|z7٬�ȼB��w^:NN�ѣ�X7$1��4���;~��Ç!�BK��Ֆ��̐t�	���u�������-���L�����"�%���W��#�#Ѡ��s�BI�I���r��Lp|&�ǒ����]ܼ��矗��w?��3j&4c�b�щ�g��u���k�\R�\a�T�vŮ�ͧ6��v���\x�HQ�N�8A=�~�_��/��/D�B��s���k��!=��3��>����o���_z�%��r\������Y09��s�f��iXר���w9�������O�֟����Y���W�E�3�&:h�D�%��6;s�t��駟�ģ������s�"��N��M��zA}��I
���΋^Y{ffڗ�_t���'��W�jN�yW��Yz�?��?�˿�K��<s�x���c��[Q���0�h�?b�Q$E#Kv<d��VF[��h\#B�R2��{.?Yv�uܓ�����ߖ�Q5�V��|33�IZ�.V@^k�^����q�����C���i��:�ĉ�R5����i��- ����T��2�eЇx��{�d�u��nS@�E��fWW�h���Z��,�7��<���Ƴ8&����	�
y1�=! d�)�u1����g�5�,'��_�Bi>*lo5y�O$�A۶)b��&���O,E����M�*2�=�/ͽ,,�`3t�9b�r��'�nx��q��!2hz�,/�ѓࠚ�ޮ���,���[@i`Ss.�n$݅c�[f|��_H,��n{k(<�A�dN��Hf�j���v"a͑���j{@���
r1��q�V�Y�!�D�Il�e�L'���IL�-d:p���~�?>kT��>�q����_i00.c������^DT�l�U��U,�2�nxe]���!T��cK"�<���=|66gM��q���XH���y�U�I�U�e?�X�ig2��2]^~<���<I-�pu{}�?�[Y�]�=x���~����xr�:A�n�l����&{�O�Ze@w�������"�@($I���-K�.oBd�mB�Q�Z��`��QU>��Ҙ������x��xL�\�v?�����d��\x���D��̬��$i`�5�3,��9Ip!eN��5,*0�3��2����s����N�t��ʦ�m?�z:���w����T�HAj��Rx;[�溡���ϟ������xDe=��y�� �'����z����ŋǱ�Zht8�����+W��u����}�k�Ν;�I+]�W���������z���G�����Yy��ѯ�گ��t����Vp�|�ߐ��w�1�ڏVYpZ�S�g?����w~�w�q���ҷ���������0���O�ȃ�`4��~�'?���56��^x-I�Pj�u��zS�9�4�L��,PS���e�2=��_f��r�#/�xqԱܔum�W^y)	��k��.-=|"��O����$�;iid�ئ��@�������!��J�dQ��m����O?�R�)�˙���	;��?��?�a��ܙ��6��,W:�[[�^����١�"_[�2]Ly�<�"(��3'����������ν{����^J?R�e���s�]z��kk��S><+<�n�������������Sdcf:��A?�p%��V�ȡ��7,t9��|�H(�Φ��΂�\��U�Mw��Y������e�C��&|sk��͛x�t%���z��.<u���zh��3���,-̴�d%1G:2�MM��U�I
�<^Y�X?zH˽y��-���\��BMa�m�6A�����@�#�?��.sqz��ʴ��n�@h��a���m�T�lyy�I�ZH{om����J@��n����ɩ��dw4ll��<�����Φ�977����,�4��y{9�Q��V��L�:'O�f{��c��5�"98��bב�L�b;��Hci��]��g�d&'��Tx>h��^#�[�	~ld4z""T$P�aA�m��p�`P呇֋{���Dw���p̷۽�"�����病���p�]`���XG%�m,iQ�(a�1-�f@I`��UV�8Јڃ� �Bm�pe5���Dk8?^��m���SK;КChd<�y������`G�jwB�m���V�^_ii�e�
����55?Q�i�TТ��hE_�����Ӟ��MK.������K�ط���P���sx:��Q�Cl4=Tꁯ����P����$:k*���;��>B8����j�[��$����<؅�{��j%iT��%d�؄�~nvZ�oq�0f�\_���-2�mZqR�����h�Q�т}�*O�n�αpVM�$�%��ƨ΀��ңu�9��!=��N�&W:O�����W_��[�a��g(B "�cq�al��I>thA'8t#����ڰ@���B�����S�]�xaqqIoC̞�A�c����́�y���ֻI"�X�Ѝ7(���z� �D!De�#C%���&�\��bUia�.�C�H��]P�=���]�B���S�y�1K�J�K�Yi`����B����E�V�ya�����A-��]W�S����5]���.��x~���t���홙�G�VL��<9=���Ǻ3f�[o����}ώn��gWS{ɼ[]���G��w�'�n�~�|�?|��ו5�������!R|��}�QO��H�@�E��T8r��:�������X�e21�G�LBO:Q�����o�������f�W��j�.���uRg�v��B��eCo�$�s5������D����ǟYZzx��Q@[E��?�/�2�m)䤯h��^O��FhT�Fׯ_?v���L|�t�D_|��۷�i��.]�y}��%y4��� ��nܸ�-񕯼�oi��%��ͨ���,pi<����䣏���Z/�(�z�]�ίm
R���Ȗ&!�z!��b��v΃k�)wc���1�H���S�i�=��+�������O�U�?�͛�5 "M�ÇkVL,ݮ�k����e���R�f5u��8:�s��H"7��Bkok`��5�e9#��X�ɖC���S$��&����{昀�Vd�90�xk� M�����l	�JF�nPc����du�G^Xgm���O^�B�F����
#��HӮ�h[tj@�T��3�0( զ������f��.CO�
����e�)J�ر#������e_U�}Rk�7U����̇�u��i�B�ӀQ�s	���2  ��IDAT�:8��.��e��[b�$��.J�����-��B�
B�+�"�!e=��7y�=�İfS���[3Ic
9��$����HH ����id���#���Z"v�G-�g��N�$&op$?lv���×$���oi� ��Yd��W�d��#KpO�H���z�7`�]�?���Xh��)�]z��v�^�qd#J#��q��,Fl�b<tU�/�08LY&ߴ}������@Y3���/�hX��'�H��L4C[� �b�HX�V��>�Yrxnf�0�Yq�U�W��Շ��@Bׂ�հ�WVv�lpKQI�]�xQ(G�]K[
١���e�x����!��ꭊ���+uJe�ѿ��R�6S0,�8�0԰iqC@
��:�F �FBZ���D �q@���B�Ī8!$������W�}@�e�.K1P��Y����I�ӆ����7��\�����J&�Mwx��-6RHS
�诔z�o��f+6�4b.���`B��U�Cb�RڜØ�ktC� >ܒ�~�d��d�/y��W_�{��Ư�S�5==e��]i5WV��ϐ�0�7�(zq���.��tҷ�P����{�Ep@r�B��d��0�IF!�[��)N�7K���2y�c��-���sҲ�����e��{��=��s8wiй��XY>56�.^YY3>��O>�_iT�7�MΟ?�O����� ,!��������I8�ʕϴ4E�loO���t�_#����s羖F����25�@�����TwH#�L4�P:4+pl���
��@gΜ�`
����� �!�N�~^�*Q�FOfϖ��W�,2�a�P��z����%Azw��7A�LLBK���7�^4��@��ڳ�׌n���1��^D�峲���@CP1�y't������*���c� U�>C��ڵ�r��y�%lv�uq�u� t@��.b3m~�xT_*yW"E`k���+�=���Ϊ�j���4v�$�I5Un5-G�~B\��]}�r����2�&C��Lʋ��������#H3J:����F��ލ�jWc�U�8�cc�}�ְ����D20=;�l���ӯ��)'*"Dv�z��@o�+T���f$�?�R��J�(�K���5�Bh)��Mv�7*u@இ"�V��P��b& ��==Y,�ǅC�Y{�P�E���θ�Sz����|YyJ+�lW1����D_ڱT��qg�ƾ�M��'���F�[���եi��^���H5��g�r_�N�kȊ't��>�� 8���C׾�7�[�%�
��eώ,�M|�4��)�cHsC��Y6�8i1�)p,Q������(��"%ܖ���H�DT�&9(Y�۞>u���E<+�4�=��~���#G�zW�~�s�ņev>�HBc�D���b<$� 9��@g-�0���zߝ�mf0J�^�;�8x5N������XA5�m!h;�|�X����KQ�KS�Rc�.Ԇ~�k���={�����n��S4rV��cO�_h^z/�p���T ��&Ѱ�VK`y�譴)�\��'��S�`t��K�`�&)���:�{0�p�c����Z[����8/�8�&�+4���ՇC�Б1�T降��&ƙ�9X��R��h��W}���i9��nh�}W*3ڧk׾�p�<�i'���+�/�y��� ���3�fϒ]�y�9'�y��ք*�P��A��"C�,�%E،��Ͱ��C=دR�я�D˔M:�ISj4�M�Mv74��P3n՝眇�o�_�]Y@�֍���'��gk}k����*�>�@� .��;�o޼�E����Hc'�w(q.o/��ҝ�{��s�V�ӏ���̎w-�Go����5 �_���+���g��^�����Yk�E�:R�''�1�!���*�T����F��8�����,x�u�ZY#!(��k`Z�L%
_8��iSP#gPG@_�{<q����K(4C+��#a{pD�֊v�~��k�hF�K�)F �S��4�_~�P���@����,�N�������i��^;;�$tS��)�¹(��F��B�p�=�glmz��1���VUa��o�3\.�6����"���+XÕ&���E�֑\E�;r�,1ݭZ�F�0�i�����-��p��F���ƪ�X�&��N=B;ф�D�1fL\]̢��d�~��#w��V\5_r�7�R8�|^�"G5p�+�������7G���+�q�	���i[@�ȩ����)S�	�+&p��Q��սm��z�&���1C��	��*���|<FIH&���'�eD���P�8�D7'��f���pJ#��3
=Q�Ю�7���$����|�^��tc}���8�n�K .�� i���&*	"��j��	���P����g��S�V��n���� �Мc4�P�^O&�'���C
r��-y�3����ɿ$�� /ʓ��X)'�����Ւ�i9i��n޼�ӟ����	���AHKь���C'��f������Z�F�	��Rɤ� �.��:��J�ՕŻ��b�#LS*��&�e�A�|:ү�ޠ�9���ay��
��^�l;�r�ǘ�odsV?�@��d�:��/gvF!!Oy}�DB-�N����GJ���'O�Q� ��i�Ҧ=��q�)dm߽{����r�2�P����=�1�����F�Q������Ú^)`���~4�3���/BE���t��a��L���M�;h���\X���
�Ѹ
X�j葕��[����GyԻ请o��<�w�4}��_J;:G�X��oI��h�[�D\_��b��d�,�6Iٺ����z}�������T'z� z�(������u랮$^2\/�[�i�=�����=�;�����s�W����~�!�ϚC�Y��cIe�oQ����u�����\{O�V��</���n��TC�����Є8���s������������5q�a��^ m�Q(����z%t��֜���nmoI������ёe"j��z�Ew�AQ2zJ�,�}(��1Ǘs�<Z�9:�8���X^�!�}���L�I(,�~cc�������
���N��EJ�G�z$�P�N�9}��^�a��2�MI] ׶<�)q/�˼2@o�m/��]��]ZZ�B��H٘L�ab7[㦱���[[��Q� �lc�ʷ��i��$���T��{O�z���1�bSSu]9h�[�/^	�R��M�e�
��9e�8�UL{�nK�k�L���X������"�����N묩c�Hx�g�6���ѿ?ih��NP9&��:����L*�x��݉?OG��Wq=0��<��B�[6�	7�$=$<��"��K��+N�ʲ���I,�2'}�2�f���َ��ΫC�r���CFftJ�/��SN/o�f<�0Q������TG�9,���{��-q��_�1hP�䩉o4"����&I`�MC�:��Qh-jo4z�F�0��N �<%sTZH_�d��*��?�x��Y]t�Aq2n�<xbK�0
�;B?:�$w�g&	�D̅l��Bw�z�5����r�%d#����>D����)E:l>ۦ�א�0q3Jt�A��Sg�\��I��l�p�����;��$C��-�L�,./!��5���ĹFA{a?t��.�1��ӈ�*�RPt9���Z�4{��h���� (�"�z@�cRS�`G�!�:j&�q�u[��D���]Cl�2���\��������أ�b�MIơ��+���z(9"�.���m0���l?�jt�c�X�֖��.~����3)J�`����RiO�� m'>��3���a�L`������� ��իW	�h��uC����N/}�Ө!a���S&��[�ɾ���ƪ�����0��Yb}Ϟ1��"� �Y�*8'G�5���Z|��=\#�1�z#=B�M�q��e-�Ejԋ��e�n�ҳt�H�G�����:�4��z�믿���.��B����yQ��p��;�u�����DU�Z�p����V�|��ﾫ;h�Z��[���>j\ B��9������,��.��EA&�e
��ZA^��O7y���s��k�]�D�!1���BJC��S{n���w�]M⋹jƴX1Otz��\�&�7|���I�'3���@���hl��d^r�{g)6�%x�\�'o��	Ǥ�]t;���n;�Irs�NGB,��Zf��w)@�3~ZX�@8��J`�G��Mq���N�[���m��O�.#��<n���54j���b��i����xLL�b�J��0bhb:�y�Q-i JT���=7	>�=ƃW�]�:�g�b�$���ę���B��:`���,~1�C��<����c8���<�|w��s��Ϩ�?�M��:�$$����ǖ���(�DЃC$B��a�.#�` ��Lf2�>̣N�S�M�N�3��33�#�v��V�/3��h�U��8�_�9��N�1>��}�l���[�|a�N;O���;w��x���LyIahȬ�v0A�Y/�}�%�:o��f�Ο, ���	/���q���������"�D���!�p?�u#��������f@����,�^�Y�C^�C���`�D���s����h�!��6p�n)��;�'Ny���8a���9��������H���?~��r���hV�͉TQ��0������,�[���˶��ffn��ܦJYo�_ZY�p�V������/��E���d�qH{8�-������_���E;"g�2�����<I!�PA�f�E��Y�Z8�J�h`��j�{�=$>�_=�ƍ:G��1���}��U�O2��w����U����M��Kب��Ñ��gB�	��!�L�����Y�������lRƑ9A<�=Ko�c�$�%�xv6杙�kĬG����܍{K[����m�e!QM�>_ZZ���{�^Ү����Es�	�]�ۘ� �d�8�����yv��y���6!�#�Lr��ua���՝�m�8	�BO^��>��ӛ7oj2���=��\-w˻_'Yؘ�hn:1P�O���c�}f{@�Ö�ѥ��8:R� :�����&�ʳgV�Y�V�?�҇Z,+҄�k�GU���!��m�;HN'�a0֦�����i�T�S��Lb�p�>HѢll/��Fҋ0�ԩ����!uAx�\��5��4�A�!Æ�� S�D�+��ŷձ���ՙ�:��chb���T;����l��u&�_>~>V9��p�P,��n�Z�^#�\�" �j%�
��`h3Ef��=MB�<Pv�!01v�ѥQT�:0�~�B�<*�/�[.�nhz�]��1�d���e�`��!����,=�I�E_�/r�N-��m�@�]�gi`�SW�z'�Jtky>�8vYr�4lH�4'���k�O%t��M"�����^�I`��C�@��1�Z���(�A�_�s�Wx���P��-~��X�
��n�%G�����oQ�\�,�bģnM䤞Y�B����o��;�p���5��As�1=�w����[�� t�!)�浥�oI������=�.$��/=eu��5�kYEA@)ב�֡�%�AE[�-ڋ���֕ju�X49��(I����|�_��Sʊ���0�����G�/hk�jI� ��'�n��ū�qr�
��G�H]iH��z��+��䑯-�;K��]�KR�Xa����S�MC|����4���J��"D�v���>�L�|뭷���_k�CQ��Px��&�(vDQ�E�C
�wB6�ҴO4T$����׏��	v�5� JYS�.(:5�nHzǝ;w���N�aaM��+W��s��}���@(�|?��O�Wt=��z۱Q�>|����!J(,����k��yA�����[��&���I�g]��'�i�p}��I ����Zm�j�$0���k~����ߏ�� C�ɻ૸u�ֵk�H��YM�S<=m��ό�&��A�V�PCff�������-����%�v�������GQ�?i�1H��.��zOn#g�L	���
�������?�٠ejTo��.:���(��X�La ���as�%̲�umY�s�H!/���0W�Zz��$zp���ڵ+{{G�uXZ|��w�������&�bbF�l�+�D���˕��7d�E��D�Lm�a\�4�%���đ�tLC��(.�p�7(s�O��!Qq��J��2�P@�I=Z� �AW�e�{{5/a����4�V?u���AI�;:�� ���i�  @w�]:77K�0R� ��8�_y�A��c��k?x�p�04�A7�`>�T��#^��C�@�r�AX#zh��iR�����y���Zb	�7�<�D�8�ډ1G���I ��z,b���j�8�l�A[�y���BN�"���
��$R��h�6��o`/1�8�4����P�./>�,�'�>'�b\��&w|�z��L&R��&aq�=b&�M�e�T����BO�{]�h�<�F?�ɟ�S�����h�(CM����ޡ9�$dۃr���&����^�*m����(Vb
�Q՚�U_d�$	X��1��.��@�B�)��R�D�Y��1R��'H7ݘ�Pï ��+��JBJB(L5Ɓ;��RrA7������/���rt�A-Ѥ\bU����@�Itgu�$�5g$�ĭF�
�@/Xt�2����`����>��;w�
��C�v�I��f	K����͛75)'��`~�]]��{�	�',n89�F!f��5��'��EI��8���IS��C��GB�����o�[S��+��<mxo+�s�L)�����J7��t4�gϞi�)���
j��c�H�P9'(E�D�����ܜ�9�'�\�%mN���/d���C��RB~���)z)����)�ԜY�a��ĳ�ȪN��J��k���u���I��ݻwus�ӎ�'�I��ILT�Ăׯ_/ysIX�B�G?Ε$T�k�p?C���?_|qW�&E����꽄G�jpsаy�1�t�p�^GJT�����`ܑ�$e��L�?�0�%e�{�y]�I��A�'d	JNhU���x��p�;k`�/�ڊp��&"�o��@����µ8���:�9�y���Xy��j>��,Z�Nj͑
\�.\�x�<�i�'
R��;���B���Kf��u|jAd˒<l�?�O?H]�X�#]|x|R���g��T1߿�Y�>��k�m��������&�P�$T06a���x�^�]�
�lH�.��ߣ�["j�~��u��_8��GDmx*�lh\H3>$Á`"!��c�4��������IVK�'�tN��>5%�z���v������|�qp��=!z��������!�SS����X!C�3�+��QH�r�d"��&��(P"c0Pn�t�Vj���r �u�z�6��^��DLpDĠ9r�F=d9h(~"A�I1Jΰ���TH�  4��l�L��&Q�^mccl��k�k6���OQ�#�ǵi^g=:��Ud2���b�rq�0���7�fVyp:F`�nD�Y �-�P\�	���g\�#�{��ݿ���q��J:��kG��!�:n�r�s�'���C����U�Y�eF
���y&_�g�[����	��>�t#�x6�����2g�J�ڠ��g���͑>�X���JC�&�����Ͼ�荂D��b�8����ױ�y��w�ʬ�U�j�����|l�4[����������9���%�D�K�*�k|��l��2O-G��;�;��%!��n�V�LnmY����w�9� ⽞D�"��3 �� �F�R��|��Q��1�4�2�i�^`l/��L���>h�%��.\xt�! �>&`�Q3wR��E��!�&�XCZ__���,����$���0ڈJW���t���}��<E�=�n$�������K{�+
�$L;����E�)�M�חA��-�ɾ',Ⱥ�2���1�mc���w�@UhK;&2��\��}��0�V�
�f� �8�<'���Swx��We����Vt��C��'N���t"
���Tgk��GmD�"���7�����>T��N��H�@8I�̋�K^�MҘ�I&+�wyy�۷���9��@d@���Je7�)���2�^�\��o}K8O�&��WO�f�آ�lI~!f(�y֣�W_�e{��#�'ss3B��j���9�����G�������G�q�8��v���涵�W��8E;����c������O�Ay��Z��f�3�G��5��=LV\�TD�)Z,z�ZEy��4��U���f`a�g���Ғ��vf�=3ϔz00�-1k�^��x"�/NMՄ��v�daa�T<�(�G=4_>M+����)��ah?�A�� ��U�����b���[��Ꜹ��3
�D�-4H�di��+�t#�2n�\G��(t�>$󱟱�P�$p���诘���[,6��J�Ed��G A0�ox��#��'�X�a�h�a�D�&�=UY(��BvWD�-E�Q/�����'��"���ί�+�����$�l�MG!�?z
��v��EpH�ҥ�u�fVI&�c�0vjr`I��,KmL�����|�G���Q6����6��i�Y�����������f��w����-A/��fq??�^v��XX�z�
�=����{Q��G2��nzb�@ ��'ٚ8-� ���y�H��ϾSn��i`�7�uR���	���f��j=��M�#5�l�s����04'2giH��۽n,3d��I+��߅��@i�A �ETu�r;�D]�j,)c�G}P�MJC"�����W
I�iX�, �Q_(#ɗc�s������R�rωac���P�M��b�1��$ec1��E�./E����A�A��)���8)�E�C'�n�H4dA�(���2ф8,A:e8�n߾��k1L���=���ǋ�U�%�&�T�r�+8M	eb.��0}��r`�K`*��4���CҌ�:�K[2���Ҽi�cv�C�d]?pA@�ޔj;p�^M�5��R]��=�o�������A���{<x7�C�E�hZN�%&��%��V!�GĊ�(E(��7�5W����o�������S��ڝv�2�����w��I?�P8��fg���������"�(m8t0�4nR����L��F�u��e^�u������n���4lu��GG���0�ɯ�{t�������<�����x�F�!��|а�N���jaa����.BM,�s���%�Vg�IW��AI�tD�r(��ր�������0�~*�?Ʉ��i~�<�����Ӧ��c5.�v�\���a�R��"��x֊�`�d�Z`�q�SSO�K'��tO�q��I�y��by><�G�k7DN��#Td1�9]�@o�&3��"G[5���!ʟM�XF}�b3��O�!ռ�ޑr�Q���D�H�1����	$��Ss��*��A(lZe!H�q�1��y��&�I�4����%�`qhS#��&H(p%f���	�Y&�!H�L���uj
��Z>ы)�Ip:��|�P'�]��u��O���RN��㒐kM�4��c\B���Ul�z���;�i�89���*�Ȓ��#>���>k��b��|�x�H�����"�[�E�����P�GB�V��$%k�k�u��nHd�q(>�$��b��`C�A����'��zCb����-�:"���Qh�E芦��V�J���7��nX*4���퐅Pt�Ct���c(�_80`�����'FLD�Q��P�hP�����<0���us��=����>�Ջ��IO��X��z1��⠆^��=yZ�ASJ��2��$���[ԍ.D �8�wi���b&YP�&J@D��%�	�G�e)��M4`ݐm��q����Fs"��"��D��Wnܸ����A�![�����2Q`�=B�5Z_���°|L�ΚS�ٳ<a�j�����]���S���`����)*/�p�#������?�	sh!0�*��4wrҊ�!z���q���b�>}���Pܾ� L��G�+:V��#�)���t��8߅��Ðߪ\�����|��6�dG�:��^\\�+���\���+��@����޺{�gG륱��_|�V�����[��w���}����h�f3fDđ52�=�7�2���!b��O���ׯ��o��?���T���~����eudt��c������,u�8���:;ⱈ�����6����~N�c�Nf�%�	x�7"�&j�	���f�!�8F�;��T��m����kv^\RR�[o��6К��е�Nb���tj��bVs۵��$Z(YUu�R���<�ᖇd)27��D?J�2��vM��i���z��Z�X�|S�w�80���FV kBK�hf@pP[�B9�0`�H{��	�g1I�)ط� ���k����De@��Y��Z���&��z!%�7��T���j����@�}`�s�Y�a9P���F�(r�)����
��&�c�9�/ȊO"���+�	J���E���acd!!����W2A��'�x�r��-�+sG_C����逿x����-y�E7
š�@��:�L~�3���������>��Ә+b�E!!83�H����1�����;''��ƴ�ze8!�ܝ�n,,-6f�8��5�BB7N]�0������d}��=��
����fj�>=]���#e�d2�j�.�Zwz�hMĖ�V��σ�#�����+���W���Ӧf�_�I�;����jm�V����lG�Zs>���1v?��UQ/������+��Վ�en�|��H8��������9�9��02�<���˒�B��4�k��ڀ���(���Vp����a�\1��"ʆ����l�N����$f%��rzzX��E'l�g$�!�H�Y�q>q��R�y(�yiȓ'O�1-T���L�x�3i�2i$��-���s����: r�1p��@��֐���'w�ܑ�����3��7
	=ᎋ.��!�V�#�u7�#���8�Y?�|k�&λA꘻]/����Ć�����D�Br
e2Q>B.�`+�T��}���R��~���n�?ݾ�%Nh�p��ZR���0���o��l���X���G���w����f,��
�޽{WX0�����9�=���N ��
�`�1'�9y0�:�7n�~��U����ߔ(�E�D�Գv¯�ʯ�c�lPhB����"�s��v]Z,L�L�!@�����R���H�Ǝ9�����wD]��Yb��>ӫ�n�wN�pa��e�I^��U�(��a��A+T!a(�<�����������H�Ҋ�0�L�lT�����I��<�ꄴԝ��K[�r�֦���w��1R`���0i`�W�y>�c�R�8F-�q�%X'�Qt"1eyZ-���+�xR<�Q�ʌ�`Ge�Ɔz!�"lKK�B��0��X��
�C���n��N0+���+�; ���x���C/f�A�1��xnp2ٚb��b �@+��=�ʪi��Za0�I,��<���F5I(����	���-"�k�/ 2
�^ �I��/�P���o>��?鮋 (¬<T3h�aӹ���#��5�$����'����,�F�h2�BÂ���5����)�8>�����H���8�Ӭ����6����T���IY���=���*Ta@2�Q�<R��q���諅��!'��v�w�܅�D�1�`�R�
�
D�鉑VH�K=�n���RpD�gL<oԶ�P��I��a��#�����5T�1��d;���?}�8AơW��6��~�e �sru�vĮ�H������ ��^�t������n�4�5�����2DnF_W��OJЊ�T
�8z_lM�wku�$�c���by(8B�O�~�)�@0r�%�2���_k�6.�8Ǿ�T��w�v����G��1����Z+ee�G�;����8*tg8uoݺ�BL��`�t��$�
���Lod���Ly4����$Q�ĵa�o�tA^dcb*[�XP,�t	����/�B}�`�b(�I�:b�H��$$Ė�'x\�<"O�I�X1p`�iPt�fB�xg�^�[�" x6��P�����Q��8UO�*j߼y�����҂"U
�"�.1܊�)����]��p�0���6��g�����h!��P��S�ߜ�ӑ�6DDы�s�\<ᕅ7,�?��m;�Jt*t|����ѭ�=��f�a�S=ݐ)�4m	s�zYa>-����ޞ�=0�|+	ġ�'TAF-�2&� �E�u��l�h����Z�����8,'b�S��4�O�����2r�Ը5
��Vu>
�X���K&�u�U*��v`M��m����C0!	��h����P���g��Z�*�ۘ'����
g|�y�0s`�vC���*�lf�.(,:7Bl�a7��S042ʺ�ѣH�ʢޡ�e�T 9���_����1Y:[���J��։<:��B��S2<7�_���o��yc��'s�j<T<2*�H6^?���_��|A������IhE�x_�S�3>$&��f�L������KP�g�k�ί��a ��kF?�7�`��Dw��Ii��n�0�Qu6	�s�N��x4)�@ҦT�~�V���W�k� ��B��MPzmI��tk�a)H���86���wYc�F_�&�$Nh��}C�b�>B�IN�{s�-�;	+�M������ulP?*
ld�}8�� �����c	I�+�D����.�*&�BN��x�h�'m���y�� |9����"��<P�DWs߻���=7g7�,��$��=¡�^D�����@���u%~,f��'F'�}�*B��
��o(�j)�`ZI~�R@+����~������P+q�0P���ȑ^�M׋P���<��g͠1��J�D�s�Cv���={w�Tn!�:�c�,	���&\=88�A������	7�`��CO@a/�I��p���~��;�:E|h�jq�x�
�m�1�>q7�j����h��g����|��	�.�h}�6���Nc�_|���m,�$�U#��2��(�塃Ps� ��v�wwe&W!-d$W��qZ��ի
����h^ZZp��n�W8I���/�W���ҥs''��EwW�K�.�$�Do�8�襬�~�;U[����1�����4vc�ҟ�9S�UA���F�Pն�9���[�V��8���NV}ytt��L�*bZ�A����)�{���26?U�qc�ч-Иa�X,���Z�Ӗ��d8摲T�MG��"��P��P�0�vs�%c�E��7@Ph�QY�㨫ؙ�*���CP�֮#͠�9�#�ZD��$�"V@�I�r0S����P� T�
 Fc�j>8� 2��IbH�r��C��@q77���J@ThU���`�E��\�^Ύ����l��+��0b2aR��?~��`�5��/i2�S|vCO�t"�-���H'
c����?
�>���~���L&��ׂ�������'�c�ܡ:}s��bG��[5��݈��!O!�d�=���ϘDY�z$Є���e��X�����b�$��IǺ<�P��`w8,"�����Q��:�����������o����o-�C�39
�`��Z�!~�;%Ӕ��7f���W$(u�,��ׇx=uo��7"�G�%�� K~��W�����/���?�5�y��ǀ;�n3E2k{%>Mѧ�ޢ{�nKA�&Pɫ�c��+� �P�� �6M��������>��S�N?Pj���~�3i)MIZb"�G�9H��;�y���׌�z8ZZ^�#�!�z�m��@�MMS?p��ѩg��NOqv��YWS�K�_�,�q��0�_}�U���i�y--��k׮��k�֏�,Ɏ0�����sd.�8�~�܀ �Ї�C�?^0����� 45��_R���<h�5Bx�]7��N|�8�!& ��]4����T2b�s��ֽ�<B|	�
� ���V�!ӮO�D-q�	D�5ɀ!�Hv�Q@�22Z��D<���~���2i���}���G���O3{���B����a ��u�J���0}��U7�����'H���.�#�0���R�Z-~t�,���驙�����S+ɬ����h�,Lٳ�R!<�Ԋĵa/�V��X���m	fE,*�s�!'��(�!�\t����,� w�f�V�^.]�|9O=�Mu�s�.���<3?V����԰�� �oij
����`[���\�bv�d�j�̉`�\����ָ�V@���BZ������,s�X�I�jڏƴw�P���,#oI��|�!��M�N:��@��Ы�V��:H&2��):�&�e�Z�
1bq#�!��;�!}���O9�Q�F��*?���M�ЏS|��Dyc��Б�x��	Y�!92B1�[�|!�\�3��i&ܹ;` Q�3�<�cF������7y~�����	��6��f�WN��h"�.��|�� ��5L�H,�H����nR�X��T���-�P��g��Q�!����?>#���\8uK�^���ܗnyi崽eΆ�`wg��';Ϸ��X�;��ă����TC; �Nw0�?��0$�A�H̑��ę枝��OݺuˠL�f�E�����e���i�ܘ>�{�Q�5�nkʧʵ����Is��f�
�@�Qe��.���Y��(-�K��c/\>����[��{�V���YǲR���Ԫ�~�}�Νō	������Bq�^��t��t�W��N[��_����JI}���+���W�V������䝖�i?~�Rӳ�ͪD!IW��
����Q�u���0�:���M͛6��3��l��T��o�N{]K$o���ua������{OI���{I9������ٓc��q��n��I��A>L�����L�����s�N3���Z�s���'թ��LMo�l��Z���j,������S�%�g�F=OJ;&+�&닿�k䷥�<�jż7ꦝ�4),T<�Xh����F�5W�Z�f�߾~������W�v��ֹ��s��W66``���he��ܜ�'?�	�Ys8��beۻB�������F�����Q?�oL
������<K������/�Y��Q6Һ�{�ڰՙY�B���ܱd��4Og��0��.^i�NwNv�a����{�W_}emq�Ν'Ǉ�~?o���ʙ'	ͮ�9�K+/�@�����uy�:���[��ҨZ.&�z�6h��F��۷/\�T��{�������K��~w���+gY��{_֊����6��y��v���*����'(���Z/C�޾mD�:kZ�H*��޾}��,��K�/j&�^�ΦTQ��O)~x�e��մRt�ҝq�� z��N�Z��ށ�</W+ͶŒ���~���79W~��G���K�̇���� ����
ف�hD�%5��t�����@�\h�88�N����&s��eieYSw�jV�5	�������7޸n��,=�'O?}Bf��K�	rߦZ"0ͦ*՝gϋ^l>ۘf0�1�J��лh�Nɒo�Rѹ�W�g��饓�J��=�W���Pw������Τ R���B"b�-�ˤlVH�-�)�h\�=Ry�l���k@��մ��Ң�&�Gi�0��A����W �X/$*� �<pZD��.�i��:���?��f-����U�훭�no ttz2[�mnmkVec�V1����<C_�#�x �0��,�)��F�e����J�g�H�2�9� 8�Ѧgd&zlD�_Ӊ�z���V�P��?�!���k�	�ܐ0+V7�*a�J�f�|W��OBNz^'���Gh+:�p@�� �P�mk>��MZ��7Œ�t{���ߓ	�C����~�K.:��5���Eߜ?�c�`a'G��hr�x3FH'�Uz�pH�z�p�k�s7s���2u�uݞj���Ў)`~��3�z�<&�n�����\0��e3xd6�T�4a�R��uWG�]��*�5���P/u��QA'i$�2��yj=�5փa`�I-��)y�E+��Q1����L��]��"h7o��я~8}�5Dҫ{�W�
ف����lwx�06(Aw�v���X���i��k�}���Sy�Q�=�0_�Tfu^�%����X�᥍��7�i��v�������̛WN9c�N���Nw`�Y���ŋ�_�y:E>�����9��h��ɳ�]c&��r)K�rr�&�?8tڅ{k��F���0�g�J�HȽ�]�k�}K�"GGcXY4Y���i�|���i=Ί̯[�Z��2����tV9�iݣ�*-��{�˦#o�2�X%�Еy
=����9kS8�NH��F�Y�=�����w�5�Q:�>��cc�sS�sY ��<g�QS33S�U>�7I:5oR�O��O^}�U��|��+zʳMk��إ�Nzu?T��LA޿�ҥK���y�Ṿ�ZG��̈́��h�Fz_��׬���z����!�q��4=z���,�`��de��/-����g��%۳���M+��_�P�|��7���#sh�Z��5ȣ�M�»W�w�w%��g��'ͧǇ�'(�zs�^���^@�^c�<K����l�,X�du9�o��}M�2� �X�4�Ta Qk��]]]i�_P�s�Aa~!ӑ867F��@���@n���Q-#���]A��v�MogM	ۉ4�dZӧO7I���B�GY�F�{,�r.��!��Bz�6�׵W=aC���_���2?=��FՑb�
hBh�G��f��ت�4��$�y�5G{<�I%�	��(�x�����8������(��pyՈ1S�Ӟ%/
�P	7S�A��Yk��ΐ�Moc+�^�	�l�se��p�ud*��
8��ܣ~��^�tQ�e������R`c�\;hMZ�1��eߎr�� ��1	��2�*��kX�Pi4tο�;�PEkK�{[W���\��/ w,�'	�Xb�a� �O(&�ǨS�uD!�NS��k]}뎋�usM �����=Z�A�ƨh���Ϛ�X����^L��O��T�	K��Q�/nd�#$�P���>�[�Y3x��ӲP>�Ƌ4��0bL���_����؟�p�p�p�jc�����|��ary��gɄmҗ�Jtm�^���T��U7؍Q&^�?+�I'��$	O;�v(08��+��W�^"҇w�q�:5z.���~`=�C#?���q{ԜcL�QH
��=I���="U�0X'�nkI��N���ۆ ���''O���ع�׭hqyqn�v�&����S���0�|��ֻ��A�g���ýN�Pm4fs��v�ܝ��z���h�i�KW�./�%�˃���������b��lu���R��LϦ�ުI����&���I��z%U�Qat�}pay���a�\h�Imya�ګ�����~�X�*���n��N�3�B����s'g�[=g]v�{����*F[:�ө��n�<yv�������a�߃�P��f/�3�}�|p�[z��ծΖ{�N�+������rV���*�J��E���;w�l��̝����}��R�6����=(���@M�6,��N�V�-k�[ms�),��/��t�Ω��Tzi1�]۸^���Uf�f,�tܖ�=ld�voin�Z�mu�y��̋���c���4$Y�Po̿�����>�ҷ.kc�nZ"]'+v�+��=x�x����ի����B���d��;+Zóӎ ����`{��yV}���7���fӭ��H�jt2U�,��(��������ji��_-v��Ta�6����_|����&��N��L�ߠW-�0�
%I����Qc�rx�7�f��fK���!��e&�M��.v{S�B��z��R��>9ܲ�RZ�����֙���l��С�|/�F�3Р�viǦ�)�0�jZZ�;88т�y"k���f�ߒZ��w�"�M�!.H���n�a��N�����[݇4|L�@@�~1PO��K<���2f�J,��`�鸦O	K�"U5�4�!�Jdd��9���K�M��q<��Y5z���".	Ui�NR����KKc�H�d9t�SĺCg�x�xi��阴�L��Po�{��25�������	H�_M�Z"vh�vڋ��bH�ٓ�O�q�����2#��M$���|��m�|xy��M�"H���@�3ބϠ+���@�$>�L<̝yY�}>(�brCJp%���j�Ν�T�#"��őz�D{�q�7�5Z��;�;O�.bTL7��IN��Z(�IPb��R'��(����.JѶ �XLó8�����&���=\e��1.O�I:��`�0$�RC���Mp��1��1� �hj>�H����7�~���7���U,�	�(s;
�ܓ!N�aY`�RU�z����0��4��@ľ߼8���f�B�P븙��D��/��b>AI���@���JJc'��j�������JJ�VWb�����bLd$@qL�gH`	Q\��(	h�@�c��?�u�����>m��]�|=�"kG�&5����Çޣ�:���t�G���}h*���`���/�
u��2�{��o��?�s��y��E����9Wi�s���9�k��/�S6�b$8�)9��0��-�Y�%����;�%�|�-�lm�p�e9��ZJ���$��)�����<X�|&]O�mLm����͛�=�h�ܶ�n10��)z{��e{�Es��?{f���_Ԝ�?(�L�=�D��3͂�yϵ�`�Ƽr~ɰ{�Vp���gjfnV�9J���?x>����UK�#�g{�'�����Q)�i}~�KE��WL�;��t��َ��DQ׉����:$v�f�>|��Q��r�<s���^�W�X���o�xEc���]���M��ӘךTS���9�V5��E�0}z�~�t��G�|�B��-�i�x��	PW��mѹ�+
�~h�=SZ/�Zݹ���(�r�<<A�B9%Y��kK]�ϬP���ӯSӮeB�"�����<7�yچvB��H�G����l�JE�GS�+7�q����K�o{_͞�4:���Bʠ���;�P�
�*0�]��ހ�N�0iM��B%�Ѓ#��4HF�G7�Qv��<�zCC�|�#v~��NB�f�j�&�@��Ϸ"߁������DCR��f>��ܫqkzs�:�F!0ݧ!%�w�.��wO��QMܛ`ɉ"��%X�R�"�O�LF�ow@�$�!�A1����A�d�ܦ�� ��-��G�˭��neI��z(�+���3h��X�y^�@�N�XZX���Q����E=��qj�^�(�]�9�^d�h��1W�2�Ix�M�r�( S�$���
}��V��I-F8�߻N,̟b�[���Ȓ/����M�)OP
��`b����{�%О}/����X������0��F���!�NS<�|\r��mL�)`�� �<�C�IL_n� �L&<gy����r��*~@#�ǐu1���?a��5y��/J�Cg�>�4�ڄ���n!��|��#����"�Bt�_ТhCXG�,�t�ü<kv�W���G���[[F���GI�KZA��Z?�sDp�--�n�n%�z�<T_���u[)+������e�� �����ݲ�ڇ�'iwT�ҵ��^���������������f����:z�}e�d�n�x�y,3A�9�h�o}�"������Q���I��Jqu�A�o�$�K�K�m�:0�������BՌ�n�9m��V�t�{�v!{�g����l�D��do�Z)N�K��+�z���b�D�R7˳^[��L2��j���K�iMi�]��+�NQ�P^ȳng03ȶ?�xP�����[����avsadfYyhy�oz�7���EF��=Լ-�.Y�1ʹ^*��v[��B�^���iR�}<U;��=�m��^�:�U�jqg�p�k^�pi�Ӝ�V�֕�9޷s��l8��)$�f��V��٨T�j���tc��O>�;x.!8s�B��:�=>h�-O[)���@����[[ý�vam.YX��k~ii�:�u���Ys穬�Ū9���N��a2l��k˽��訽p��lү�
��ay���������Rq竭V��ojun?{4sq>��z���fg�թ��,-&���0�P�J��ŵ�KsI���[͵Ҩ~�j)%I�Z�Ȓa��`�6�m][���`�`�p��&4/7O��4ٸ<'yy������z�2�*秛��ۧGK�����jV���i�ìI�4�����Z��2~�w�_�t#˓���tU	�$Dmd�<#�%`* ��iL�P
]���,.�a��/5	BQ�PO0�lc.P�E�'،	G�5��Ro���x�6v��.�����5ڥ�����߾}��ٴQ�z�-������+V��p�ȃ��
�#(�$,��Y�So7�ی�r�}�8uN}�6$�����S�Ex%j�y5���..7]@sۢw�$a��.4�h��t�T#˘(�FH%2�@J,--lnv)��(�Bk>�p�Q;I�9���n$��jU�;���t�@�� 06�V^�[ �
�nTe��GEV(M,�����G����/_�:X�2�$Q�Y��8�`��
��7w0,$6u�g�I/�@�jI��zC��V�[x|��D���c�
�i(?Ĵ&��� oY:V+LPłP��,�/'cb>~����طT$$��f�+�~P���Ih�T �3wN��hff��ɓ�I��d`�2�4�[F��W*s��Qf!��2���g�l�4���Ĉ�0B<E���p���0Q�9�?&�F@�l��2:\�x��raPa����SZ.�)��	D��O�_����_����]*b|SZ#�����[_3��'_m|��g�z#��ϒ�ϲP�e)�+ئ�|�)%9���N�5��қ�cL��&�
�άj���@�v���
��V�G@��9$7N*��v��߰h��uI�+�H��r�.��v$A.w���r��uQ�_Yw��k�Qk���E=^�jh��uf���j#n߾�O��6(g3���ݚ3t7w��r�fVum�L��ц6,5uO�Ç%�%���4{�;�Z0��T����D�S��q|r���?�jS.m�ȳ�)��h�qi�z
=����ο~�J�N��\�I�y�%�F�^y%)�0#*+
ҽ��$O�o�e�Z��Y˪��g��ԝK��a{O㜙����efŬ�D��Y)��b�ƍ+�˚�G�i̫���]�(K�XFo��onn��5��AKF�#�i)*��������=�~�I=���%A�\��_�ؗ�.�ܷR5�B�W�b�zd�?���q���=��]O��Y���_��%$�6�QKE���Z�zɃ�����JC�������{O7�ux@�hC3����s�3�?�O6Mj�����͛g{{���_�@/L���{ɲ�Л.Df�p&YӰ�81�i�~����8�Y9ΌG �Nt�s9!��#'#@������� &�7]w ��DF���Jd�A�׼6���|���0q��y�}��t:}QU #���1���g��I
<�l�	8�Z�`�Aj��[=0G�[�adr��#ަB�#&S;�	T&9�d)e�;� ݡ��nL���,��d"��f�������a�F��$�j��:@X��$j�k�x)ہ}�Q�a��A�z���eEh��Ўx��؅L,ޚ���Rd{�'������ c����1M;�qJ��D��edz��و���b�a��CD�(�a>O/#�>&�	8iV�Ȝ5N��#�"ʒ��(�$�o�%�HJUI`ijc)4�;��Ȕ����[��WџG���*}�:��'B��ɓ':zzܯ������� (�d*B�}�i��XP|H�-]\ѵݨ�D�7f^D?#�^4�?jn��V4�(D�D<��a2�}9�P_��3�8�@l���-.#1�@pt_E䔆�X���$~������ �Q��[c��1���_D��b��{��c�?/H�PK9N�7f�X2�g�W�\~�l���@�hq~��ʺ�u�v���JD����Y0A�@f���_Hg�l���GwE��	�h_�\�O���m�u��WkW3+#��EW���W4c�\+�[[�>����������W/^HZͤ�NjB��ٕR2[Mʝ��$ͯ:��~ki8\^YN�N������٦�Y���	N��$�.Η���ZRM�45�~R�>���q��)��G��8l���,05������q)��؞��y��dvQ�7����݃[�M"�����Baq�,��I���$O�mn.�f���/ƃ�lS�t���Ȥۖ��;k��nw�a/����K�Um��?\[\~畫��F�6i�<z������-A�s^ҕf���?"��4gNgՖ�*[razp(�uP���a334��6�z˫2��I�r�����ɸݎ)����o{��^�>o��mo��|}�R�><�j�jZ|��x����s�g���_���3�)�3�a:����s3���|�u�z:8�۷>
ڼ{KK'}K�]_0~��✶ʝ=�z�m[�|'I�^�ڙ]���O��-Yݵ��T�V�L��f�3���ͩa��������7;�c	��;��]W�4:��1��N!�0}g,�f5'���ϴ����ӿ�O���i��N�\������d�pca����������5�sf�{���\�>z`�^��7.����^+k�V��R�����T�ҡ�]�,�c�k9۰�r�d�S_�T�hq�s��V��6R�th�$�6�p,'�z� +J�["jf�f��Oh��|�C�i��$ư��pE	�8[���ʛ7o�+����F�����ly�mm����wce�NyQ���]SB�y><�z8�b �Ǆ�"12�'��@�J���Q#TQ�M�H�G1`|�?lL�4���G�AK�i�ę�I&���8o=��
��+�����$g~X/t��3��,�����i��=���c�@3X(��Iٵ2)x�����t�'����#*�kf�M�b,���na鈁?��jU�ҒӅcpТq��׮]���&�Z�J��F'�G��ȇ�;gt�v��4��D����]�NF�_�^j�2��b�al�"�f�^��i�w�����?���?��?}�y�6���������?����&A]63�$sg�Y8zl�<����}s�8���`
!�΋4+�l8��0�N�v�&Jts]_��)7��H��4�y�W$,!|e��E3#^�TG@!`�B&�$N���.�3K� 2)�ܶ����~q��&��w�E-�̛p���'��]��B64EW��a�!'7�$Pb�:�p������C�q�	�2�fvV��u\����~o�P�F����0����(� ˤ�0n�~�Rzg_|�����xf�3�g�V�G��I67Js���k���?����whjl�j�����Yi����_�:iu�|���ƺ^��O��\_[��z��#��$���a~���k��m/
��]4���̂�벭��[�iowue����'������1���:o�޽q�ҥ�?��r��-vui���]�_���Xs�X�ॲe��K�3�/��L�����dv��fu�k�k`��Yε%~I�nn�_Eǈmu�[�n���w����R����=��Ʉ�;6jZ~oh�szfn�m���+V��ﹿwd��#�E�Ly���<�=����_����r���<W�V}f���>�fm�o�.������)==�dY�+�q3�O��
�f����N�붩��ZEჂ�
�Zf�ݶ��ϓ?��?ZY�hHSN�e�����Nz'�?�����G���������qk�h��/��t�[�Վe�祂�/��CӼ����+���9<�_�7��`�`?����������?����������\��ވ�����yf�4��ݻ{�������c��2�7�j�[{C�<�e4k��ⳣ��C3I�>�$q?�t�Ҕ�����F!S$	�P���N�S_��#J3C󱂳��J��ܹs���S������4��iIr֓�T�;u��e����$ԧ��Rd�#�2�AC�h�������ȝ���L�-e����K�Ν;zЛo��M��A(r����PS/��l�QQ�1�s��̛��ȝ��<TR4 l�3�õ�5���B�֫���|ѣI��X�Hآv��N�A�G�,ܩs#Sի��Y85U�1�/�&��MkCʿ�?	'��%��%E�H�����B��%�wv���H?;R�0Va��n��ێ7ICk�^�^���j<M�vmZɮO>����~�l����{���v��坝]��5pc������SKK#]o]�]D=�,�u���1�Xp�(��&\YY�C�^P��ZZ2�nh�I��d4��0�����tL��F������$�k�D�'i�������o��y�b�<�EF��=�' :�\7��սC/x�+�D�@ģҫ��E�g�ٙ�2gRA~�(�&�k��1͈@��T�Ґ�6	#N��{E�D[�4tt��Tj��;_�ů9Ͼ9�xe��i4f�$É�qxN��k�/���}�����@��	��������W��7o��=�K:�G�w����Yƨ�!,3���H�J�]���d"˩�J*i�+�R8����2�����Կ�m�o��m�5�>nm,�Wsm�R��mL��$���>ַ7w~�ww{o�w���O(����-s�J֨�	�M鍤Zel��<zO�4������Q����2=˼ln��;��`q]�g�;���[o�f�������gG�4\Y�}z�\���G���_e��vvֲ�я�T����e܈}d�y���ޕ�9�4T��oMO��l�n�LT����O��	F���������ͷ;�����zZ�������:M�G�Ӆrzxz UV9<|o`�r�8�����.���*�l�+�����+3�4n��R���ݺJVT<v*�Js��Y�f֢�22���㣩���=3m������������ޚ��7w��t4y����x�_z'�����/�ŅGO�f�T����tv�f_cΏ_aԘI��kK��M�6����j���Z�ތ��+��1d��w��ʲa���be��2{��[�ot�f����6ӷ�~��ç��+��Ҩ;?���>XZXo啩a��e��ѕ5�ڔ����ѥ�g��O+6�l?n?{��ѐսs�,�ݕ��߼zs�Z��������7��ޭ���s��w/\Оl�{S����v��Ɔ���L��������X�DR6����i�I:\�p�y��k��&�.-x���JJ��
]+����g��#���@1�Jr�u�(���(1˼\���V���&�"���kW%s��=��ҹs�p2��XA���%�F@@����Z�Eć$ GF���3���M>t7���e$ߏq��c�)�]��lz��^��|��`.e�i�(�$;-�jJ�-j����0��&��}`4��[���[�:K�N�'�CD�{���m�"��7�Bt����n��� ��5WP�� ! �?��o�:�8/~h�PE�C}ѱ{���+χ���~h�l��R�EB�Ơj�+�^f�y�����7%�w�iv�s3��6�֖�<y��9IE?��O��?�m{�6jD?��7;��?����ߦ�Qˑ�m T�Ȍ�0@�~�u>&�,!(R�p�.//� 9�ԣ�F?��L�$jR5��xd�vrr�V�?��1x*dϟ�����^Mf��\��[@ii��k�L7fa�ы���Ү$��?t�ȼo�����ֱꎨ�	Uz]^g���G�c�4qC�@6[%����E�Lf�TB�|�BhI�#!�K� d��vэ�>�qz0S�.����2 .7_͜b�9��PJ��1���cB�W�Op9b�I�	��P���㤩�
���Is����ᗇ.���!͕�J��l,��d��<� uW�=Wk6 �"hw�D#� ��F9���ٖP��P�z�*<�e��o��C<�4	")�5�k�c�ݻ'`L��:i�ס{���;��##&�<���4Po~�O��W.^��wi�Z&���%g46(�_Y_����;��;7�D����L�RF���Zh{����&�� 1o�o��N�����S�e���=�p�d輙��z�k�/�Y}e��7o~e��Ǟ�����ys�{�����z����S+9�Q��/Za$�����/�@��%��;�Q.\�b*dd>Ņ��Ķ��>��CM�;�^׻\�9s^�V��zmY�`��=Y`���k׮ն�L�l	:�K��X��ОR�������v%��W�u,����1cZg��P���=E=7&��ր3f��R��{�'�q�{ 6-?�~fFT{|!A?��Cnk�6�⢱�f���N�b�/^a?����n���54��J����7~ro�`1\o#��xb]F��v�2q�ڀR�"��P%�	\�x�����_�����+������3�M\�s�k��]��{�?*Z���y�v��/m�f�Q(d�v��N��F�V�����"�1�4��#�C<�7nܠDKw�U��Nd5�����$��ɩ��s�$��Ϸ�!us�����#od���+�ǂ'���%^��9�D���|��c���V5	��Ț�4;;���3B���UxIu�L��4}^���"X����:�H S�4`-���b�Wc��?B�|#�*�����$��˴y�6|uBr���`�lXJ=BS��T���+�ݫ#O�
�hzq�Q�깒�z�գ:���5����ny`�q%��{���ǧ�u�+�|�лUo��V�3POv<>C��	���́P�F��w����o��w��]��nc ,����)�O=T������/�?[�Ŋ%�H(c+a�$�!�b�֕�����8��OƑ�ȫ"h�ײP qp`N}�5����rI2��l���?|����x�a e��X?"�W��Ɔ�2�a�˄��w5���r56�KO9��Ώ��X�1J��>�\�m����(�)������]J��h�3�c���͈�b�1��Q�/�N�+M��o2 �Bw��BRV_�$���6�`��m@�$#�/�_���hjj:&�:Pd�{ξA�6��3�}���_O2�$�|||�'�r�x�����{���L4��J`���ǂi��8�2@dӧ|ssS�ĬG_�
�,"Q��I0)2��i��>�۲�K��NT'�at��a�۟||�w����࿺p�+:H�q�.kb�� ���l.���j*��A�,�\+��ѠWM�G۵���t=���J�Y�����g�ե���K��v�ܹ�Arr��;��z���9�<{���}���t�����+�+g�`�#K�t�Z�rk7G�/�Y*�ta8UN���Tm��5;y��A/i7Ϧ�A/-����G��k׮�b�#_��w�����l5ۥ��u��:_��~�ٓfw��ڠ2Wo��;����#ԶE�*�b_B'K�Ų��¶���ֈіfu%='U���Vӭ����w�q������C˭��_{�k�������D���y����/���?�����Z�}�^�l�nk����2#3/�3`� ��6_��I��_�[_�ז�㻧&���~*�X��-���+^�p�fR^��N �9Oe8f����`��A[�5�����zc��gW����i�e�Y&x��/q�}��Ƚ�2ks-��6�=�ۆD!��P��?����ب�FئZ��n0��U��*k�}�����}��v�y��9狛YE��JY7�=�;��ϻ=����zcKR�#ީ��n>��{ͽū�KW�O�
�J��ҿ}��/���ꆛ�ONM�T�$7y2Ӳ�0-��������7'{_��U۝��5l�SGN4q�lg�گ���r~蕊�-�H%â�U�I}�;x�s5�ei,><<��+i��p��h������Y���8b�z@T���Y<�:lL$�9e?�d�NN�F]؏����ch�o��y��Bי�	@C62�[�(̚����nwccW3��cD�o�1�=��a�QUi���e�L�ǅ�=��n�����b��6C{Fף1�c�T���.��$rH�ull��!r�&Ismd�ب�3q�l%�鏌J��89��<-�H�A��l����*��B���*Y1�'�TVR�cč����-���B|fD'l�Gtk�|[��X�K���'��R����E�w�.X���Ҁ�03����������E�SV���Ǥ�M�l&o����}?Q˄_���N���~L�A�LZ�
}d`��,t=LP?A����|�F��;6��X�8��k7B܅>L����o~�o��6�#�&͜TvFI��p�g�y���{��Y1��}ED�D�!��F��6a>��4h�q��2?*�Lrr?�&ar�5��������~s_Kw�}oC�p�:Ҿ7�>H��!�i��>�s"�0gpJø�TC�I��$♌�e\�%��X�
f���Y��큑F���xS~��e"Nǖ�/�¬�2�7'�Nu�\�J���]��҂����:}�E���þ�t�+��������J�!g٨��_if�oNʃ�)��HNKS�������76v(�
�R	�I�S4�$�%���u����8�-�U�ꭞ�KX6>a����\)T�X5�d=|.t�h���C���k������)��\��똜r���	R�Hu�昨7nQ���m��~�0�D��1P����U+�1�E<�
B�[��i�m�<�����㍋�|Xr�
y��IV��0�A��~�Ž�W_}5m���K	m"��h�`\v�����ll�(:��@�H�7��kw��R���d���ѳgϞ�i����֮�����"� ���Hw�d��+��3n�<��@�aZK�*�=��v�&6Xyx����|�əG����7o��п����t�ؔ�\Ҝ`_���z����q`N
�tB��t֜K�A�m#b�<�vfጵU���?���;T~��H����NZ		�<}�L?�����u�à]+��>n�w$A��t���N�uy�dR\���&�%1q�v:w���8O�>�V������`��A���t\1� �ĉ��`Q0?o����?,V.V�ǔ�4�YWH�
�������J�� ��t'H�
�U�e�)�L�c��"'�!�
{�Ul6�a��|��c��Q.+�%*G���ʼ_��G
���WcR�b�FJgvq n�|3��g�䁣K��t/mll�/S�|ctx��p����&	�c[��-��1��g�YUZ�AxssSN�ܭ�?)�����a%�4�j���2�ӍIz��ғ>����/PVs��jT^܇1��m>��(�ee�+��u!��l`���sVW7^x�\���2d8�D]/��4.㈲�}%+��)j����vJ��!���&���yq�%_;��KQ�j��Jrd�3if��0��	&R	ѽ���7��_�����}����7��|�1Ł�/<h��U	������ՂD�"?n�ٍ�C�8 c\���㰭80�Ʃ�EJ�r0ەq6��L��Q�W�����S�����-����e�ҹ�8#mJ�q�U+&��m�>��A�k<s� ����}�*�d/,,��U��ō�^�/,���� d��8E��0q�=�B�JB�л�I����!�3��|6]�FJ��99����ʙ3gpl�,/����I��!�ƀ6���2;X���t�&����sʃAӉ��b�p�	�b9^7n,��^��]�ڷSv�'^�ӓ�Ė��X��r*S~`l.�v3�N�VEz&���|u��Ȍ��٬X/;����z>x�u�3CS���Vwk�����8T���Nuӫ{ͻ�������oKLd476=ٳ;�����ݝ9Ǿ���-��w��A)��:�]��N��P"��d�R�9�yWC��$yaocݦ�R�LkW��04\�	�db����g I;}�p{[k���Ѳ�u��z�o�G���=??T<7ZO�W��v9}��xzjl������_��_�,�C��n�u[����^�m{mI��0&Ώ�)���N�#Gh$�L���`qz۱7�f~�<^��|e!i�����v��l��red���
�:63~�G��ùbB�5��=�0�[�ʦ3M;�B,�7B��ck�8�$/TcWkj��饻K����S�����������#�Pg������lނUm'޹~#���*�P0A����C{뷒�L��-��������t6���'��qw�?b%ۖ��v�����|���31V٫�J+;֑��팵�d}��W������vùJ����I8���X�\�7n�]���3��Fyxm�n�T��/��fkGX�f�%�+�N�3�^��l'
'�{���snݺ�cr��q7.���Q{&;�N���~�����'�ܹ3 �tT`+^�p���9e& �H{'�p�o������G����L#|&�仙V�G�@F�E�V�Gq�lL�,>%�>E��.6���LMM�9��$Ĵvb�n�W�J�W��7G5eֈZ�9	1w�Z��C�(wpS�3�W.x�Lr�S��53ņ���#�jR-�-��'R���%}P4�[��l��*Q"�Mщ�MMM�G#��p�2�K�^Ba��٬a�=:�B�+�P��x�<�[���'�Ǹqq"�?5����	m<J�'3���-�D��ShXO�4ޝ�gGMz|qf2���W��W������F�1�v�G��VBWn?�� �?��[��sS]ec� �w��H���qJ#�q;�2�5�T#4�/3�l�xF�Wvh��p�?P�=:�o��������cް�k���H�U��#��#�F8�8�8>��h0�h���$�";
q!q����3R"&곢�5����hD�o��q>���v�e2@l��ս�@hL s�ۜ�� { �9������������p���p��q��qK��nL�e�B+,M*���ܭ��� AVeގ݁��C�`t�aր���ۊ����+�f
��0q^z�%�Fl&�E�Z�kdO�W ֙1���
y�-�FWoӄIi=*]��.�i=�ꍷ�h��W��a����qc5�o(V6���ݔI�f�q&��7eؒLPVs������ 
|x���0�{.�R掎�p}�'IF��d.��t[Kٔ�铮L`�Z�Y����rwa��.�������7ϟYp�5
V:$}�ݍ���:�F?<lt|���\cɺ�* $3̈*n�;{�,-9I�^\�LN��}ome��0�
0'zΑڷ���;���U��ѩ�v�'l��Y0�@}2t��L1����O�<�������Z�c�B��Z��)K���EMf�<��BJ\k�,�LM4
��|��`��p+@�d���u�Z'ki�[�(��>4��ON���W�1��U�9�̳t^J��r2yTÐ�Å"[�Q�n��+"2>H!9�j<Q8Pbv=1|I	ƹ�k�~����OX3������_����b�0��T�mfG��j�r�?KJ\���Ľ��	���'�<$�#���+d����f�($L ���l�j��ж����މ�R��'�VI�*V֝�P�Ѕ������7d���4��89�-����P�Rgll���eB+&�Ⴛ�� =�q^'������fLQ�O�A�
lZ<5Z*3�m�?�+������A/����_�n3l^�&d��I�d���t�`�U��nQ<>q>O�y��	\��Ce#N�W��z�At0h-B��\}:EdX�O%#?� *l2��b�_�J�8��\��/fldggo0���	G�
�K8�D�+�?1�R��B`V�Z,P�iM_Dx�Ǆ@8v�(�����wf7�2I�5�z��W��տ��/��X��j�26!=+�T�2�����\&�C�I~ �3��,u��Aj�[*2��V�3�#�b ��,�;pdM".�,!��BK�ҵS���.]���������aD��,^�X4����)D��N����h��,�h�F���&�[���.s.+A���w�"F%����q"o�l���tJ6��옢,�Q;� .��B{�L��0=���$2{�mv�1`��3��᝹�y�� Sw�'n�����:�,)%np�E_���#�&����"���[){�yf��Q��KI^�w�)�k�^�y����lFMUn0쏩�	bv�Zӧ�X$��%�ʣ���r�F��%=+����+�).9c\�S3�^�Dn�t@���N8lP�Ù��&������Z]�/,��.�d�L�
M�Z�fA,�qON��W�ys�y�=K�yv(?t��S�&���&d�z%s�������G�f����T��X�9w�ُ�[�s���N������'��?�L��?���·n|lxb&Y���k��B�hU�n�$3���;0�S�����z@�k-�����k'p|�Jfr�����s��lw;�L*�I./ݚ{�qew���9��l;���ڹby<�v�x����m��N-,<�K�򣾶�����L�J��F�qS턴�,��~��]͐���N��H	���O��GG~�9|�F��^�I��7,���v�j�\*���].�@ҽ�r�g��z��{;5ǵ�D#t7�nM��o%�6}�N�$B�?�veud�G(����s�cY��[�7�GO�wz�ח����^��r�~����JA��� ��%Ryi[�o�;���D����ce�b�림��	�ǳ�v��o9�~ж� ����F۱�~��v�?�h��`���������Ny^n4[*e��˳�D�vn<7���=��:��-�gf�s��nIM~h�������z/��ŕ��	sI�VgA�޴��'�_d�p�6A�TWx:�V�E�#��J�$� ��ر#KK��<4���Z���&cѮ�G`���b||�f�� I����*{����3�8�@���Y|� ��M�7E<[��Y���y�<�ԅt�a`��[� ��t�Ǚ^Z���JL{e���;�ԩ��!]5�:|���2�#�U4�J���n̓�Ȕ1��h�	�O�qT���k�=�<fe�-��P�1�<J;�Չ	JЧ��R�0Nt���Kr������ܘ�J@�F�8� n�F�m*]G+Y~�~k�W3PE��,{��vL���~����tt)��oh|�y�?��?~��W!�z�)l����V���J�(0w�(��D�!�^#tS}��7	3�X4y�$�M(_ Zu���Mnܥ��/�wH�K_�e9���T?������^x���&��:9W���ӝ��(�����?po��T��vco�9q}e��<��39�$���z�b�)2��('7$0.�0�29����!���i	(�]?�G�������&��2X+`��g��^��р�3�Qf4'e*��IZHG�]*����I�+&{o���ǉ��ZRޙ$����rhH�g?�q���Kviuu�L6�f�f�� ���S.(�%Y�࣋�+һz����+%�%���ǘ`���j�-��ث�m-H�A�X̛�M�HhKZIW�ػ��<�[��{R֔���}/�TF;u���[	�45�+Z��2R�8��O�x��g�~ڪ��<6 B[ն��&�����b�����~�ļ��K�)�ƙ�}��lZ���Ζ$�4$U����z}V���	eN�*zzr��΋��k�"�@;LbV3;;��~3tp_��d�juD�`C��bE�O��O�����; �����~����/�rra�w������u�n��)����ϝF��1u�F��)�����~�ҏ�������[��38XY!\`I�pl-Їv���"=<��\,Bf�)ڸLđJ1W��v]�������n���˩!��
y�Ɖ'n�x�y�ɸ�p*)B0�>-�u�_Y���@y�3�����4�ɱ�������ϧml-2&%�S���d�W^Z��o��?=-a�����Li��{%�D#�z߷Ԧ/�$�rP�c`�]e{qOFb�I��7�4��>E���(����)V._�ζH����X*h�:X�(km'�Y�|�Ƴ�����؂0Bcff&��u�,�����/bl������˥�%lQ��@��E�3�eGQ�)G���^�����}� �B?�ݤӂeR��h!���3�����	�d����bzz��$ݳ����f'~�ࢻ��Lw������1z��P�Ɠ�P2-�9�jq��`x�V�'��W�rA�zvw�T}bZ0HiC��]�t�̙3�@�'?!#���?c>V�<D�*�f���}�)� *_.r��q<���qu��f��ta ���E���q�@V'iee�����>�9�W��X}�s����;A�5@Ġ7z+�W\r/��V?ث�$m
�=] D��6����Nf�
u+@+�]�l���L ��4��+�/��j*i+81?��>���b�C��cY���nb�*u?��~c��nH��7�|����'bf�dL�o�A4jv�aS�6T>N-+>,����{���U9|X�㳨,�֑�,�J�#�z��b*�)��Lb�N`���Œր��>�f��+���)�L�C0�����g*�`49�˖]�䚑���ؙ����'UD�B��Jaem��+�Iqt�����d����g^8	��H�_�vmײ}+���o��?:�}x���`qqcokrj4����f���\ԑ�);M�`���N�
%s���+�u�*�(�Pinjs���t��Ȧ���.7ﮋ��q�^�'�N $�#d7�W��a07d���	����Y��������w������xA�
�V��;p��B�x��v<ߒ�/I]���@�{��Ń�}��E��83++#��O���f���r�j������bq$�Z�v���޵%Y���H.UN�v��q�,��_z�����C���^>]n׽�#&���l������N�k�F�7v��Ο?������/OTw'&*����^��'��-7LZXl��Ě��pT����Y�z������P���Ǉ��7����n�^l�ܞ?3�u��������N�N�i������X^��+g���me� t�b/v�L{�p��H��~�9);���OeV�vg�d����${�������r�X�
��LK#H���w9uzzl�ɟ�Y~pײj��vv8�t�4a"�s�&tB�'����~�e�]�N���"�r?hom����|�V�T�A��XYj�J���Lq��x{�.g��72^v3�ё�����S�P!w7���K�O&�8�t6�Jܳ�}�@�x��S�+��c�����n�2l�f��F�j���܃�]��as{,�z���z�T^�Z�'����;�3�;؟z]zN$F�<�@���,`�)�p�lq��R����|��8�h66���-��Mc� p�tm����ާ�DxiB���	,l����D@H��&p��������'�y������=̌����NX�h���A����={#�h�/ڄ���$1�͊i�n߾�l��R�0�ԚL������#
a~�i�: �Qy�������+W�j<}�8.HQ��WS���x}}W�<�sg�K��1���<[Lز�2w���#�.�i����bQ�R��f�����v�*V|���`����A�UϤs��#o'JY�XT(�P9��ɦ�����֮߸!؀�1�X��q7��(�m7F6�V������H��rҸ4�RW�^��L�g"]2�C�.8v���f3��
�.a�l�$��*��n��M��w�V���O_���ͦ�O�:`���NU4?�y~r.��z�	Ҳ�-|o��#]0�XS����ɵ��i1�2^ܖǊY������
��4%�u��ˑ"n���^o:� w +t�)�&-���2�Yz�7����`lt�\�դa|ljmu�N?��	_,u�)$֐���%82I�-b>�E�GI^B����^R��J�V��OjMq����
D�\ �9%$)׎b����d�"�R���f�������7�0�	�a�����QH|G���[=��X��!^E5QsHnN�2���&(��=�]�_:��~*n��I�KV#�V��������q Ai���D���w�L"��.��)s�,���~&�V�~��r��ˤ�P�6F��o�Rn"�؀j��ώ 8�(T�@	�>Зt"��e�䂈�� �d?��?� ��jf(��93�D2�v~���n5;���$[ȑ0�4�=mшEg/��O@������%�A�����ҵ�
��m���d�'�����M��ק���.�m ���Y� &{V�Pͮ=��#ǟ}672R�l屜h ߵ�!^{�~�=r䈣��3��X�퀕RV�'֪���Ռ"52���kv�~��):9�س�>69v�ر�����Z��z>�O��N���-���j�i�@���1��j�[ۏ>���;�2QIx�Z;����ӧ����AXU�&�;<�=_����ZuM��%0�/��5e!/�)o�s�F�<R��H>�c�C_����Q���SO�|�/}���p�*YàO1�b��紡����;	���ڌg	W��5k�I�zлP!7nܘ8uW�F�^z��W�N��w���]�ߨ�Ut¸r��}Fϻ� ���+f(��@�v���	�6����g~�ĳ��:�xv�zrr�Ky�ı��m><=�T�$�S��cB��v�����~L�HTy[U���DwT��LB2y��S�,u"�ɸ�3�!��1㞼9�~5�� ���ѣG!�~�mhP,�Y\\$���ɡ�_76��Vg:�Ldsaɳ��b/1w�\<M�h�p$���f[����lx�i�0B-,�C��Ƃr�ݍb�����ԕ�`�P:~�����H�2��ZŹ��Z�w��\>#�0�ɓ􁋢�(#� z4�b���W�)}0��#`���3[[��~����Ӫ2f�*K[A��*������@d2K�>�{}��>��Ӂh}�+�����;M�u�=Z�/��R�3������/|��B�,1u�H���k���L�h���t=��E�%�q�*\�pS��5h��#�ǌ��t���&��L���"\��܊{;r�S���[2J�`>"�\����Η��%�5�s�CFA3\�EL,�0-+*���DEX����X��@��%q��W��ΆgR��?6���b[j�����a(�널�)RaKx���D<-��
b3�U���NwЯFG�5��f��*��{�90L Ơ�u.I�����ߥQv� q�wy2r�\/���OįpW���kh��Ar�|2u�Mg���RNxz���8Et�'���G���;���8)�V2��ɼ�Qj���S��\�su�s+�����פ�$'�I1�d���1����,~���T
�2�ß�$1�=��qWZ?*���L�P}@G1��OE7���4�\���^�|*���k��V3�Ne�2��7�`������� �ځ��	ғ#��欉��>�Ϧ+�s7�6�����&N��NX�fR靍]��)�t�v�
9�7��#��	�w�׵�$3���B����џ���k�r�g>�G����hH[QZ��P=T�ƶ{�6��M޸zM���~��խݕ���F|�V�{�
)t._��09Ն��݃���p����~&����F������O���@��-~/�9�aF�=Q�:13��IiX�v `��_|�bM�v.�grv��0{���]����  F��0�>�baAthB	K"���*M��o,-/����ֶtQ���Ne�P��v :Ɏ�y��^��|��cl��Df�aI�vL���h�#�#?'�-$�b�J��艣��2���B��>���ʦ¶?�0���l��+�aIe��c�0ӀאJPI3��.B���2�q���]���q:N�3;;�t+f8a�x�齷�����Z�(��I���U�WV��@�8��1��S�|�Q9v�֭<K)������8�ԗ[@������Lw�PfRg}}�dL�U�3D/Z>����פ~`���5�tjܳI��D�N�<6*�K L���U��tO��Qu�W�"��御mI��F���Qع�2�Q�E���'��j7�.����Xz�R�l���i����>=�lu@צ��K��ĸ FH���[o�����@�vۥ��ttR���)���ϞO�$nN	7;��_���)\Մ?|��_��׿����9q3GQ�R�%g@��x���[��R��c�'.��	[S� �p�|��:�,�u1J����d�1z�B�0�=�!1F��7��g���We��x('$myq����[���7����.JNz���)q�WWW���Z5�F��Dڧ���m�l궗��0NHӀ�=s��j-z����?8$�:�`��J�F����������-�^�y��^�iÎٿx)7&�`�'�Đ1�߫J�@ُ� Yuo�w�鿙�i��Xgc�C��dgһ1���2�.�9՜{Y?�8�V[�C�B�JYq�^�v������������2�k�3-�	N��ak|�K�!��>�i�_�揝�~���|���I�����m�B&�
r+}�Ν�5��_��nD�i߳tُ{���$Y1�#-�h�JWr�(�9��~��ի	m�0<6,m(-�iF�235v��z_�F<6Ÿ3��S�ts���{B+_(	65�������qż���*/��Sz.+�Ѷ��rU��IY�fK�XeK�ԉ�[^v4WO�EGY�����n)*T�M�u)�4�.]���I&~�F��l�eb���#�lߑ\�4�d�x�41ןk�7>��I�_�8�"䚸.�&�Zk�f���T�ele��o����O>����V�`oy�{/� T�"�ik�]"6ל�DN�Fl�K@��lvJ[ %�ya����}�b�9>��Of���D_M�w���RR���n��c�ƆxZ��jz�RQ*��ht��O�����@!U�{�%2��G?
p���[k�:�I�Wj�=XJAӥ����b~�9��ف�f'l�3;9��=@��Y#��$��M��������fn1��������١�Z�$��?�#Ts\���z!���^�v���T���ׅ(G�s��5h�� !���3�a�b���aZ؊ ���q�r��*A0�e�OE�Ǽ������I�g}���R�y1����s�*�D�Vԣ��@ɘ�A|�x�Ӆ�V�77w9 �<8�}Bkz�鉚�$��X(VkU�7P{�����vG�%�d5E�U�t�
e�|�QK��1	C�vƞ�#�������1ϝl��"�Ĺs��qL5���
y��777���#%�qgd\����䌍A����v	��D����|�O��O�z�-m�  ː���Zs�-�&E|�׾^��3���)5�O=������X�����=F_#_��A
Q1Ï��'&#Fi^��	�ɸ�&/eǄ��Y��;d;:�?��?��׾�����G�FB�}�^"�2�&����%�&d}�.n��c�ʯ��?�A|��X�)q��m\D�jԒ�-��eړFEZ�UK�#7���0T��l�vcv	�t:I�H��Kh Ӡ��1���f �;�cr󱲑KH9��+��Ro����D��x:��Z~���r��4T��<_f0���x0@�A� �I�/e�m�  ��\���{t�/9N�s�!��r��h�=�$��4�94�M�\�r,���X;�Ն�'a8��K�F?�3?/z~;���HR!6�fE��38���qӰ���3P`�����>F�	ɾƘM-7�f�-�{|'Az��X����?8(��山�q�>21���}���Ŷgݻ���dꀕ�ҤKq{a�L���ӣ������'!vk��pk����0���p�w0�L�����=�K��pjrr<�����^O6_J��b"��,'L�N>���N+tV����l�01<2�߹������ J�4?(��"���^5̃d���*�%�0?�7[�TjJ����9�Ɋ��+Aχ�|�P�H��Zk<���6�vdV:��T��;[�+ч�6K�n�F''�������.���/�H<�qPǞH�d������/�".��K���(t[��uq����$�����Iu{�kA���,����G�V�6ۭ�[7�ΜN���j��l@��={VxՇ�陙^ʮT/^����:�L<y�*ڊ��ǾZ\Z������o���I��`�Cd��S��p_鱓Rv���v�ڝ���k�Ƶb�n�y��G���A�O����Zi�aAk�1	����	��u���,H���H���;!>�Ĳo��9��<h�ZP�v����z�0���������|b�$�~"�'�0"3fG$gd���L�j��{�6����Pz3�� �1�_��f�,T�A�S��E�tB8H	�a��`$4Ԛ�TI@����K��.Ah ��0�bBD�tFrE����Ky�*��������@�~�}G,&��e�������T��,G�����D��m�Ĳ�*���O�B�P,HQ�<5���|W`)��͆q����؊�ݓJ��LT�|A\�e���gϬ��]Y�c�_y�9x��c/�JGGVr���šò�����˵Z���6�U܎�~�[/|�s�{�w�E��t6��K)��؞Ե$�0j�Òf�(�o---R;��}�'>�����8s�ɑgh��4�\���Q���a|�>Y�
���M�r�v�jOFy/~�kO6��b������G�LC8������v�_Ù�F%_`&�q.����g+i�̳�(��G>�}�c?�S��������1�ig`]S�.��!u����:C��~K=���$oO&�T��T���@]�?�LB'0
��&.<�K����w�(a�aQ�qSiPUFB��k�b�6D~�i �@ʿqPQ�1Øe�����BSvg�7�8fz��������2J�:XG����D�ғ�A����,~z�T������E��0���kGg���28�<����ܺ�B��������l0�t����UfC�3#D�@��]h�P�0�c��"���"�f�:,<�:���6�DyR)��3�*��� X���]IB���6�";�2�� Hܗ���j(�=j^��պ]�|��iɫse+��s��.�Oh��8�v�¸2���������W�lc��jN.]�V���<�/��}����M'E��ʒ#����[�vM�S)���3�46�<�4��K.��-�q�V�@�Np��,���C|�։����-�L�މ��_Wn���,oI��b� ��:­@�|>W��B�1ʓR�����j7Rc�ăQ�����:���շ�b�1�+���w}ϻ���9rB�ޕ������͍˗/?���aN���ɤ��8~��c�k�2�ڌ�0D4'%����^��2<;�}�b��Q�rMJ�N*�*���J�dj�I�N.�_q�乲����ø���ױ��y|��J�.�4���0$f��JL?>>F�9>��7�	l���q)z�8��#"���-�ނ�ʁ� �7n�3I�n_�4�hX"0* ��Q#���<}���A�T�=F)�ό��I�+���n�4��]���C�߰$\��Լ���5�}#bl����M�}�@x|�,c'3�J�Hj�����\D����A���Z][e���jW��W� )�%��b0��*�����%FMF�ÒU�(���� �6
�Y1j�ً��.�*P���*Y-1Q�%y/�����`��.F���O�[���F%a������o~�����h��|����ˏ[M���&��	�YԌ�㲿����SO����chH@K2�(],���( C�m}q��FuN���z��rrx I�o�0������M����~���?�<�Ȉ7�f����F�01�i+�'����y������}�����NpQ���,N{$��Qi�@ٚ�l�ܘ���B��ѪzX�h=+&gf��o����*V�.(N�m��Cb��C�ǹ��'��~�^�����2���h�q�L��k:Wj��hЏ��q�	I9	V�Tt	�\+��19���H���O�+�� ��_S�s�7'щ3̬8t�'��M\K2i��0��Ԥ�|��9� ���]RKeE�3�C(0�L.
�u�cf:�b~1	8tj\f�0�CfEnq��µ���_����'=�t�2L�fØ�	/�hO<�c����4T�x�n�
	ј�t{�n:�doj���jv�v91g�����	�%7�l�3�����>ŷ�V�������3'ﮭ��2&�[0[�z�J�%����ݯg&�>�U�_ma�`�ݩ�<�K�8��nah4S��v[m��w%�,�*j�DH͓ڗ��d��^��^O� ,��S{]����Q���N`KC�L��Ð���<����z.�k��)�m^���l˹o��F��S󷊍�S)5{����٣��L���.�����g�y�R�-O�Ҕ��R%�D�cǎyk@�UI}-IH���A��sċ�0��pgC�B�8�ؖ�}�_�Ԛ��ǏKo�drgc��뵺����8U�fe̮Y��P:}�L���Z߸x����9r�̃g��_�)(�q��-�s����C�'0�L~���:�]S/�7r�(�=�^�"��/5��?���=ws��%�/�������Vh%X�a����#IA��f�7���7w�j�]�|��(~z�K ��m�[�HJs�=1���(�I$� �b�����8dɇ���ȷ~��I;���cں�	�T�`H�j��Ɔ��Ӣc�:�ܘR�Ĺ�N\��!�ح����P��q1wB@�Z�`t�>��sW�E��F��ikj�:m)]"��l �*��o��Z��*�)>�u!^�/͎�}RvQ)�9{�iyK$����)ߙuǻxڐ����/~�ō";�1fF��W͝�˰��"��#�pc�u����Go޼�X&HYd�i�U�!�gE}��Dt�NP$���X�����_~�K_�ҍ7|�A<� l�$i��f�#'!��el���dE������?�����?������ŋ�P�<��L�����0������Il��*w㖳��a����&���Z��nu#(+b����gv�ҥ��c:�R2��oɯ�]�����[ �{{�7o��5�7���!�t;e[mq�5�}ڜv�[bbb���h*�(�}��n�4�LGΈ�$ҹ!�Ùpir�� g�>��LJ���{����4�������^�z�`k��պQ��\0�7���:ڔ�P�eN��I����@�� J�pGZ'��g��!��g�L�Y��;���
����x�B��	�fS���c2/1$����t�����i��������g����Gl�W�B��<�	����*A61د .�M���N~�i2���r	�������|צQ��@n�%�'��oŽ��8�k���Q��(�˰�5^[[sӲ���7�� ���Be�U�BU�<P��Ip��P��Z�u��(��ቖ$�ڶ����$�[�{P'SSS���J8$N�FW�v����Tov��b��D",�������ӥ�yN���w�����$h��TN��V��Ԑ��z�����`�����,��b���^{���iF{	��L�¥2#���9�踢��)��j���rkqiQ�Hz~��K��#4�%�+��ׯ\'�IIWʅ����z|F2����=3��Q�v 2���Si�Ⱥ^�ԟ��B��wl�bZ��Ќ����Rk4�0�����ӧ!����;�F�q�t��Z6�1˘�[)�n�a�Мs�<�̞�s��'>a?�DiW���s��굺�i�י�ċ��^�l��S��P�]�~���5W��/>e�KIƤ�U�8���Y��",*�䳋���'($  ��m<&\q���Soak���ϵƳ�?������8�YpkV��$<��З�M����=hk�?ޚ9��{�c�N;�m�(�h.�1�]�$�Ś��N��G��Vp)���������c����-wma�!>�f�a�}yyO�9yUjw��03�;&J�@!���bgg[i�(CISZJd@�.K�T,�����%ڦrR	�^_���2Z�2�4��'��� ����0��m Cc�#3م���H�+i���
�`vgg��"ɡ!��i���9��\~0��I_Eu&����$�������Yc��RE��FB�Y?AI�I��l��_�e���'��Ò\^�@�8f2���j����Kf���Mcy9�����e�
+SLѣ�e���7���d�e1��Η)jY$���_z���]�&�㚐��2G8QL���6���>�}ag�}���]��N�73`wX��y$�y�Xي�kRf�Z��EB5JG2-��;�����b�1���F�jA��;-��|v�%fLz�)�q��0v��15�K0X�+D($0��x�(����1�2$���K0G<Dlĸ��a�qE�Čh�@� s׌O�� ǶvP����W��8� ��_���!2s/n �D��e�3����	+n}��5Z-�t�fA����/��A����o���ON@ּ�����ҩl2���yV��j%��LS.��XI����´³��w���
,|�4�e$�����$q}W2'�4İ]IC���^��q�qX%jo��q���m�oj��O�ޛ2h'�T�jK�Xusg}k&�N��Wo��;z��\�<\���;B��9���;9;S�RY������HV(���Z1_ȦS�j�����:vDZ#��K�%��A�-whr�̩���NK��7.�_��ډd*`�&�S�Cǵ&ө�mI�$%�4:�S�~h5�aR�����cQ$:_�6�k�H �`J�n�a-^y�UȈ�9�?q��.`�b_ۖZfQ@6��u �l� �:={�Q|�(C�����o��S�j��v˵$�<7Z8}�L��o�^[��tSB�4ud�V��[I�9:9q�܃?����#c�[{�ⵣ*Km�%BH���LI��]iv�8�/޺]��<�|"Y�~}��n߾==3!!�v���˾�FU�6�ju��/���{Z�z7��Q�ۚ?v����$�����b0��S$�PBˈ�G�GM�x_�q���q��޸S�uz�=q'\L�������y��F�省�L�;\�`MS~,���?���б,��l}��7����dI}�dX_��:�H�D	&x�U�'L�ʒ��(�{�1���-M"���vgҺwq��6J�U��+´�d�75��J��z�Y���`>+�>KT)����|v���:�j͞�R�H�N_���Lyq���K�����f2	M6��.	�C��`�f���U}GY�%bra�x6�~�efӱ�?1L�d)���l�&+�j�.V0�A�x�=O±ҕ(!ŭ[�0����۷��1<D%�.�d���_�v���&ȃ���cj<=�$��!"�Ϥ4L���kk�n-�"�}j���>Bx��aM�u��O�K�'a�|[�d	�ɟ��W��U��@I�|��$Q���tX
EB��ͭ��1������?���X��jKޕ�Ǵc16v��rsb�#i7 �(q����T����n&c6?�!T�1��7q��1X�t���e_z�%�KX[bV��q�-�av�^S<���^¥~�������`«Uq�LL��Y13<\֤���2�$N�'���[�vj�B�i��$b���Kk�z?w��N`x���ʩf��	;ݐx�ߏYx�8�|�Ɖ=ɘ����j(G�=�-k��_�@�����\��A𺭝��b[ᠥ< �i��[)���Y��Ѻ��;P�(��gSNB$���u���2�(д(2���4u��~&N�u$t�D=���d�ð�D�O�GqhO�p$���ܹC;�u��TQ�%}�>�QJ����>n�ٲڋ�-"D91��('�D�0�YiBn�j�3�[գ��$j�O���"�)"7;�|�7_��0i�[��{���T0Z�$b�������.l���3���m&��V����2b��z��y[�KW��ݞ�1&�5̚ɝa�+6R�~ܪ6r����I���ZY��w�{D9J���.�<��A��D�ڕ����I�ax�B�h��V
 ����V����h�NM�M�P ��@�zϗIQO��k�RIHaW�W����ٳǗ�6��+����D�D�� �c�����Xz�]~�JY�CX>��3_)I\�I�
G����W^y��[][�=p^�]f���X�s�o�����͡�q�۷n	���(���싷��E��2346�ڋn�vW����|�g?�)<iuu�4�MEٌ@<v�_C�}-,���W�~(olu
F��Z��S̐%4�p���;I������G�� ���ټ�`�o�K��=6��"n8Hk��l�?��k�cB����3�,f:�*ڝ��8Y�e>7y.^�Ȏ�,��C7��=p���������#�PڃH!�U�XZ��ϔ&�����y�a�
�
k�k�J�K�H�E8KGF�퍳F��h;v�-�CA+ے���Z�$��P�(�ÀW���K]�z	C:~�spll��3�~MG�jӍF��XT`�<\5E�)zU�s�l2D��L�a�����ОR�r�jB�p�ILBc����N�%��v�@w	5�R/�%����t�pl'����(	l���M2��ܹs��������O@���yq^:�SD{���K@3Q�s�	�n)�?���Aߎ;���M3o���EU�p�%V�^�ي�Na�~x�͋���w4�Z��s#���B8C4��Q���~�������0%�(�X/��:9�jc��8<�K��Q��,K�[�6B=I�8e�AK��<	��r��xܸG��<��~�/Ѐ:�t�e�8���Ȋ��%�h��JN��,�� &Ű�}qȂ�pn�D̓36�� f�5�f��@��}w1/'.��b/W���/b�!l%W�.q�t�����kZQ���WB� �A�h������ta�0Ā��w|H�f�&f��ށ�e	���Є"�^a,�9L�6�=�D*�ӧO�8f���5J��4	7L�b�>���g8����s@	@/uwU�2m�06��w�w�g*�4v��0y���:��{C"\�:�SRH�G
Co�|����&*��a��=K�����g�	�8-�LJ��َD�}�ѷ�~;�������P)���k��F����l����h���PƷ7ַ�\�2�H�j��J�h`(p���AΓ`V%'Jweo�u�R���%�ycB���p�۷ob+��E�<�щ@�%�:`'t�)�Z!��W��u�ED�cX�b��Ij��{����P(���_oք��rϝ;�L�|�~������Ύh��x�אַ4Z�N*���Mgr�����c�!2��t��r{�)��\ߘ��T��o+o���t�ݹ��X�ךmٽ�l���7��m�o���ugc�&���%�؉r�P*��na�)�V.��6�n�����LDS��fD[ocG�~h�Ɍ�5
E�������Z��H:c�NN出�n&/����t����6ezz�-�D@��t�7nB����A�H��]�)F�¸���F��+qGi<�A�����YDt?�Q��oh.c�I`�� l�8��Se��
!0��d��T��xd����(5B�>mi��FsRYg�����X�J�7�X�1��� ���\�-p;
�Mk��v�׊�,�����ń� �''UGx+0L���a�%.n=55�4UU*#��G@	=�;Ĩ�u&r��ŚY��(�d��R���g߹#���g1L��)��h��'[�q'0�M�B��;�ʁ��W�I@s�����-�{1�B��7E�i���ܸ���ן��W�]P8%�h6�d�1�51=���U֒��_��_�����ٳg��;�/)}Q
�]��L��B`���D٨ș^�u�v��ʘݓ�R���L*��D�0�)1��b�sڊ�b]���N��~�_�-ĺ.�?�0yx�b�/v������U�1�3�����?
�<%�����cfE��1�\SM�C�|@nޗ��H��� 4D�EqK������5��%��̊Cp�I�x�~ء���	wb�03B�����w1���uk ^i�<P�Ɨ�g���>�=�?8?�9~��D^	�6'�J���u�Zx:��m�G��PIN��kiLӕ]�T�vF�+)")��2HK�N����,��*�*t���7P'���- 1�fi5%�K
���e6�4�(G���%W�:ɇ��zvim_�7I��o�l��v�D�<J[����?�
dl\3ו		t$Ͷ�9�@hM<�'�S�I<�I	�W{]�Yq�1���=͖�@Zն�*�\�a��O[J_.��a
�&4��#bX�c��ˆd'��H������)���Yx��s'WWW����2c��0z���N�䚞;"l��Q|~ks�5;22<2�>5����P&^|�{3���6x��`I� �=gqnM9� =I�.c�����9-�J:"�0B�2J�����w;��E��B���|�ĉ����"
�P6I|#ow���0W�S���|�-�K��[o�wsss�ixv�Z��s�_�Wݠ�{���mX���q�9+.��,q�Μ9��G?�U'���Ŏ$��HO0c6f|*{���JI-��0��H��F�
fjK�,uП�Tn:��?pA��{��eM�)����[3mTXٴp�ͮP�ZKKK8��a�|���&�M��8,̚g\�$��4,b�����L�������0���;��>�sK�.���3K�o�XX%	��7Z��`��u�+k���0~җ�Y��`�{��2��'L:,F�nZ�1Z1'�6\�T���F�\ƃn�:J)�ba�����i� u���1�Ng�>�ԩS@�;�a���69]�6
�D9���P�Ց����hI���D�2]��<'n)ai���� �li�\��l�!� t���KKwԟ�P,�j��7���o|�/��"{�0�[�E�Gw,��V
\\\�<������ṳ'����i}�-e�.��3ˊV�������hø���)iOPR���q� ]��D����]��V��P���������3m: �`�΍I"�69�����>��s���۷��0����A|>��Z8J��J���e�}�#&�L���m�� {Y��)ůE�r=F{{qg'~�&7	�'Ԟ���σ��F�&��(:�ŒN���<�Mi$}�ԛ�wf�ֽ��\A.a�{�(����4puR߉��J�V��og`�A�� !�̬��HX�3d9�Nv���ǔw.D	F�p������7n���q\O�<Ij��Ps(>��d�d1V�S�9%��Ʊ�e�B�3���Ў�$��N1Az$��`����$RIVD��s,gtX�5��p�O��|��9iֽp8�c
!|U�U�߶���_98H� �������%fzc��f���
%[���;=q@�MNL�L�]f��j��.�6�.��R�.eM*�H���b/a�5��L��s����  :������^s�o�*��&] �/��|a�87�r�;��J�{�v�����5>�Z�8v7�P ���7�������|��-7ǎ;}���pj����;�\��ˊMp/i� L�ԓ�1ٴ�N���t��'�J�.z�����]��"��\Q==�$�Y8z�q�4���EB����R�v+���꩒Mm�](�ZI��@ɑ#����MO}�8���w��%edbdum���MMM�lo���#sSu���r�xa&���!ͥ����l���Bu�
��R�Q���u00?��;����Ѽ��pE�@�v��%��v�'>����ի�%�7}�\�?��dU�_K�wI��� �IC���$�1#c����k*T��`�[����OJ�U:K��t�*�s��"��؞¥�p�ZK�fz�� �X�Rd6�D�:�h��M]b����u��$�d���o_bD�_�zf��i�&��.ɘ���o,� �`\����Sf0�";7-��c�"P�_��`1����טFM��S\(I��� ���$�DL}Dh^(���Q���:tz}0Òfp���l�֭E��V�K\JV�cx]�Ĭ�1a�b�={6�����晘�)���X�cc#{{�$��E�,+��䨏�C��-����k��Y��;z�RxhRJ������|�����2Z�Ә#J��q�������J2��w�������hu]�a%�������x���0Q��Eِi��s�L������C���Í��������!��j�J	�iK�A�����u.��T�5�+"-�3`䌍����8�����?��>�����D�,�`ޛ�zQ�p�j:]�IG�s$�Ֆ2�N5j�4 Ê3�� (!�HD-%"J�x���d�����"���F�q_��a?I;
 ��&��c�ѡC��U�Yq����B2i &������p��j�]��n�� �7�0���j&z���VR/��4�5cX6�����	;&g��BB����:c�Z���0�eE��x�is�Ɵ��hQz�1&��8E4ja�2�O2K�[�AN
> Q�w /�ym��xSx덷!���<$7B��0Hi�\L�b[�r�f�_�Z5�u:'��GRb�}�?��K/�������ؔ�y��կ��E�AM���2S��r3%`��̼��۾�H�h#��5����-KD�tV��T�*�\����X.��2WI1��Ͽ����@6hߏ�=�./w5��`�	}�H�Z�_�0��<-�f�NZ�!���K��q	�8���n_뽝XRo,ݟ���#.<�իW+�����֎���Rė(�uժ5���E���t�����G �X��Ǹ@�R�0L�-A���q��;r��Rgy�&YOVw7��{I��0���i�[�2ޙ}��$�/r��R+䦂8]4~rZ�{��i�Q���I R[I.�'ܚ�txjX2g�A���TXD<4�0�[V�J4���ǏՑ*����0A����y�G�A��C��%#�!?�Q�=�)������i4��MeFih�p(2q�K<����:a)~��w޹BS��o$���ǘᔉtpы�b�$];�����1`R�3��mҒ��q�۷o� hrRzn^�rev���.��J�"-BgST�Sf�aO�<Aϐ����a�KbY0==*����sJ)Ix�<��?�區z1�Af�4��書��㧈VY��^�T�~\g��֥�5��Ct�@�Ւ�ommho�ŕ&�C���'K12�A�;�����lVf�xzz�����k3n��,R���� ��
�-$($W�S���E=8t��'���� �!�����BV�=�]�o5v�R��o��AܱV��s� ;K1�1m'C4|�R�?k,��8�܊I¬�D�Ro���o}��3���mF�D/�"��O}�ӟ���.d�a@�b��Rܝ�@j"�,�Ĥ��k�9�5u"3�*�n4!B$��x_RiY��@2;�� ��TF滖��x53!�"��d�Ѱ�#1�/ah�a|�]@��,]��Ӏٺ��kP�l����frD�J�W#���eE�p��}ӽJ_�@��wk���=� �J�M>����I�ȤWIbvz&�-�{p\���qj�	ALY�O��u4	���YxB�W�����L���^9�fdM�����р��P+LIz�KK�Wq���P�������=�-�5qq�C;�eif�����������':7<>z������������s�45b!��������̍K{��b���y9KiWN�&8�r���~8��2���'�_ߪnn�=ڱ��߹t����d�f�rފ�N�B�{�Fh=W%��� %�㻭&V{gG*�'&ǵ|I&��@��c�0�R莵�>�z�"D������Lrk�|�̈<;|�F����l�V2tl�9u�����p�<6Unuee��Ww�y��d�omK���ȹ'����-M0��B3�N��௜�>C��b6e�	�Vz!�=u;�����ȨU�L���]��v������V�����%�}8]�wz~B�&���A:F7|?�%�~B����@{�XݟPਡf���~"�����]ީm��7�Ǥppt�ޮ6v���N{?LyN��f�����zF4��ˈ|1�i>���Iz��*ef��+а�gnn#�WpN��)�gf&vw%��9�~�v����_��Bk�y�N�`�s����"�Tӄ�寧O�ƐX�I?��:�E	�z�!:2@�:�ipq6>���ǳ�MH��N�zx¿�V3� J�B�Ҡ���؊y��<�R�j�ZǏ+��,���ã82l�I	h��y���d�d1`-��X@� �p�d��6��S�c�5}�˒������( #~f
ף�5��<G�q�Ү,�9,1��c�=t�t����jv�*�͖֚��\ժ��Qˁ�	���$��QMEC����)�VN�d�����zG:���0hoܸ�i��q�Y����|\.ั��'���?��8� `�J��Zm�J�LV��(lֽr����3�/�ƛ,�\�B�'��t�_������τ�$�e�'ޤ��8�y|��o���k�7Cg+�G6]O�^���srw��i}�ӿ����be�,����}���1yx~L�o(��ǃ��lN�
z
�-�v��p�c�x��˘�'�y�9��jK�gng�`�e��}��`�T���<����+����7��,����{��طܗ�ʬ�ꪮ*��n6E-J�Ʊ��)H,�����Ր��"�o� Az0�b@@�%yF��h$6[d���-k�=2c������FU�h�##��ￜ��;�9�!���M��9�$d�q#�޾�<�Ϣ��٢��r�Ѝs4���4�H_AN�Hr*~�}R����W��x&�q���m�s�����en8
,-�+�3����+,�f�y���}���3N�2��MI�M�E�K�V��H9~�^�
��'�!�	߄�Ǉ�b4ⷷ����TH��k����ޞdM�bC��q�K,`��d�̜�3O�6�SB�~�R��+o�z���T�_��W����v��E!�b�k�n~N��$Ϭ.ز�o�2:��HR��T�����pј�շً�
q! ��@������k�aW
� ;��k�)eq�![O��k��v��0��5�)����V�`E�ܹ�[��G��IMn��:�k�ؓ�7VP�2>���~f=i�9FZ��i�wT]���I���0W�m �|��e��'?��?�X��!k}E��d�!�_�K�={�y�cOCW,F��ܤeEU���6��Rk7��وq(l!�+�Kܼ5�9��h�.Faag��\z����_�]�(_D��٣�vRJ�Ϝ|� �h�eI�}��?��Y^_��_�����÷�z�O��5�a�oo?ai-�)��ʐ�@�?�D/)�n��K-�6s=ْ�ڵJ�^g=m�P��g/��V�&l��L�i�� kcc�����oݺE�P�A4�������p��;�k�ɗ�o��_����������"�9
�g̔޻����C���yc�)�XA�!���*ޝ'�m6��_����o�1�h(���ƍ�믿NX�dy����4���=--ĳ`�'qL,�'4��!Ƣm)@!�c�����.�o�M��D�ߣ�c���R�6[�NK�Sj��|(�	����&	�u�_�t	���lnnP�c��f�=O���gΜam5�*����%ݥQ�0DHB8�l!�;@��7��?��?9P9��L}O�0�l�(ؗ�_��_����������>~�-��%!:��C�%t�-��Tt�I�0�|`����[یD|F֚����(�i��D�����Bo&,��"�����������L茴����o����plH�����悚:�^�5R���X�6ך�u�t��h���`T������Im��j�U=�+F����I�6�����ؤ{/���h�j>�t��y������ ��|t�z֑�͸�O'���Ңm��Q�-Y��iw�RN�9�����Y�c6KӬ�E�N�l�JQ+H��j���~�����H8��4b�,�-=h#����nn?x:M�+��i�	#����orʋC#�Y����F��%�#�`�] }b�E.���y?za0M�u�<��F�7	��}L2�^�,�4�Ñ�wOF��j)�/�w_ZO�'^��8o�ay�N��\��4�j�pl��}���O�K�p��-�9��l�m<xt;�F��K������4���fz������!���Ʒ�w�7������8h���N�Z8]G�e�RXLL�Em�${�^.���ˍjxW.����zvk���0+���!�X e�+��@X)�o�D�����nr�|���B�Q����� ��=�'n��v�8�ů~�t<l..��w�Z��Ʊh�9�`�Mp�kR=�:s�P\A�^Љ�\�\L�/_��������?=�y�����{"1�W^�
���ݏ1��������������b����|�IU�vd+Ԧ��eO�Ė_�T��t���I2��@�k��	=s���>������o{�ͷV�˦YJ��Te��5?Y�~9������K# ��'b�_Y]��F���?��:v��q�����;{G�B6A
�bO��s^���rVi�|썄j�F�c���yQ��4y=W�|���?�?6��%��]�mc#6[m�h�$��������3[�^1��qX��0���O��ǻK�������+�~{�P��8�+|L���!YxH����x���Z��j�5��h�y����(����`&Q�s�҃Q-ml��kB��5
���pԂF{��ȼ���>��H���a�O|eO~��r�"ȩ#S]�h"y���D�TH�;;���i�ΝPc��DIF��hځ{��.��x|�	�O� :��,rde���.F���Z�W��ϟgy=�r�Z�s�X^<�.Ht2���t�B�i����\�5����J��oyY����ט�!�g�,�9��I���}����f��y��۹���ss퓓�o
%o�\�+k�h�4-�K�r@b�?z��t!�7�g7`�6���� ȲzȰg6�Ǔ������f�^�ݕ��Տ��O��������1אM�󶼸��ڨջ�f���?_��6j�+�ƺa�;Z�R>>�n�$3�-��M���Y?C�X�8#��4�S�n޼M�fs^�d#|8������Geh=+�c�Q:K�d�,>��w��W��_��Z+�'ʣ��KU��X����0(��Nh������8��o���3��0��ȏ��� ���G�n�&���t��9bԽ����s��g_*(�Fb���bP_�|�r��Z���TS��:�Hm�Ƕ�xe]F<���DW��6��/�N�b�ӌ1����ID��}���Y�i����%���X��m���.	İ�ü��Ѧ�MJ����~M�����Tcz�$J�A�$���:��Q^�b�I	��j�b��B���0A�+��o�zF�ό0%�Z�W>W��<����	>HRgd� 7D*�:L
I���`Q=�g�aH"�,��c�4B���9v9�"��ص�KR�O-B����{I�P=sl2#aQWac���?z�{wukE�ki��G���ּl?>�̤G_迊^���hq+dk���5����P�A��B0_�ҵa�a�3��g�'h�3@38rS#a��P��XO�Z�i��<�����cX����ɕ+W��-���95
�S$�6����q���o|���ܺU��_�j4���O���[�?�#< �4�h���<L�'}���'��ٛF��~��lv�f�mFU��O^y����&6Ͻm���tLZ,l�d,]�?��P���f<���s۽��<k�$�/����x�חW���O}|fkk9(ݸqceuA�����k_붤�����	Vp�|�xp��'���ΎY�C%��Q�=q��bvg��}�V�8˫��3��i!Kb�Ju�����m�W5Z�BUqE߼!���T(׷;��������kHb8vZ�%���( ��uѩ`$�Ĝ����~�#���a$����`�I`uc�q���I�[ܹs����!c ��`�p��}��Ga��sܸq'���� ~�������7>��cc3�h�aP��"��c��{����! ��`�Ѭ �q������x��e� �������O��S�ĄP���S��^�ʺ?�RK��z�K�.1>�(#�>�S� T0,��M�WS�`���ט��������71­���\�qp*�H�1�ꔲ��GK4�)2�2����/|N��/o�f�)�h;���C�ә�_������Y=z���]XYk+Z�R����Ĉ�%g��[��d��G}���������x��`L/ �Yz�ײ(�ˑ����vI���t,�L,f�yW���&����S�l��T
������ܙ���k�
`-�.���|p��}<;{�s�(3��	+L�����]��6ʬ�Рk����i�u3��9e�q,�l� q�s9ϖz�Z��� ��}B���;ѡ}�|�R�H�0N���.�v%��AxO^��&���߱���v��K����$�a[-?g�bS5$���c�j됫���5�lM�7S�\�=�p�>�뜆 %���W�FXNJ�Fb3�GC���(}6l��Hg���͸ߌ�N��6?N���t���"���[X�ʇg%#�m�����̽���Ķ�>S�s�x�R:	��t��`��4��x�n�� �7_\����#�m*0
�ʏ��9�e$�Q�S�ќ��?ϯ�+�q�����R�
MY}�+?�Lg����{�]ڒ@����0\]Z�㢠��^<���iR�W XOF�f���^!,7���!;4=(F�5#�"�5������6~�3��ʓh�9��X3YB2��߇i*z��Y�u��~���^m�p��٫IoEs���4�޽�-�ۇ=�b����G������^i梅�d��a�1`f�i���0��\N�"�3��aeyi���W�^�k��F�ks��9���Qw:I��nn�D3��y��J�>�=�<R⸭<K�ǀ�V�6.����_��w���Az��W_mE�{���5�믿n�$;�{n�ŷ�z��ׄ���Xtv���Ví�Y
��x�\\�/à?�Z�O�ž�s�B9!��M�Rb�i���ũ\�(�zw���:�#�3�bR�����onnV�6�oƽ������#���_|��~n�Q�jc��P�%�FX.�]�%�g��\L��l�9+41t���P�8P�,x@|�IT>$���bE*����t JL<@����`0�{�.G�R� Q��Fw8�3�O�P���	��wcK^Ef����,J�H�T�*NR%np	L�"8�*��p#�W�P�ʏ��jr���o�&{Vҿ�`����6��Ԗ�����ڗ,���J�Z��
W���>
��`����䴏;A*� T`j4���Gl��KAk&J����:���/���'�h�*my�V�v�A|��:i�lV+un��Ƕ������������7�9���r��	�چ\�&����ί�ʯ0�/�R� P[�� ��l@D߿h�����t�<S!K%��	&�q�k�-y�w����E�q����C�����l�S�(�8�V��q���RHUE0�������N��_�Z�3��kvP�d4(Yf��1M�S
R"�]��G��|Έu��yZd6�Zf2�EC~��:W~��27gҷ��:��O���lu��
x��}0����G��f?�NKD3�����03���EH�n�͜�㺤O��`E����xf��0�κ��|����e��x[	eSɊ��Y3Pc+'��bi�u�QY�|e�a1.G-5��L��4��2�O��\5
+�ܿ��ɌR���!
�找]�%|�ڐ0sP�!�ҘS�k��㝧��4��p��!>�PX�B�-$�*���1��'�ؘ��8Ҟ�W�a1s�~���<N�3E(��˿|饗���!����߽�����}*�.|�K_j�|�a�έlI��H��65p� ���2�M&Ǧ���I����9HAb�Mć~x�hz"+���/���2x�2���2t9hz�s���.�z]x�M)��s!�#ϭh�xz��X�P`�C)���2S��I�r/�x�}���|�L���������͛b[,,����(ץWiM
��������M�C׽��r�gS������)��	�����_�uǌ��<���̯lH��;o����Qc�\W!�ꜰ��t��0�?9Zބ����M�hF�P�Z�@�Jg��	�Db���Wʂ� ���IQX]z�������Z����'���}�!d�D��'�8�D���z��w���`?%�nkk�!˩�i�FV�
>d���pw�ZlLY�v�C�P�R�ѷ�:x�42A@3aJ�hKK��qƣF;e+�[|@��X+�O�����QѝF�b#�iWs@�@�����)����0�V�4o�=®`F��xe�dЫA*
�WJ*6|s�0(�P�ڲ����\uLʑ$V�'ЍKC!����S��c�jPr�"�����m�
Æ ���X,�	�TSS��1��9MW��b��cT����|��K�mI�0�`��`�@����3�񬯯�cu���3���Il��-!�?��������g�O��+X���}a	.��tIO��2��W'�)���+~)�D�Ę�/�4�+�ya<R��2f������N>�~.�����)%b&�མ��&X<���J1���8L�v�zH�h��Mc)a��%4q��T"��Pr��y0��,Vb��&�mpL���f�/�Lbc�cN5�5�~,���nI����V`�5�ǹ�� ���u§�2�L�;k<��ytNA��������Բ~�t���ۧd&�S���Fs�s�3wG�vu5FAN�c��Ӊ�I��v:CA�=��6�����\�8[W9T�	�tQz����q����r���)�������^���d����V&�\���B.��X&�غ'^�NEhq������X�f��G��r�T)W�my<ѻ���u�>�L#kٝT+O�GVMҏ������G���߈�!/�=��ǲ�R�_9���>�7@ '���)z*�����ٳO���~��<{f<�/MDʆ"1��8�ǉ譧�����@i�q����/��m�y���x:N䄰�1�n�4×����9i��5<G`|2�����a��t:9���)c�p��7/�x���@
��>n�1>��̻Lf�Z���p�&ʷ����
�0�i�ʅbI-�i�㑒�J��h8��ǕJ�������9/��Dv�ז~�I��c�:��=����%�,
���x���Q�ټ�}9�����8�L&{�̋�ƹ���������c�[����"�<����\\O'��(�%�����iΓ��X=���D����K�	��j�QÞ��iYs*U�/�D�I�s����P�}}�M�ӵQϟ I�s���aG��K����n��f]i�~�;��%?F����q�֬,W�y!��T�7������/cp�j,B�*�*�m�+t��0i�@}����{�\�%��֟M�1dKVmwd�.	�6�D�s�ѣ�.xi�.�}��
�՚��(g(LY���qS|����1)���4Ϩ��J%���w�q�3�W^�PY�G����9t����������=dysϙ��|> +�H��Q���As�ޣ��0?����X�Ag��2�
PИ���8��0B��0��J�q �O���$�@��($�J�_c�,��I�M�-�<<�%5�Fi��(�R��"���XkM����?���Q�J�v�9���_���W/AQ@>T�R�x��Q�M.4&��+�7��~c����s�C����	+j�DX�K>�Tu{nooc�u/��:A�NhHx6`J������w�}���G#RRbF�������������2C�fb�2�K�A�V��Ŵ4XF�zJ'�#��G#����=C���Cp�]F��A���Jt.Φ�6H��0Q��? <[I�<[t�r&�
h�E�;'�����M�Y΀s��"�K�����f�̯N��pu��R��|u��J���J�.d�'�T�܂Xƃ�6	M�i<CE�S�wP̛aD�����𩚛QtA�=�B��.q�1�N���̥�!eq�:������]]]��@J3�s�NA�;cj$���{]���,��)�i�y,�ո�����h�6���B??�s)F�N䜔�b]�P�����s�(3��u��_)nM֎�hf��>*���W���v��_�e��-؋a��4�S!��ׇey˦��b$p>6 >6�#x��
p��֖������.���V�3x�;^X͚뫴���Kl3֙�5�۴�nFK��&���u��D��}�3:�L��K��촥��Ȑ��W���噫v%��$����(A�NW˻*����F��ҥ*��"pɐO�9���%s/�C�H��|���"ZP���@�{��u�y׮];J���ٍ5�?k^딇b�J�/�g�o�+-�fCf���H%c?�D$͔;YVE�S:�q���4	���O�SV>���� \�x�G#�d��$�i�,�#�yc���3�(/4i̘���o�Z���Ip��z�lg�o�~��![O�C@8BG �&mL�16�H�\�~ߔ�^��	V�@��2U�B���	'��3�vt���d]ϙ-��F���U��777q)r�q��ё@����% 6��\bGx���l�dù`yb�ꐵ�ˍʛ^��Cdcm�&����P����c�<ܺu��S@�Q7��B&�1�ee36&���=:S�󝏢���gϞ9::fԂabFf���64��^X�T(m4IĜc�\�O��Cq>ݹs��פ�0�m�S�k��k� �~�7~��W,j�*�	E����&�\��	��S��c�PM2����A�L`�Ÿ	�|$�%!mj�i�sI���@���$����٥�s�qd ��{}��ЧN�������T��ل'R}�$Iވ0�{�p<T�f���)�K,�lէ��3��]͌?���0y	8X1V���M�w!�Rg��7�sJ����Y���>%G�����s�=��n�-����3Iu���p��Y6������_\u-��y� ߽foj>��r{��clI����3���%����e�+��Lw��{6Nd)���f*���y�j�|����� *������L��iC ��u��2}R\��^����It�:��~FJ��UY�GMO����K2L���BF���%���ona�p���l��&ҵ��.�sA;�XT�9��C�T�A��s�l�J�_�惹�ݜ&Ikh,I�Ѕ�4_�y���Ѩ��-�h0-?|���p�D\���k ;X�30����\���^�k,����� �zǒ�0�{�ϟt`�;G��r�֮��^�Q�V'��q{=M*a`�6�����oO�1�o8����S�������k/O�����IP-{{��I�)l�yF�g���ؒt=��\P�j�J�T�7�r�K8/�D�7o
=}�g-���	���J>dJdѾ�i|3�gf��<wx$r��+��B UuI�5&�����d��ǥ�8G��^�����K/� ��'ݠT�t��B}~�Q+�e�:>nw6�Wˠ A�Su�&}��a��x`X����a�g��4J�(��
�B��Fi�^[x)M4�ǐcy,C�KF� 8M(���NF]]�n�O�y|�n�,��
��R�8{�zu���B�����<h4��`���G�v�c�&�S��4�%!P��z�b��Q��8�S��lX4��xc\�~8�c��.�p�F@��N�\*�\��R�2o��9Ciy��~�6e�)�a���g�V�Ơ.���V�ҝp<��a& %�,..01����S��,�-�d���N(B�� ��LxZgl�F�b�c�Mz�|K�ua��LBj.�H�Ѩ�5;$b��6�#m<�0�_�_��ZL�E�F�w�G�C��꫱��c���|��$�	c�_���ﯭ��|G��@h�ON��%��uL���$�担���`4��o}s��:�uu��O�>f��T*�Z}�:��q;O@ (�"�&:A�[J�n����S5U�,H?>�C2+�0��b ���J������ +z��pINc�m��Y,)�跆��[�N���V	g����+����9@ϲ:Dbݺe͋�-͊Wn*n�$�2�[�9+	_l�qJ�6�%-��,��^sQ�̺�xG�gm@鐨:2l���e%M���y�[G�Z��(�4kH��9�u8�
y�h\��zݞ��6F�yfa�7C����pm�^�ގP�yu��ܤ�Q[g{#�g����76��4���g�Ĝ�h���YN?"_�6���YB�߃�H��(
G�Y�,�b_�g��Ҕ'��څx6\yo7��t��ʍ��`s!�K��e��0�����q<*��p�ۂ����")#s��� ��'�ϟ��bəMuEͿ�q�=��<�2ɒ"=p��(���0��U����%�)�n2t#���Vl5�h�juر�O��y.lq~��H������O/]�pa	����
�-9ɚ��t��� _T��/��\��Y���HI��vS��@K��!5����,�+_YX���Wj��dV�����o��EE<�������S\����l�ӏ"\���0Hd�~W�h�X![����l�F�s�9�>��w��������Gcq�<��yG� ͂rV�|htge�޽`sc��؂�.�oW���ɤ���*wb*	1�=?��-����1���Ⱦ$P^�i�m�o�$m?��Vw��aW�n� |E��ĸi1��%��/l]�<R&�#��l���).5�$)��ų��}��6�nc�K��]��Ƞp��1h��L��?����wM����pY:3�'y$fb���NF�p����{��X��FW���������k�0�*g�n�ss��L�u�P�5bDT*gt�:b��ŀ�1���%����q
����̰7�8\Ȼ���� ��7�-�Ry�����F��~�S͚P�0�C���LZO+O��81���E�t,�'8ч���Ff1��D�K�p�ɿ|��6k0[�lyxF��ŋ��fS�"$LN�|��
LHV����P,w`�.�	/��z�;J�[��X|�ڵ���������H*in	u��q���7��@��.Co��1�ܰ��t5�_lTց69�'��l�F<���b�qd�5�ќi�v���Ad��ڮr�����I�G��v�K��Ʀ�}�6}���F�i��I�8@l.I;�8L�wXq@����V�'�鮦}blrg��%�e�Vu�d�ft�9o���x����qփ$�pwYh�r�IF����P�z6����Y�8Xwi�մ(ߜ�3���s��j��(rB�������J-�aP�s�X�L^��,��s8'.�#�%�=�rR=���+��B�(���\p���}^�g֑ff�@�;���OʝB!?����M�{��::��Ps.`!�������B�c%��,���2::������	�(�
eQ�jq���@����� |ۍ�Ӫ~�ʜ�_�J"dt���݃���SM ��%����CS�J�$qR"e�����$ΚJ�V����1���z<na�"!A��K~��tp������/|���Qn�v�O��76E��)�+.�[������+ ��b�Qϋ�Sp�Q2}�P*N¬3�K/�49�՜�{��Z�<�,�gϟ�����J��5�J�~�ܹ�ߖi/�����ʲ����Z�����Zo��5�>+N�Ã�/'^��H?�������O .!?����W��qD$�����I��.ǳ�J�POKj�i4�L�M�_S\*o�X�����N���R �铑?������[��������ｇ%f'�He���?f7�/^�$P.\zqڀ�I�tYR���+���@�?�qC�"�7�yg%I���_~�`in��m��Ĭ�� �D&Nܹ��Ƶ��4?���
!t��L�z��_a��A���F�Q��V�|h���������_�nܸ1�sO�Փj�R��?���_�e�4�}r��R�8��bq����A�������ڙ����  ��IDAT�Ӈ:�|^7����q�q��K�Ov���-M-���P�����+�JfQ�0@C�N �"}ss�>i~��9=d8V�	�
>a�N�$�e���H!��5��;0�6}��&~!��/~���ߔ4|N��d�t�3\x��#�ͩ(0f��5E�6�"m�D�DYsI{�H�Oocc;��~�"�����	1�]���I�7��Kr��T;p'�?d��U�1��2L�޹sM΂(���p ���V�Z/F��l���(iU"m1��nn~m1��L�$~B��T<�+�$@r���^L�{�D�7��|�%ي�>��W1��Q��,c�j,�ݻw�+��t�.�\.�*SMj:�t�T�����&��h�����˿��Pj�N��Y�����(�#M�''���o]�P���a�x�&9�EiA�!���T+0Xy�.�9��e�^��\.���<u�1CF���m6�I�MI1=��������c���M�f;#��0�X(�,�1��qVf[۠-@��z}^1����5�2ɷ̌4M0l�7{�M��فT���6dJ��C�0..��[��͢"b/f��J�R#BǪp�s1���}�h�ۜ9|$��n�,��H=gT��A�̌�ų�
�+��[2�V�6�g�u�u�8����u�"�lKM�A�@ʒ��sw��������&���ɟ�o&f�{]5	b^�B@ȆF	^��������(��tk���:��-i�_g��ިs��ߥ�B��b]���`���s��\����jSC���!�a�h��q��x)����3��8��J�J�����^�E�������)��\����gyr2�~CV��xgtƳ,�S`G����� �j'�1�܄��hbcQ����J��T�Ad`�W�\)�n��fu���q_�c�q��'6�, z �_{�m��x��a�z衆��(e����ؾ7�Y�ZKv����������
,���H�m $��q$�^��U`�yQ~q�����(�EE�j4�׬?V�_"��4�H�~���EV%�#��J������D��'Z�g�H5��,K��U�A��l~�쭙��#����l���:?�3?���fҰ:�����,�dj����ss��H���Xj��&�i~��6&�g��nݺ���{�T���L��.��]*2._�0S2����|��w~��~˼�6�9j�{x|����%��r��q�j�g�y�tL3�<\ZR��\��d�#[8��E&B׾��,��T�f�b`�����/��H�&�9=�a��
�`3�XN,s�x�X���[�8x��i�P�a�	����������ƻD���� ��)V����Ҡg��-Ji422?_��į��6t�P�-�����g^c���&�������)v�I�BL�a�Gת@���|-�I޽�b��S�1����sƨ^, 'Π"a�.�O(9� #U�`n��Z` R�% t�<�BZ�jg2s�����<�O�u�DϥԼ�5�r��
�{F���;d~~��e��K�Lz��ѷ/�~jb�+3�<�T�/�y&��Ʒ��m�u��Ź#�J)_�N�=nH)�֪F�Fcr���1ul9C�"���r�1.���.�� ���c��tw\�N�j.M�nݺ���#G�� הal�o~�F��A5@����� ���-X��S����S�i�,1�.�������J�ڌ-��Sù���@�0�Y�&\e�{�l���DMz.W?�ME��>$���Z��&�'Y^W���8O���v}N)xϦs���U��g�y�V�جY��K�{&��OX���*���C�iU�)n>A�T�+�J� ccf��b ����3��Q�m\�E5���#�\I$LO�%���|�h����n��z�7rp@���%���`\ �Aۆ���a�a��Q?�T�da��rOӘ����D��qG��j��V���.Uʩg`��6���J��T��S�H:_�d:;�EK<Q�������/J����Vp�����ݺ5�ldK��K�.[�s��~k��M�\[[�~���q�-<�}]O�
n�A.�*�8��B�7�������d:��Ø5i\��M>��iD�;�r���-���M��d,�[��oma	�<�H���&�|��e�*���}�w�[-<V�2�KD�$4��a!_0�ʐR�&sE�~nk����K�j���2	U4DA�Ta,�(4	w0&V*�$��>4�+B4��0"#�:��~�p�Ţ��3.��;�9Sί,���ݟ����Z
fЕ,��|q�P���f��B�H=�^y�Ճ�b6V�m~(�KЋ�i����L���~��G:��4�z�����ˋ�!����y颩��c?�PW�������;<ܑю��ިs �E�'���6�+<�W�^:I�T�U �*�x�v�����	$u/�ƅә��Em:D��3��=��A��b���)�ZH�[���A����E�c��j_yqH@/�C�%����iIﰋ�y�3��d��P#�@]ʸ�i��.���xa"�I��y�� ���Q��I��Lc�袾MX^�� L8�0Q���ҁ�2f�@X^��89d�au�/��f��r�2����mt#�#��'����W3�f��"zE\8¸Y��Jv%֯q��1�3O�Ǚ�"�Y�ؖAlĉ-��C�Z�����Mt¼|X�� �[pI��7�:܉堂� �"˝�q{��R����k�B���؍����,(
=���8R���	gϞ��M#6�J���K�����0��Ć�2��ٹ���Q/2Pn���Z�0��.=:Ta��RJ�DL/$	-a>F����p���O��O���/��߇Q�y��������o�d��AS`b?���j�L7����/��p/<i�u���g���`H���5F�gi]�~��.(�/���e��YF޳}-��l]oG�6�)<�)�..���1:����j�e>����	���m��iY���S��8|FO��F�y�-2���0'��ݼy�ut��k�p�+���/!#+K����'�C�&�?�}(O��L����j�]8;�|Tڔ�+�b�3���7�.�1���Rj�O�86�`e�l�<4kh��F̪��9�؅ܦF��$FS�H�f!CE���$���Pj��TD? ���f=4����]<��w�}�o�a�^1"|C���G{�׊:��~�����C�;�@k0�����GS�P�22�hN�K�JM��^�a��������R}�!�Se�&�M��>+U%U"A��&�K�4j�V�
�J8��IF}y�O:|H���r�*t����Ӝ׷�
�R�Q����[�<�$GA�A�O�b��HΞ;�u�چZ����o�HVͮt�\{�e.�x�+J��84�ٗoK٩'��-�
L;�? ߕ$���b�R�;�'�d�$�|�kֹ�X'hҌ��(�甎_�?�ĝ��T�ؓ��G�O��0v�_a0h �D׎%�Z������߾���~qeS���(�"/�X�'>�ۨ���^� ���L�ZŨ�GT���lj�d��
��Ο?����r�1^�KϱȆ6�l�M�b�`����"PR���.��b��޴�ɇ�b3��Q�`��AT���/�)$t0Hx��N_ �R +��XGn<��JXV�j#&�(/W�><�R�%Z�Ʊ1ˇB���"�,�p��>��KtEX����T<L(kO_ˢ��@&3������=fY�� �.n6���t�M��2Q�rU�d�����2�����B�!)�n6�;��>����A���^8���,a�!2������*O&6�%��>�*z��tؐ�J�XKB����(�E#k����a���ˀ�DW��-�q'�$ .�޷̴��FHD��X�8�0��޺uv������M���+�㓒����_|�E\�U����G�᩿���鰙�^��iǔb�s�T`�?*uү��۷ ?C��/e�
f��g�9�=c]�� �eE���R5(�μPPf&lB�9���m��9�(����C�8�T��-)p#� �3Ta����MsK3k{���TR:Ӑ �Mf��s_�`2�7w�8�9u��ܓ��\���%6q䂊�g�Jȃ*%�1Ҹs�O4[=`[���� �N�bv��|���zp	����wj�^t�ғ�@5F�lI�4Sr�{q8�D����8/�0��O��<��l�~|��JS���FiX��Uj�j����(L�i4��k���s�g,��jɣE���<y$9�W�����)5��h�%�F�a+W�JY�i���[_^���w���d2|��7�{'m`߅有��$<&$���]?����Ρ餽��0M+�h0��y����K^��9P�RNmY������[ģ	i���ݽG��;w��ܹ�Bh�,@j��t{������tttx$-Me*E��P�z�ܨ���ڨ+�����|��;�A�4CPH����'+ǭ��$�?����N&PM���ރ�R}ee-4���ɞ�^Q̑,ʯ�$�BEO4S3{������ջt�n,�O��R���qcn���B�XO����Pj���K�^��͛�j�P��	���bڛ^�q}0����Q�L��_�����Īy6MV��������ƕb����N^��8�R��4L{���5+o}�k?��{ߟ��aZ�'x�r�O����N��4J����d�ʒYY*�Յ��}<�yr�������BWu��R-�f���3��j�R�Ђ�������D	l�M�U���	,�"���q�G�[�0֯ѹ5���chB@li@:hI�.�F���d��UU��`L�����r�L�����3J������E&�k8�E�?�Z�*����2�2 ��b���bԨ�͊%\�.r�:�H�[��{M�K8�5�L>�s`�\ZDb�<s��(�y�"q���@$�)}l8zP��2���uu��A p�tnY�|��ƣ7W���><<⍤�k���؝��-�x����u�Z�x����{��!>��W~��_�S�y��'��yI<Nci�M��nT�r[�ڵk��k����+���<�����+��O��"���o�g��!N�;��}W�C��M?��#,��/�̄Hz:I4H;��с,�:G�o�Ч�#������ݻ�h0��*W�\�]t������������jH�]B��V��^�廟�ޗ����9g�#Q�Vb��Oǰjm"0�������<_�Ls�%p�ƺ�hW��]�M3CV���n����0�Tsn0~�̴��Eu���x_�������*#�f����p���E�&bfY�"�Yc\�o�W:s�UNI�g>��+�OT��7�pO�y�¤����l5E-�a��(��cIJ�.�J4H��4��2;g<�r�������S��J1b;w]�Dږì,dE����1�;s���gU�*Mp%<ImsS}x}���D�h�a�i�U�f�z��3^>YT�1�B1''�z �z�#����0�a\m��3�v:�_�uк}����J"�Ւ~S�X�V8+�pNm������G;�[_�,���$�|�yA��Z����4�,{0��żT����\��Y=:x*LN=�=�%�N2b6�H��7��/_�lΝ�����bE浆˕p�"���iMul�q�@�ݻw_�u�x���ZSҒ�G�ڮ�--|A�kQ�&s��N��<k3=����\h2���B`֑�"!�]\d
�ښ���cһq��|CB���Q��5T{2'�DZ��l�'Z�g�NEjx����-�
|�k�&>Q)��㖤�YYŬ�����ʻ����~�w�Xr��uٍSY�6������#�Z�wd��T��:��se"j ��L��w ���JI�/�0ǵ&�4��qڸ���s<��ȡJ�T`;�p�Q����6b� a�"!�A��a;[@ 0ÃYV#��|
f@���K2�P��+L*]�$޻w� �=+�]p�Q�O�`�/��kꕨVKP���%nD��aD�5R�.%�����2�	a|2����X8>��\��	��j0R�N�0-�o�������p��=�KC�ə������;���#L&�!�]�lX(H��4�-<O��R5m���ݿ��>+x
l-6w��1�ۿ��o��ʭ�w15%F�3.N_ 9mf^5�Җ|�[�ܰ��9O�Fe;�.��t� oi�i�������ۯx��&�z�3�B؁ �}Y�X��ծ���y`�t�֭+W�ܹsgee��y�<��8?��GtL�ZL�Ѡ���9�<�ɑ�{5���-�qlC�5[/i�/�*4�5�ϒY������;ͳ�eNұǽ��U.��a�v\D�,)����$2�Ei� �9��{��D`}�<*���fG�Z"ߜ-&�E���;>�F���A��2U�Ӓ2���
X�~���k�^ٙ��tz�<t�&Z������u��6����������K�4�w�{��N�0�T�$w&O,��w�bwe-ۦ�K���Ç�IL�}V��k곈���Yf�����f$ ��l��|�����R���kS�3�,7S��g4t�Us^58(�����)�Vޜ߄8��{���wxD����89y��B'��$�!I?|t�=ߜ;*T���շ�=�?�L�O��3�;��+�Z�=M�����ëf�ՠQ2IM 5t�QW7�f��T��~�\5�t4��+�¢�u����gǮV�a9���+���W5R�� $�n&�Ņ�
���@�J��i���J$�I42��^l"lŹfsk���/�P���~_�ǃ�����K?��'���>��`v��=e��D��p���?s�#��1-������Μ=k�ǝve�R[i�MT)��W����Q*�������a�x��R-M�iA��
a?Ii��+a���@˔��熞Wm�z���c�M�n(��_�׽�y�b��'�tO��֖��?���{�;ز��0�����7��zaa��R@�| ~bߛ��}i�Q�t��+�l&篔����r:n���Q�G�ʀ�(9�����l,�sny�/I�@s�z��bf�3�G�F �2@'�Y�����	�֔�̸,s��� ���zq��_(���8�H��q5@���CU��>}�����6��`�"�GK;��b[*�(�h�c��c����H�.:�|�u����\�^�Q��(�HO�3hH�� ���㡔�,�b�f����P�1DW�;G��fΉ�fP��O	�/Զ#e��3��;8,�����3H�^-o�b�쮯�c2�CF&O������1;f͸�~9˞��,��_�Z�W��Y*2(Y2c��4'�gϞ�}�7�ړ�{-~#|dB�o�c˳��'i�F{=<�A`�$Ll�!U�ccYE�
�ǵ�}�ʤ`!-�#Sz�s��g�M�i�Wza9�iAcD`��ZR�V�j7QZI�JERh\�R�k8 �i쌹t�1�x�i�҉8��3�q�c�p'���$�3fe��[���[�2^�9��\�d<��F�j9'8R��K��є��.����s Ɂ�Y'V�lds���˳)t`x3��;2KJa�Y��gkKi'��$R��4�4��o������`�ɹ�ir�i�9�1�s\��h�s/B�����]2C
�\|��ׯ���}����}O^pG(uئ���K����Q}��%bИpY���`Kɏ>��V�������Rׅ��`5(�fdf��J��-����_
�A�:&��;��f:�Ѹ�q�y%S�+�lGLK�:'�4嚤����&|K++�I�rM�C]��L�"nB/KG��Q���3�Zs�I��#MŠq��L(��`����S�0c�pV�e����=�y��nW�]BF��dm^�/`���ZOQ�-���G!'�hN�ʟ�R�M/��Q�&rA�|�\�yQ�I�:RhB� D�I���y|�x����3���_�lm��'?���^���\q�}90��Ƌ߽{��Y�f�up�z����c�� ���{�%0/abI�Ml4MX�uN<g�4Jj�q`����| �_�I֯4���͉�
�������ם#���\��Wvx*,q����ǚQ�ų�(��>���$x*y�S
�����R��q&����gb(�w8l|�OD�O���T�ya�}Z�^��gq��&��JW��`�4�)7j�fZ}olkC=�HG�r�S'��F'�g;v8#>��I�����d����d��D�q��p}^	�)�?k�).H[@��tx|H2*"-w�=n�O8��}-�f�w,�%}i�L��O<�EcN$3�H~�'�Ęj߭K�.��;F�2�]6��p�8��.��壣��D����ڍ��JW��������q�/c���L�����8�j��O�-�i< +%���ҥ+n�H��Grc|�T�$z��a�oĬnLR�O���v&��m	�{��âe��ϒ�U�b{�!D"�_�	v���B򬮮�T�mnK�v���6�t��z��a�|�m[��G� s�A8��LPc��0Ѳ�h��O_/F���������¡��|�6�|G/a*��s�obt�	73)����VN�ٳ@���^@�q=[��[dcM/�����[��w<��eNN�E��r��̳T�<���Kc�V�TЭۣߔ��_�f=X�Ol(��rK~�?����K9��Y�A�+��3j
�g.hԦb��0��`�P�_gY�DJ�Z��X/�9�X��O���D�(��q�7�(��}�?ES4L$�<��p2�ХLd-IKg�`�("|r�%Z����;�(x�t$�}|s����� R�pn�]�'�j2�|q�`�Xf5����:�-�a_J�ܢ��L3
^�S$Hc�+U�<���B��D��d:_�3���DqNJ%S/&���I��4�4�蜌`�ۥ��byc��������Ӈ�	��{��덹Z�wZgV��<|gm��wV�.����8MZ�Zs12�hMR?�{��+L� M��(�B�dT���R�t;����ŋ��ju�V-��� 3��8�ZJ#Q,.��T�r������T�Tsa>0i��pnan~~���#��'1F�M���A�קwr,��xX�W��q)�%�i��)��bX��i��9`��Kj1�xx�I4���.��]��w��_��W�KM�����5ʥj���*s�9�.-/���ZS��՗_N��Ao�;L<���Yb�Oͩ��(�EsGS�Mc����`:��wξ�o_9�R�7*�����fan������e{���n�$)U�Gm�e��uA��K�'�ti}n:�O�/��Q�J�aI���I��h�\�p|Ҭ4��h�Duo�f���ͥE�w6c/��qf����;5�0�D��������o$�ƇC	ܘ�y�?ޯ�4���^�[g�'�;��Ja�D�d�$#����	Zլ@��kJ����5=���,����m��YR�{��Ü��f��O [�_���.��G}��S?�S��_ =O5���'	�}e������y'v�xA���,_��w/_���,��AO?KM��Xþ�"��(�x��Cq��Ot;�ʤ�I{I�O�c:�pk��ʘ���jr	鬝$�+���h��1T��D#����X�*��FCr�Z�C��Ԗ^�z$����%�T�W�dD c�ϝ{A8�|�M	����҂�EW�֕E���᣽�{xp ���%�v����X���tj�z.'
����8�{{���������J���֪T���{�~�,�$ȅ�����n���6�s�+�M��O1EgϮ����+�raI���'Be���mi宺Y�>(��������[!�e@�@���ܹMfS���#���@-�Ls� ���0u�;��h#��ހ��Q&�+�YH7��T۴L�%|��� ]���� A�A:�q=z�l���K\��q8Ox4��*��c�T����XJc�f�Y �"-� ΁4�����8#��X�mZ��lj�u��R%* � ?��r�j�XyU垞��Q�r������f����g�o�\��f.��� ��i�mE ��-�2A(�˚�c5�8
lx�&Ca Q�ߕK�K8��hs�����}���~������w��������
A>�jQ�7���R<�9_k�s�9M��6�b�፫m���d2R8��S�b��Z�<�D�'�D��t���v3����X�x6:W�7���O0�pB�	��_���蕨$`V|�-"�mgn��N���*e��ʆ��J��J�M�xKM�ݻW�^�C�i,Y
c�RA� �QF�Q4ju�?�Z���wr�v;��__Ӊ&�г.b?�6%�CP���<�k;ׯ_ǥp��2��}_�zq��O��-�t�'O���/ �9��K/�,\_�S,�;���qq�|���=z���2V$�iG�p���x������5�VP�׮]{��׫U�dP�8��;������U������e\(�~�=:�%��#?|ޅ��d����<3Z�̉����h"���!�����ئ#�fS�g��d)o��6 ����=�>�e�&Zq���3�jIN��ؒ��`,�4�f$���kX��+sUp���@�����>�bF"DL�絢��@��K��ӧ�^�k�&
�qb��stҐ^�^�d2�I"V&9���� ⯼��Ml����t�{�1����k�?w��9�|d*��c���#'}E���l*��LGX��Ͱc��lt�@A�u���Dt\������è��K����늌��h��2#-P.,
@�Y}GGҺwqq���o�l�d'�-�lڢ2�紉���P-EF4�B(�}M`r&+!#U ɫأ�z)(�R�"j/�E�ޘ�D'�x�vw	�b��4|G	��$tÂbZ�j/*`z��5'��ɣ��@��;�@gdA�.gϮ����|��]��&@s���g����^,��Gn����..9L��6�,�H[^�^�S�lf�s麀��0W�B�st"�V��D�˖:+̚O��$���7�� �OJ�Y�Fϱ4,�V�$f9��hו6�2tsˏO�!���ͦ?R�A���- 4pXX��2����&�	��9����sD�ev)��b�	�<�Li�搨����Lէ�F�y:�"�je�l��˓ǟQlV��^�L�P������f&"�N��j��,���W3���>�f¦�*ƽ��Mt�ht)�P>��n1��G�(�`r�'��ț�`�"��������aJ�V�	�i��JX����u�[�hv��)3O��T:�ah�T��fZ�8,<QJ3��c
W�*�3�8�8�,�����).�J��Q�4'a�X"�R#�J�fd+�0跥� 
���Wqk�Ϸ�ʞd�'╲~�rY��dWI��PT��G�T�9{}������4���T��ymɕg˗Dʪ�[ɬ2"�qV��u[��s%q�q�DY�2?I#ml�6�	��FIͷ���(�b̅?�7�4�|��A�l���������z��9;1�V��&Z���څ
�+W�/�������盕ڍ���uj���I7z�����	�`K��+��~l����;*U�%�nݒ%�]���|^�Ibˎ(�D�D^�ZY[]1�t�Kw�$�Hb���,)Po6s�`ymu:���^i\B����K&��M� zn�}����N8�p�|U`c9�؇�n+� ?�g��^����f�������Oz}�(Dd��J�}���L�HQ!�٤�1N{X2�t�q�^RUС�U�a�RN0�d�U�L�8��I��QbR�����f�%	/�5ҊNm�c���\�)�H��vIw�ޥ���d^���F�s
Yf�R�s�I1 ���&��#���!&���A����������tRpEu�}qV�Ή����ц$8v��No�6���2���B�.��a8�%�ݦC�Id�� C�Qk��3|@�W�\2fOG$������W�SaV��@�*��L������Xq^F��(�R�Dͩ,^�:uà!�����2��Q�%��h�����aK����C���;d��+�C23������H�/d�3/��xt\9�C@�Xb��v@*0C� 7��2oس������O��h00�*�}��?�t�RPq`<���r�p9��v�&>�	��x�<�p�$=ļ��Z�F~ǽ���y��X�わ���W�6n?M���G3z[���	A�Y�_bYg��ig�9ܴ�Q�b��<�T8K�A(���т�=`�i�M3��{��A�ٛ�i�aM�M�V����"�р薧@,�x�/���Q�^ �М��=_g���|���I�=W�9K?;0&!Ӿ{l�J��ln���W�����]M��i\��D���9M�}�X��QRK��t�ܺu��9'5eQ_x4����.�<,�^�Ô��l�UR�?�����csT�� �<�)3�K�T�i4��:گ����\+K��h*��r�1��
��M����S�x_�S����v��%��$c��[j�d�Jt�J�}�V�[ַ)2:K��f��s��iR���l����9�w���x\�i��L���ˑ���E��^vbu���Ű�f�g�o�a���P"J����X,���	f����z �I�f���6��N��������"hb��W� �N0 �>Zn!6Ҿj��ի9? ־�D�RL�u��V�~�:�Y}Cx��DLv��j��\c.Tꋓ�^C�����&7���zG6ݐC+�	�666��s�n�_z	0�*�����!	)B?�UP]Zz��'��"�㱪I��M���`/�i'�/f��}��ו���)��'��<���9eKr�N1�=�"��+@����
5�um���E�8�90>!@�(�,��o�䮞�� 8=�����kf.ӟ�e��r���C�x����4Xbr㱽Rb�hG���S!�#�{0���6����QV�OIL�!K�8|��a	RK�E�.~΅ @����*�Y�nV�`�aS��D�����׈�>$�$�|�O̲"w.�"���H$� ��gsɉ�Ԍ$r�#M[�8����j�d�v��C�4��)�rN�)���v��f���Ą1��H�MK��,uQ������uf��L]���}	�m����G��uj�X'+1}�j��9rP<�: [`���ݣ7�e⧶��z?��}KK�����)_4���֋$\��c�ꫯR
q�����S ���`�㬣F�^.�ƍ�5�T5z6���7��^F	iyv��0c]�,� ����N�r��&fŵ��7�|+�e�K-W�C-�d2r�?����Z���ճ�Ӊ�0����b����=�ڞ}?qCB[,��2�ǣP�3�񒭟��b?w��^�(-}����6��R�a'-�M��RJ%u�_��lkk���K*��&����"40e1���\���mn~��e4�D���i:*f�B��?�_i%Hr�T��%\�P{�?�V�ז�|����>�f �z�?����"��__��9nV���t��I.IǩH��틯������[���_�Tnݓ�|��&��bS��O�������jT�����jnA*�B9O�^��<L�ss���U�n���R�Q(��ڑ_��e���pY��)�l�v��z����wީ��E�:�A�מ�XJ�:/$%�:��b��@�|�PO�Q|ZQ��l� ����؛�X�^Ղg���Cč!#r��++��.C��v�Z�� !@�Z����^#�?n�e��F~��r[23��.�\eWee�rb��Ɲ�z����ɬr�å���s�iﵧ��8.JR�F_0J8�8I�ފ�U�Rf���n\bMz���,/��z��m�f��G��c��Ѭ_��5CKX�����~��W��J��:� Rw(�q�ln�6v70�Ņ�R['���T �^yccs�]�t��}�p��	d"��+HW_GMd�E�]���g� $��l���+��6�R��H��a������33���O��_~!J�	�Z�3�'I�%������.�ދ��I�O�a�
�ܔ��n=��$��6Ww	��kC�u��k�5r�*^p��i�j��o:�R���决L�]P�6����äx��X��T�u�U��QD��aZ4愱 ���f�E�gr�z�@��#�(��ek-����s���S���]zD8@�O��p��aL'�ޅ�"	�9��$Wc�t��M�:F�)�h�SM:��*/pW��/��'���ⓜ���ۣ��"�1#킊OJG?5�c��T��>Q��Vk�-_��3n�_�4�h'eB�̬,�F'Զ������ʂ[�ĞQ��'�ye���y!TF�Ϡ�������	I��{6��M�����ŅX;�j�{L�g�F���e��CCQd�J��b�-����~pR.'"gXPC@5z߈���i�;r�pc��>c>�EB��(����7%ɉI�b>���J"��;C�;3�ȣ�C�H:Ñ�*[fe���6���/|�����y�u+����he�EZΣ�º)��>�t�@G�Đ�p]�,�Ͳ����x��1WK�ϖ��8~1?"s��z��䚊QN]��l��ب ���o��{ug'�'ƝdD��U�w�҆�2D��^��~���?�������oJ<"�D!��+L������2�$as�}z��D�H����6%&ߝ��� ��$}`�1� �5�� �H��o|�$�Sڌ2U. )�쌸���,m�=��o(��#.��l��s�I�O������?V& iuum�Mc�
2�&6�ÏE?X~ ���,�+���j3e��ɓ{�w0�3SӢHT�8E�
���C{��ٙK�66�@-/��~|���O�HkK�k�y�����cǏjm޹�yLćo޺E��1ĉw�I�#�/87)޽'���a�?���\f���`����})V-	mK�HKz��ؚY�Gм��ýV�0��Jf�)���޵�)cN3/zf�n~\!�cI��l�%7:<�A���2y>1���X�S�1��Dh�wDg�������d(P#J��7��G!�b��#�b�Sj;8Aa�l}��֦����U,��'�IY��=��<��=�(�OI�e:w�/��>�vНP:���y��=��.���p�ڒ(`�D�)��03L e��X�}u�1��!3�0�G�#�1������0����51���̰�ޑi=B��M33�nw�ysMK���H�v�kv5pL��ȴ��*S 3x���i�g�a����_����P�3x�8,�@�b���P�ʒ�j
}'�J��IK�Oh��R���=g�i`��O����C����@6x遡�e�.�ϸ��DH�LF���g%/��p�#fXK���R<��_������+#P,ҧg���8���.���$R�P���uߨ�����yS#���Rsr2�d'�zY�/_�(3��D�]Ì�h�uUb�OG�A�Z��}�T�(&���'��
��W�\���g�]�������g2s˦�'��g��(�YI5����<b�5[����ˮ�h�*Wx�������Lb���.F�Ϛ��I�y���{�{25���o7'��u�S���Iu��p��,������g]����O���l��E<�!����G.'���\Dت{���𢾙r��(�:G�7���H�S&&�����lty-fu?��v��*7�B�Kl��`F�g�J˚k�ba����iHY�JC�'$�����ܹ,I�^�{8Q@�h����3x���S��@�'��Z��0cw���x��O>�j�@�|�Ǯ�N�u�	�u��-%��xY�A�S'Vq\����5<�8��.�y��J�<����(��^8���0�����D N旖mG���á�@�5�I�1���in�B�x1��"��
�{��N_�Z� ��:��H�T�ó��M��R������8�Õ����)��l�mn�kD�'K0^�O���M�����7o����Dޑ��GI z[/���7�"q&I���& �x ^�zU8A<-� aR���A�R��H�ƅ�1c�`R��_��ǰ[X����`Wٝ�(��x��r7�2M�f�"�����\�V�I�@�vk����ʉ���U�;����`��Jc��s�ƻ�{RT�#�P�FG�Ƣ���D�7EO5hRvC��Ix =Zjδ���ޛo��s�)�+�Z�#=�t��V�y��!g
�0$gYw�8��y0�k�dm�� Z�f��3gX��h�3Î ��g3�
Y"6*	��X�s�(s!t��H��X�ŉ�$L��(����*G���f����Z�Aj n�E��A��� PV���
��	5l�:n����2O��a�Kp&�1�"�D�?��fh�L��P[���y�0���h<�2fc'�����*�t�yƵ�EPf�|
�AE�(\`'z 0�v��N�1��0;;O J`QV�z,z�p�z��?ⱱ=�9
X��R�I���ĩ����[�n�3����,����ȮtNp�7��%IX�a#�b^_\z3��m����Je6
3��7���J�BY��v�	�\qk�Vke�$D� m���nr�V��Z��3�w�:ضOK-�X�|S�Q�7�7���eU,�l|o^3߆.��v�#F���-�$�h���u<�]Ql�y�#B�3!�L���t�$I�t�����)�e�N;��m�C�t�L�l?���
�<$z���5�}6��~82m=m�61�s�EӴäT�X���g汚�]�H�gN���/���Am��pa�eGq�N�:�D��<걳3i�w���m�X}��g���q�H�9)���G{�~/��H݄��Ի���)g�����C��DJ,Q��Y�,&��V�P^_>I(�D(θA%��Hv���<��%�T��q�'����/BpO�RnA��TU�w�u�oj;`J��ͻ���q)��*�v`��c9H%���E��]�p�I.H��:uj8b朘�.]�F�%ǂ�J��Nw���˷� rs��ov�U���D5�J�ĥ7����� �3��ݾ}[�]{���U�j�[�������5�M)M�*Pw�����ƴ�ŝ�S]WyF<����}o��E�,�P��������[�w�y�M�w�����f���3e_ ��n_�׋��W��޺u�/j6�ʂ(M�����V�$��zKo�ׯc+�+���$lM&�����)�%b��"b����y��[��{�1��<y�8tm�l��,��ɠa�1�T�U9��!j�����)Ƣ '��*�1(l��f��ݻ�J��NM#j�(
~`�9|�q�R[$803^���J�ɶ�:~p�c��g/�^��˄G"�J5B���{�E���v�o������&�f��IY�h�7�>e��_H3����c8)��_�X=�����(�`�^4,>�׸��l��!��&յ�&�::��� I�F��С�r����q;�E�	�Q��]R�$X,�'H��4�\�٦��hګ3��aw���{��볳S��R����{��i,"���ʰrl( 0��"�E�K�7F0O�\�����9��t��x�Qo]h�h�2W8�Q�SgSq�?�
d55+���5�u��]0"���O<�M$7�c̄�-�4���>�O\���^v�b@��j�rEj�+t0��xgB��[4���= xx�%؊���c��=M���i�U��C���������4�s�dFQ�W����-�bCo��U�;��^�v&�Z�,���סyS�+�4�
�~�gM�������S��_��{Ҫ�5mà�l�f�f�e�'W��n�X+�%,��[Թ��;6�G��g�+MZ]�wMmfj׌�=r��؋X�n@[�ǋi��ƪ?��R,��g��q3>�L�Y�G�
�,�x��a**>�49��-�%�sg7�)���j����,��f��S7$u��Ts0�I��4�6�%���L! �Jy��ՠ(k���m�@�\�y�a��++(Iwo0���A�	�@Z��M* aT�W�~4��/|L}�uZ��Tu�����F���|�#��J�^K7�f�R���-�[��9&��e�BYU��g���ʱ�u��z�%^Ù�E�wc{{ii���w$]����w��.��?yl~go7R���R��s�$�.�Y�����-�;.T�!ƣ��R*��\�s2�'	΃X2��|��$
{#�2�m��^q��z���8�3�u����+��Z��4�>G�|F�)�����B�;���FT��[�޻0�0��M��x��*����͇���1I4aD�0��!q���Õ��Nci���+�#-�L\�;�7ɓ%��DÊ�t�j�.&o$F�h(^+�K/���_�������L��rI{�6*��W���{�]�*4ͰP:_�xa�]���n����XL��Ǩ<pq'i2�A,�oѾQ*��ĕ��Dyt`k/_�>������
5�Z������W��~�=7���R�i��d"jc�,w{�H5�A��;���[ĺ,j��0���0K[[{t�0�h�Q
>�.�N��H饞WAL.�z~|��͛8��=09xf`)Ғ� �X���06h�ǆ̂J�>��q\ӟ��O�(*�h:c�&#A^�O؇x_���N�r�@��Q	aɘ�E~��T�Mq�5d�P��dd'�ӋQW�����~&�a�_x�;w��2��yM�r��5b1���	�gH�������w�+T|-b`N:C��k��鿤J����*8|<�ٳg K��u��&��Q2߷á2c�M�L�}8:������N���z[S���`?Z`E�f�9��-��O�����#���$U�ؖ��FS_J���?��W^y�������T��2_�{x��%R�k�xx���O���J�iH���m�%�bO���fE3�@7n�����d������H��)-g��1�ؤ�L'�(κ¯��`h����ŋ��.�Q�b+w���4P��0R�cOi�9�6O�u�$m�)`5I���e�J�Oє�305R�Rt.��A҂i�E'��%M�GgsטS��0���Xj֍ժ�}l�A$���ڬ�S�QSM�$)�X����LM�ɼˍ�ɂ`9ߛ΀�5�w͇��*�Qlz�ۛ���GF���"���=_�j{o���z��֓Jk�(%�O��μ�~`��H�(��G��
�oj:Q�� {���[]���g<g��"����+8H⁋�)V����� �#��|��<wO3�]��J2
��\�N�%���z���LJL�.Q��{+���-q�ܼ�Gm��*��y������ٕ�!%I`/�x������2�4]��C�S
J�7<�LC� ���K:�����~l�c��$�}�}P�$����B��^b>GCuH�{�J1E�+�����?�M�P��aJ��b�����w9��|_z�:-I��<J�D�߃��[�ǘ?�D"�\��!�$«�?v�#���PD�N�@��=�*��|�}��Z��?u<r���]J����F��,\��X,H޽�-w�"���N��Q��e�=Y\/�S�*|������gf��d�jU�Xs]�ǽA`��9G)��J~���<6�W�jSH���_������5�z�dFF����+����'d��u�b�L��J�w��.�%���%�y�VVWX�&��66���D�w�kT7*�8��e���p�xt~SC3}�)M,��2��u�ۭ8>C��$�
L�'[����̌y�I33�f���	����8���]�� �`�=��4#t��qq� ���$1���?c�Q���Ŝ8��.��S��Pa�[w�xLO�d�"0&c z�ڃ����D1�!�U�j�a�}���+F�S�Zˢ�!+���D�x�ٶ�6RrA��R������$"&Z
Խ�l?ܔ�����&�{��J��kt��:L��2�fJY������16$��� ���0��d��H�Ī�!d �UPˁ%��s�Kb�Rm�}2d�٬�+����_/\80!Nk��!���P1UjqeWl�u	tilo�-���c�>ܴ�r��֝��05����+〚ϳ��'�����|�S�����{<9]��a."�6��ܹs�>��6�Ёż��b�A[`��(�ϒ[K~��(1�>	(���U�g��YM0��
���-%9b3���/^G��G!?1����u��-HM�ވ[[��D�M| 1��|�"�㭵���Й��^�5!N̊���؅&��|I�6���jac��}u-��z� �s�_�Ȓl�(%����.��wq�����29xB�;����Q��&�u�k1�Ƃ
�x6W���	���8��V��eޜc�/1j�ޠ�"�͠���ސ�&v��VG�PG��$u�I�F��@7,��.~s����Ea���>��+x]�\�����V��Q1�#�m�2�*��4�}�$�����x~~~����;�S��/_JbAz~����͛�����a8H�EI��i���NB�M���!Q�Hf)�4g�u�&l�^a���5#�슧&E���i���ad�r����*�N=���;oloo�ꕝ��]8q�`_��jպZ8�Ѥ'���2%��+�Y��V�$@�m�R9�t��j-a{��l���k(�����v�{�;iӇd/�����Jn�_x���?����j�A$�%(+#vzt���uY)�y�Qu� �8u���t����{�������L�T�`��k�{��2?{'�V;�%\��tD���LU�q�F��o�8Q������2�Ʉ�@P�x<�A�y��w�қ�oa,'�ڤ���Љ�����N���BQ~��a\��ʲ�����I�9�Lʮd�'��p��[�K��P��z�0����VWW)��ED7���(�)�Iv#�m��Ư �l�(�7���G�4�'� \ӈ�����v�a䥔��K�/NK��Y&);��ͼ�6�["��;��E���!�b�'1tP�:�����R��g�$��Ǧ�b�r����U �W�XvI�����4��b^���`��l��<���&P�3r��Soa�4��E1�Ȣ]�ɚ>Y��A�X���|R5Zn�l�N��'�>~*i.����R�d�x�
s8������:�]���M�։�`�3`����d����WI�TX�3��{�z��!>�aSKWݷ�ጵ ̰�2�L�Mq���v��"9�k�hd�!��>`�Q0�|�t�bat׮]��?�����ߟ�jb�|����vvv��2�T�"m|�>�'���̈�a���4��ȼHs�$ ���[aq]�p$�l��G#q6�:90�:v	�H��s�6�������}a��f^Z�]lz�����y�
�L:������ʗ���mC�E�f�qfd���i���r�qD�w�h]yD���~ 9�QX(e�xrq��N!.%�b��1���X��}��"Ԋ<��ixHHzI)6+mY`�E�:5��')v*��Zt��J��-p.h��Z �к���绬��X,љ>�J�L�C+��v�޹#{A������4U��h�V�3�%]���	���(����R���ō}�瞹�x�����Wԗ&Bv{W��fU�(ÞU�ca��!H�d;��yqy����;W��nm�=|��BӣD�Zx)�7��T	ZU��_e�l���AU.����ܮn
�Qz�
�A�L����"��h�^�8q>�'1�~��6��Q�N�N�/0"M�\y
k=-��g���$�"�����nH�	��դz �\�Q�f;���CNM�e�gj#��^% �� -@@�W6���1��tS
��^�=H���6�e#�2Ej;��3d�_��#.�^�вn���`	bWvo����^>wN�K߽)�J�_T��D�'��)
v=�pf�<x�pW8�g�����=��p�����"cp��h���sH�02-k��I�r�����T�0/^�z����bou�
�)˻a=�T�|ײ!zJUEA�/�~�A������gp�NO(�!��tfx����4�Tᦐ-L{���/)�5N�!��W��B��Ͳ�)8�|��a��
�)bl��&FBSmK51|�t��I,2��B���c/���Ʌ���jU
=G�*����ų�G��ù��ҔP���P�;�`]�D� �q�nܸ���C�VPB/�����p�TK���^kb��w���le�Q,V����#	;N��.'��v:s�'�,���
���e�Z�{����pL&�6!��q��Fj4�P�
�~d\�~_|�sx@�K���K���p3k#t����m� 6R�1��X�����Uf>':�i$��+�Gg \V��-}���/|���˿[��]�W�rc�^��a�ؓ,�H��5��J��%�E��k�'���:,��po[��Hz��(�bCE/W�ie�ƋX$D�a�5�,@�@�;���+�T	z��ʺ��7˴��=K^�S��.�@�8{a��r���G�a�91�����dZ�M|����5X����$����+�L�A��r���R���A��Ŋz�A�f�$&��W�w��]E;�S"�t�\A6ɳj$((���,H�w���IfkX��ѿ�/�UN�8I��}��.�`0�mJL�𔇫;� 'g�O?�\a8p��T*����遜h�q���N<g��S�L�Y�p��69y�8���on�@���I�fg{��;��RY4}urx�������o0!�\f�#�$�y�t������$����������@��)5��S�s�� ���Y�GO��с⡝�2��S0�:�C��NW�XcGbS�m���6U.�B"�$"��O����e��E���Q9K`S�(PRd55b�non]�?���?�|�]�ΪU�̢���Y�_y�ד@���ܺ������o�i�!�G���<f�bA%�Оa7�%� ������`(��q8�j�Z�v# ���JE���D0X�fU�������e�eq
��5����ɈpV�W�<�m�T����x�%šY�)��������4,�R}��9�_QF��~w8,���$�W��N\����d4�YG �j�}0�f��aPd��]Z:yguwv�%���1@-̳&�>�k$Se;#i's�]M���d�({S�H��5�dU��8Ѫ46D�k0i����Yb���aAh��8JOlD�Q�QY[��'����4Ԉ%c�'�ط�Mfy�RM�4y��������t�|����E��/��@J|�ZNX +��1�3�
�l�; � ;>�2����ҥK�����@��ӧyw�#�T�ׇN�l0@Fc�Z�:ۚ��&�x��O�:�pM|c�ד���� �|ͣ%) m!v���k�Q:NE��1������ �)h �#	���G�a�5��ad���LA���͖y�'|4��׾���|�������F�P�5��s��n�	c�������j;��d��N��QW6Ⱥ�:t4�"�&���aϴ�$R�r֛���D+6�	q#a,�&��Y�K����`�$�V:��<�4/��O����Y�So81=9�GC�f�zz��\�O�o,>��vr�M��"ãk�I^F$[��7˵wmP5ɵ���z&�� �cZ�9W��h� �6��%��>�K[�t����4M���	�~�i,؆����YՊx�������˽V��+�A�Bk�fi�@31l ��Tx�(S�N� �d-G�c�KHJ�p�e"BE�lr�� ���3lJ 	3�Yyz׃�����O�}�^�NUxj��(Lia��P�cZjD�i�&�xN�G��;x:i;�N�g�[^�wI�5uUf� ���/�m�q8�j_}S���A�VBF��H�Pϕ5�&z�����Yi��àV�v�;�³Ϯ�o�߇���5��^Ip_wu�|���W�q�B��Rb�^x�x����j5����u��Yv�e���.'����:�ʭ[�0�O=��<y��d	
j�]�xQ�W���8���|�0H?�~���U/10���$���+W�� �n�Z�z��͛�@l��\M���P���ʅW^y�kS�����-tzD]�I>c��ٱ�J���u�^ jr�I]��k׮5g�c�V֤%�V�?��ڔ��P a�4�#Z,��m��m�t�2z�_w�ȞH7���*t��Z�^~"#�{���ݻ�pً�N�?��߂��P)3~$j)�s&U�P���	���x�愝�p�<ݸqk�-u^�gbe�g�3���Ќ�a}S��+��^���M�D1Llf�|SGѳ�>�d�H)I�bO��:��Y�4H2^��.K-:�"�Q�^󭭌t�J��!%l�!�e����to`~4o�I��1EU����r�bgI�Z����pJ+(�i�����f��ۘ�I}ϩ�bfP��)jr�A>LO7���L�f�?ƺQ��ذ���?1%�E�xH�k���L����~#�+4fŉs�AR�
B'�ړ{:�ҵ/�+v�¯&�D���[�|�ĉE~2Q�W���l��nO}����G?���㎡i��m����ܾu���~��pqn-z[;��R�B�`ُ]�Ҙ@�F�t������ѭ55�<<��s~�߿�I������Z]]Wr�J>�g�*����Ω�x�ܹ��~���^�Ї>D��R-ZN�/~�?��?�٦���Z&_�Q�C�0v8b:�����z��Q�T��ݢ.2�/��]Q�oZ<��ӬEE�#�x�\��fR�3gR>J�������mn%�*�7Ǆ�mUo`���|8���*mE�̎�%��48����o�!��\�-b&~%}��Bo�ZT�sw9��V��ד�{;��NV!�2��(���q�Xֲ��Г�q�	
�/��Y_����h"�@7-~f�)l�6�g4��' "�۷ok��ta�6Jc�z��M��R�m�o��:yh���I'��EúS	��L��$Z���M���p�7���s����hyy�����JS���}2WV�Q�5��yE	~������'���`���Txm}�)2b�6kt��������?��˷o�q�����#C�Ud��	F�Dz���Dvs{I2Wu��\ 9�I�ZB�k��H�V�V�/C���9<~���ӳ��,��v ��Ik�G4GQ�̫Z��k<�;	S&�˺��v��uy��	��j|ӝ�c��r�� �L�U�)L�7Xg"Mggf�f�+�k���Æ�ãT���R�9��� *�X��Xk}��'/]�N���4�J|�_��:]��� �S���S�Xӛ7d��./,?��Α��nE�6^�7�(�#�+^%�gkX��l^��u����I7���ߓ�@�5 �������x�"U�[�T,ת��9���$�F"����H���:㩧�F����WH�E�B�ŕe �f��ǈ���������������S�&|�$��/2˄�}��-"��j��D��)@(��+;�c�)L��"��a��nd\/2\kĔ�"X�;w��C�0���A@"<z�%�w�(��U�,���&��� leox��i����aT�T�\#i���ҥd�k��Z0Dq��SX�U*U��+���[Д�Ç��zP�"�U�֠���1��U �ؙ�G
<$�u��$��R�6A_�O]81=BmoZ0�-����l9E�J&�nw���O}ꭷ�rc��F�Ɇv$�U.���W����� w� �x��W)O8�,aQ��(��xet6��kNM#�#H�HuN�M~Ҿ�U:V7�c!glcKlft6��s�=�ꫯ~���ƛlhk�-t6;�9����旾��_��_�N��d����b&�I�v�n�z��l�Y(fqC.4�n*G��8��fF��z!�u��KL�����)��mJ�c�$6G��ђoj'�G�p�q[�����Â������LɔMwK�k|���G���M-�̿�r���H�r5�A#�8�	��[�Y��pе��n?�H~�����h����qsQ$Ѡ��U����t�P+��q6�)�X�����g~؃e2μq9O��gM��2ֶ�o�K{��1x��g�Ҝ��kmM۳Y�<��rlaw���'��o)2�@{�wa��j7�����d�MSS��'��:�
@@�w��mu'�O��R� ��/\�p��igM�0�H5��2ڝ��q�~������ZZ�uH���=X~��%Ry���լ�;�k��z"�qkєZ@G1��o
��D��Fʳ��S!��_|~K*_��w��v={����Irٔ<�$��5�b~��ᡪ="��JS��z�b�t�*���-���뛞'�gS��
��m�j�V�"�	�(E�z��=q�lo_�~��
x��l�œKɓV�ް'���1�,�ƃԥ��ϟ?�}�S����MOE�Xa(m,3V��؊e_-iA��xX�7��+c��wmm/H�Wt�)�v�6{!Pa���A/2��1�9�iI^j]�p���h���Mgv4bbM���d����H��5cbfo
S�ޞ�J&	����?�h��k�e�;>C�7���\%������R2O^�������%MŮ�up�p��@ZK�DS,b��u�������2��"���{ril+��qV���r3�ɖ��
��ɓ;;e� c�toа��ǎ��d����XO�H%����aef�{���wl��z
�:�ŋ��ݻw�Q�8ZHX�!��l���@��("���� Z�g�D��iÅ-,�tYB��h�!SJ�i�כ��t�2�[c�D*/����8�FtDq��#��\�����>c���9Kt>��c��XᲫ�K����r�U<;��CRӁ��F"�U8R�٠ø��Z�c
=�"0�Y;
�u���V�\b��t`n޼I7*�3c+�%��}����?��/��/�ZMlr���oipS��h$H�oJC�ϖ�C�qM9��h�4���ٳ@��&�H�@�a��`��W��Qь�v�gr�NL���.5��EC��va N����"��\
WѴ��|����0y��B�tG�ۄ��Ȝ5��h�4�z�������X�cM�j�{�M Ż�N�r�͕��G9'�����7��BP�bM�	�R��TƣI+M�Ż[ۇ�&��6(�"LO�ƣu��ZL� �<��>D�P�|\
JԸB\��+
`��9�עˤwx��^����0���F����,�R"�����s���鞄o�c�ƅc�w*~��>��Ng�܉�V9p�i�P�x�8'�P{n����sr�n�x[*t�*�M�pn~~�<XVZ�������h85�J�ɍ�����W�Oow:gNKk�	R��x��S�{��ҠRk�^�s����+~��3xR���K���8���:�ͩ�'���ߺ���%�:L&�j�8��V�)*|7(t{�ɲ[F�0�z���h͊�(�^�`���i,k�Ҹq�F� ��{ې&�����v�^n��{�d2??+�ѩ@\���$�.z<?��D���\��i�g(����AF���w��js�O�n����P��ݕ�\k�=si�$,���{�O��Օ-ܨ8�j�����[��O�E�5�F��q���XDjc��+0�[��3��Z'������^�ONJ�Y��}���#�*
��x	��:���U'���a�}�}��:�U�]�y��jՆ��uؐ��֨�:�E^xI	�:b{��P(�b�����w;O����d�_��o.�<)-,k^�S��̔�������8�'�S�rb����S��&����B	�=:{�|q�;��svv�Z):�������s�$�y��aB��o}K+"ݙ���1�`���� >C?�s�B\bE����0"*���h��G�.꼼�����I�0�Ř�@�)��fhx0�W�T�?���_e��'\@�5k#�{ｇ?�+��5xځ���E=#��&���!�M���JZfi���2�fN5M�#@�5��d��ў,���t�(eLM-�-�Gg=����_�T%ŗ�^�ZI;��� �Yf�������F����D���6�W�FXb�1F�𕃃,����;u�D�^��چ�J%�:6N�:�9���mnnI�Rig�1��4~���E��I:��±��G_��_��_��^�*!�jY$ �%T��/��@����}�>�������$�<���5-���*�ȍ=�o5���#I���!��h�D�0��(�0���%h�~��T`1�v�>�z=+jn)57�I=�����w;��%<����o�����"�c� 3��g�~�K_����O��O��4)���Y������yl]-I呛B������˓=6xHq�l
���8������g]�	I9.�2"�(=A.��ӌ����i�*�r���2��n�lJ=�
� �Ǝ��g��R��-^爎Y�je���i����#6״�
L�4�H)��<EK.[L�W�����o��iE���'N`w�J�	��&O�:[��8�Q��K\�M5�el�+c6����Jz&�g��9�f��rY�tl�ki��#��H��cM&�Ȍ��,;m��U�Ü�TRn��H���
�	�c��5�񉶉t�uF�w�f43�W �8ЖM����)�*i"������A9b�*���W���Ƀe�d��MO�K�Gj̉:�9�� w����:w��p"l�Pr� V%����Gr���]�d��Z����,�^K}��ǜ^oIТf��V�mMK9Ť��P{�8���g���ĝ���~���=�j?w�#��V/�3�Р��hL5Éb@��'N !�k�G�����Q�%����ţ���;��U<unQ
�jeh�Ɏl�^؃�<]/�4�슡(D$\�Ԕm��|/�&-���_�����W�)���-,.��t
w���6;�u�w�{�L8I[�F���� ��hJ�%��M]����&D6����DL�F��dg'?3�����J��Ngo�%�����}���>-��V��R�.�aF�~I��n�'�l$,2T�X&�n��o3��=���
�ݞawK�<^M3c�o	hS�-&�
D:�l`����I��m�\7�Q*�5�Bو��&іJ���0��%��m�p���=�=��I�Ű���|+����8>��&Ļ>���`67���|��פt���Xn2��-.��`��������������o �&xt;�=F嘆�\b����#�T�<�ML{�t%��π�$�#�0���Ң��D�9��+�;/�������luz��L�
9�j�;�����(�A����}/	e�آ�-L��'}mx�%�}q�?��O�;�a.������-AY��776>�����O�85}NRR��:^��n�_��sO��8��A����3F<���s��2Q���L��!r<Ij�Z�k�	��KQ�r�u:��O��O���k��%�n*�(=S���گ�������~o/��`���xXz��H�rW��|q"aMd�����T��	=��D_=d�iE���j��{��z	ײ�v.�ətr��l]DD��o�ʂKb�9��G'ﳺ�w�Lk)�|f�O��n.Njø�p���ej�X6��~���$����0K�2����}όQ���C����4�����R��b��D���XY�/
LK�(pI~Ȩ"�"E(ZY-p'������h�dՌ�$���������X��&03��1�'|�%r�]�gܪ�F�ؓ�T/�� dU�����(�
��W
�v�Tݘ�Q'�l%���0�z�|j�l�o�T�tP�D١y<7�Z�?IͪOz���ݰ��NMO/Vf��ڛ��{���7�Ʋ�'��
�6f�N��x��7�ܺW���X
^<1ی�)�`�s����T��J��`{I:�+-u���H�@{�bټ���O�<^��77�^oss��~��f}E�hmc�,�`4����'��+9�3N��S���;��rrڱtS�k�[-RX� ��a�ٞ��w*��ݼ{�~Uu&S0�?��v�/��{�ĭ�cO<�D�Vu�$��dN5[�xĢ�d�{�;];}]�!�2��ZT��a)8�ֶ��bz��?���0.L�K�sN_f�Е���H\A�����ޞ4�k��;�޹=���l�m��6�R�3�B��,���x��L(I��o�rh�b��x<q�B"��j���z��;����P�=��'~���g�&_����ܢ(�F����K�HUj0v���0,b�
��S��u���\��U){�kH��xH�s�DT��stސF�Jy��JX��ާ1�c[1$��(�фJ�+�81.��Y�ᙢN)��!�/�R��ϊ9׸,^3/c0�vj��a.����!��������7�r�)��ܯP?xN��e#Y���2Ӌ"{h�o���x��!g���>L  f���X��+0�ld��2�����k,D����7�MV��b}��&]�%�CE'N���%��\1= ���r=�v�1�Oj4*�Q� nǮYxI?�P2C��v��JKv&�B��r��++s�2L����I:J���cz����'��v8u��f�:|��϶���իW������W_uMs<0��1L�aX��[�i�����kb��Z$G�A��45"!k��E���-����6�Q�H�MZ�����g?�S
q�Y���gH��:8M���+��51�|f���F��<ņ��Z�I���,1�L"93�YR�3�~�F�<�q��@7�C/l� C(����GK<��ٲ֚g�ɷ��5g/���di��D�}χyԄ�s�7r��ِ�]�<Z�c���cа�5,�[����@͢:��4�N�O���.���!'���3Z���<����aPO�e�D����tM~�M3�*&�Ϙ�KFY��Сh#'��%k+���w=�亚.JG�w��t��U�X3�0��!+��I��<��fv�4�HRK�Z7����J^�wK2\������]-�.�"�����4��r��X��7�����%!��H�,�9���?��%<��)�w�G���NVo��Z�.��͝P���Pp0�������=�b��h7�x�b�1���F�!�^�!���&�N��賊�ls�T؅�(���i��U�D�p��%�ם�6�>�۳��ο���m��խ-<���Y�����H����T�hJ2���.S�1�E��	Z�#�+uΟ?�O<x �u��� �pZ�!R�������B����;4��+Wbm.��K��Ht1���}]�<D��םCm!+�et�5[МZ:�4����9��ʋ(�F+��> ��u���5A}�-֜�t�aO��A,�ۢR��A
�G������2��S�'����Ьi��tr�>r^зMS�n�K�t
������ԚL��Uf�PfaA�5�	��C�D�>���<X���Aq��)E�0��v��m��۸@I{�F����Y@2<����3f�`h45q_�p�á�}Y�K)GWr����_O�:��3�H'�؜&��Jf�_$m�h|rS�f�ϒߩiȃO���cc�c��� �8��ʊ��-�1�/#wtovTL�HN5�U�DXS�`��֭[O?�$���&�"�:�Co7�$��G`Z=���K��Ӭ��թp��Ie8j�ά��%�LDƳR�x����:.,~�ԢF�~�Lx̾b��c|���@�F�`��H�y�#�E�[�s�_D匍�@��Q��o�*!�$����jV.\�^����O���'>�/|��YPT��s�[�?��o���|�?���c���X��b���!c �ʞ�L�#�-r�s=�-� .b�A�z��)gz7�
�d麣Q��o�1Fi�8�X�\H��	��܏e��O��h[��]��$G���1���$&�p�[���k�i ���c2��o2	lT�D���?��Q�;
[��k���H�h�� ���nzTfdŻ�+�{T�>��������Y�\��j�$��4A ���ING�4yAc"����@�!9K�b�|��e*e�á��'�D���HWLC�m����Q����3F=(|�$h��/(�(t�I؞�@�p�sriɻp�P�v:U�"��(����w,zl��w�:�A�)v��p⋟PvL}Z�7[k����﹡$�������G����F�<�8���4���H\2ra!�K'�Ŋ�y�4A�qK�,���914R�{�� +-<�9F8.�~Y<K�'�Y�!��@x0(�)�������w��m�㔧D�T�U�Ң&�L��s���EA�U<IPH¤(ž23���#���Gr�F�A�T������͛7��}�M�����\ZkA5�$���'n�T�Tk���\��~���=��]1�gWnތ����Z_HG'	��.WG�'��R]��c�jv��&3������t�ԉ��DҬ��u�N8i���%�;�n���Y��(���Z�ٝ��F�aF������ɋ�y��������(,y�w,��awX�;V�������I���V�ɸ���V�u�X�4g���?vo���Μ=q,������E�3,J/	�@)�� �R<�ҠV-����x�����t�i�t��~�G&���Z��Z�cZ�iȻn���eI�xu�28H�u���0��k�tP9��w5���ǉ�N�-�.M[h�ܐ�����$�v�G��F���$d�5@q8�R�2�����v��g*WL]���ю����`�6e�+\�����1�(ǡ��D<������b�'�]���G�T�øH`xjr�{�`��_���T��,f �U4.���`BK���d5�LaGQ6����w�R�0KA۔ż�4�k�ɳcY��~��*Df85�� ! �E�Ғ��v�Sңb{k�8����	 �P���3mh�_~��_�2ݮ,�$�><��.Mq 0��׫�����������:�Z��9.px�F���w�+��ф������t�rc�&"f�+=j�iL��y���\I�M�?R���#��+0��錸�����_�%a���Ԕ�������/_������� �NF�^��P]	%@u��ɬC�z�,@�+4Ռm"*����`�����R)Kw�Z�gF��kzeZ���5>�QN����l0�=*_�< �Ǜ�Q�?&A����8�v�(g8'�S��fl��k����^����9�C>���\��*Ä\��T��a���I�s��*�
%q�S�� ���x�M[�����VXd��x48p�$#J�C�'&X�y�m:�EZ$vfyAZrI������Kk��V&��@L���p~�5Y���%�&� �Ytf5sV2�W���.��=~�`u��������MOΞ9�b�z 	(��p�{xK5�.�I�(W%'����l�;+�}yr(
�RźO���G���/<���=�FεoK��v�Ƥ:�X��'�<�"�h�'����wF��r�h�y�"���ѡ�rh��K�'�gsm��J�g��;�L��$���Tt���ͳ�WiJ�˸"��� zꩧz���H�)�uEz^�P�G�G��P���|l;���=a۬�TS�bB��g� J W^���{�	�k{V8GZ���1&�5����(Fu(��r]�!�|\h�*�Zg7tB+;2kң�_�R�N�I�?�}߇տOZ"�w��x�	�tdK�Ϯ��(�&�ݦ�/(v/�F���T���3�/�9����	�R�����O9b��iC4����Ve��},F�4q5���B�"� � ���L�B�"�=�Lt�
��1<9�=�Fw���E�����e�.]�D�eÔ��0`q
h����$L��������;�� kXbɚt�F�&NB��j���Q��q���[���0�H�܆�(40�đ4&�r�
��m�H)�r9_6�$�k��(
@^�-�����f}x��O
���e�W�� ���X�v�]"���Νc�ߔ�����+.:nff��I�}�Q)*�W�a�~�G~����Ͽ��q4K�p3�q1� %��������Ϸ�2�d���A#��|e����:��z8�WJVop���o��jb^�M,6�!�w��枣������G�G�;����<S	����;����q�����{�g;�Cr���!
VZ�=*"9���udx[h#	��� [���R����n$�7�u�Ld;њ���Q�*����u�q)�\@��ѡ�XP�k���C�#�5̷�	U�g�,�)��<Ŧ�Ҿc/�Ü�Ja�e��A�(ѭ-n��w��}�99_�{*թ2
��xB�2ս.Iw2���is߫s��:�s3��f�fB�Q�����L�[,�ه��� �$Αk���B��e��9W��z�����U� .���z�[�w�� � �Wh��Y�RoO�nm��D���$MB'�����z�sX.�ժ���(���3�=�d��D_il���A�x�Re�.�(8?���`����hB�4Iť�Q
�(H�=�=U�=���ͩ��bg0�c��qV�;�["��_·����pX����V#��.���;ol��'p�4N�/�B��$�S�ZpS/
E�&>��-��A��ׯ�9sf�uZSS�.��<�no���%vR�R��pR�6�^�Xȸ��(�$)��D�J�·�h�&O�i�J�z��S��(	D�o��D��h4,�^>�����L%�\7��qK㭓�??5_��f��g����¸���Q��r�w��A��T�c]ֺ�yB�T�� c�fv�����v��1�룡3=�?�[KƋ�F�^���k8�����k�z�_��t>ǃ��;��yA�ޚ�[;úX�{��p|jL�6�sXJ4WCMâ<@��%�>��L_u&�s�Nsއx)V��q��_)תA�V��Ozn�X�iv�IS�2��6�t�~=�e��%��Tg����T�`k�}�sT/�R)�rj����ظ�������)5����S�R* ���E�F�؂r�2W�⒁KZ�̗�9H'֝;wp#SlC��Q�%|�1`�QN��]cB4�[��ڂ��YY��L��c�����`�r�vu����[X�e���6����q�iG �6&�L�w�]�(͈����κQ�X����Ԧ���O^��Y_ߤDfS��i�Ð��s�t���S����T��>�"^`�\h�bU`�6��ϊ�*V��h���Ӱ|ce" GJ�J����K���'Rm �����gǣ�:&a������o���kcG�^��Ub>�
em7�a�����g>�����r�	��0���2g�{Cr��Y��3����sDŒ�����#��?�1mI[V�]�^��_͆D�jX+�!w��jq��o��o^�zU�r����!d�鲀k�߿�� ������U�h�m�F��,���F�D�P��DA�PN0(l�#�T�.Xޢj��2S��#I������^���9B2�t��')g���# �Bz�Ʈi���ܟ�����2fR��t��0�Z;?�c/MM֢={/�&��-z�ԩ�})�">�9h���u;�!��Lo ���,��m;@O=��v\�cw#�����@(���[L�/�"�ИJI�-���R2����f �'G��8��Ԫ���ģîvJOHDDc+1�.�/�l@� ��������܂$�ֈ�d�y��(8{�$M3��4G�,Q-7�ն�L��3O�!��ٳ�<�pjA�2ŁV`M�8#sq�@5�SΊ��#�Q��@�f���ō_O��(�bu�"D�F@I��Dz���UU�W�+�O��/��/�Yf�2��XhgmY2���`Fs��^��M�D���.Xۈ���uM5��KK���G�<#)�@�6�c�
?��H���P�/�����^^�����|�E������k����W_}���姠9�����14�z��7g�sd�b[ZZ�3;&9�7���/���u����reA�H�r`wH�cߦX��:��З��_�p����W��O~������C�wan7��ԟ'�(WwB�ggU9&�#�2,���5��W�)� c���!�DҌ��`<����v̌��{d"�4���\���a�C:���W�8y�˦Y=s�''�`������E�_ƥ+(k�	�
����K,
�;＃�2�&�֥"�`'r�>�c&Y��jb�7+�#m���/�������O�8qL���0���FG&V
��UG;Sڱglpskk��ٳ�B�=��s�,�gT�L�"���x0��v�����ږczZ����y�	����>k-���Çkx���9b-�6��m�59������i��hgg�th���K}����_��p��#a�XdJw;C��:��ƃݸqC�]��!뀌��~����ƛo<��s�L1���4!+
�_a�������������H���,�c�L)�ff�q�X�(`ec�������݆�-S�TŬ�&��l�A�ޔ��šD��M���7<}�ԋ/���[o�mj*��p�~h<�3�<�����?�������.A-�o��.� =s��ex��f��bI��^0XI�#i����	=�K�'�&� �zj5�;=� y��h�/�kj²�Wϐ_p��:�E���'�|�d3�k}�%�Kf�Y�Y5m߱�lXmHW+���,��>�}$�*�y��J��)���48uKˑ���C���sC�������SȀ�O�8�$2�q��	0���n��M��)�;v�I�xJ���*�Q3�.M�@�rBj`�t7pB�y�]��=3'm���t��v��.�sg��lss�f���tD[���~g���f�������85�Z|k0*�"bL7'�ǐp�����W��%�Ğ�F@ g~~e��X�m�����w�g�;���؜��q!.N���!��K�v��}����VH
�Rs��z���)D��	��p��}��PR�fԫ�������$���踍�l֚StFI�T�&Q"��r�W��s�4���6��W;�4�j?s:P굵)��IЭ\.:�'��;�nO�j�f3�&gϞ)�^<�����M.^
H�(�|-l{"*�cOĞ�"���R�/Tpܶ;;qٓ�$ix) bZ�~��g����<3����J��@���P�<uR�_���m��h�I�wa���T&U�fT��"�/$�,�Z�&��B I��{�Ὧ��⩹��^2[.��0������$�Qg�}|���։������ob��"i��d�^{�/��%ظ��y�;��sB���A#,H<�?q:���+�ɑ4gV���C��u�^�����)a4	.^x�c/�o�*�1��p4Ll-��܂�Pܹ����S˥���[�������@���]1�}�	 f;>����l��hW�)�&lA@��c^�:��$��)�����u�{�=lB��s���}H�QG�)��{^KO�u).���W�!�n-JF����j�S�<���1QB�kh�i�]�t��$u{����gH�i�7&�ҖeVI�q#|wuuO)��+��,����<Jyߥ7qzZڙܺuO��J�\�w<О��d�{��!�]�[�+���{�l.�v�f�FI�v���%0Z[[�]z=U(�)�R�Eߗ(v�^�����V0oP��!�b������F���.!V&��N�
ݙ� }�r��a7�IH����adV��?	�X�#*e5�X82��/��/�ʯ�
�@��ح������'���_��W�7~��~����I��u�:�z w�3`��L�+�1��ݻ ���p21$|j'�_Y=t1R[qX�V0=���Ah��y4f0Q����z�ڵ��~Oh9i	MX�����ǰ?��/�o����@�cJd8M;���4�Va+��!�g�1�'"i�3�8�l�$3"�J��[�
k�6>^Q����UL��@\�cT�8Y��
�ar�e4c����P�-7�\��I�/��5�3��-A��D爳-b\��}�Z�6��R�TB�H˂���:�C�dS��-��q8��ŭ�(��y ����;��`����M	(�% ���ͺ��y�a?��ᤓ64�Qc�#��(�c~��`2� ��P"(1��EΝ;g��W�\�]�C(/��6�`�v�$�8*�ϟʄ݌7!�qX�b�����b{���b��6fݲ� Pc�ߵ�8x|칓'��7]5��Eֹ�f>���r,KAn'��z>q߮V�O�%K �_�{1k�D��t]*Dxf=�+^�0�:x����W�չ��u��Y0Q�(ɹ]������s\6fv��M��`�K��>���~j)�n�i-��|(l���%7�Q.���8p�:�c�8���$pz`��6��u�yH׿P0~�Z�{�(���G
�a��^0蹎L�>��)Y�]�NX�,��2-C �fh�k��^{�ޱE,p��O?=5ۢ�p婧����w��pO��Wn�e��3gNyu��7�XVg�ӕ.�C��*���	�PVCWT^0�g;$i����pJ�b�`��>�l2����={���̬�ܗ0w]\����� BL3�Gh��.��ߤV���eq-")����26��
�'N0�}�9Q$��ժ�R[�#�#C��1U��T�D?�|�Q3�ig0Ή꜌v��x=��U�x����S�Ǹ	���>=�>%_��:�@��ؓ���|�}2����������<M��<!��Qr�b�ڋ�b��q)m��<��vr�i��#�d���r�����<t�cz�IxK-N`���"yR��heѨu�a�P�
�F����&
��߸q�w�zQz�
�Q0���XD�7�?�_�"��鵢���!D L`��$���?��ׯ_���>G�c����qԬ�c���ַ���������������!(�!�X��@<�^���
�cg�:��[3��L4��[�WbY�8��G�T��t0���� ��~�~�g~+-��S�����r+>��3��z����~�������AX���r
�6aL�L��{���uMoSC�pr���͖�"Qd�z4e�E�#�	�K��y��xs�,��<���RG���g�ًڦ��JN����11}����\8�1��4W�;���=?1qm~ ="����(���Zl`#��������hC� ):�"��:Óѐ��TR�i�aő����0�>�Y3�E�8�i����ٯ�/_&�7�/Թ=�s��/̸My�Z9�����G8u�T�c���B�=����"�P��mH�hw
���$���£xБ���҉S'G��p���ؘ���to�ٲ9���I��Y*�x��H9����D�d���+��KO<����w�-�œѸ�vE��b{u�v �2�䀑ܛ������'N^y�V�{n0W�5J��C�k�Lr(G�/co#iz�~{�����WVuu��n��n�v7��m�k`�F!,4�#61��e,��t��#~�B`��k_�c7vw��z��=��\#3"2c��y�y�}+�1�jUgFF|����9�ٞ�����ơ���[��g�dNO�'�\�j�u��j�B�$��=iA��I��T��
��f+U����9M��\N���`qa>鶞��G��ݸv����l8�����ηZM�'��R��T�c�l:�x]Sw�	���ȉ �D��Q����s'�Fƕz]E�����i<�4��q�v���A����叮�?=5�޼3�8�n�� ���o�T
�|�S}!s�,���|bo�	E,m�����w���+��r� ���8��eW6����;>p��Ǜ��:�rr|v:�c`va!n���N.Y��^於��dへ"��ϠjT>j�i7L����8���������`�_9�\��v�A� �clj���nǩ���c����=��Ҹp��h.c݃nT(���^��m��7S�q����:N�S,���:"���JJvCء��]�e2�Ɋ9)�ɼv�����xBNi�7Ky�iv6$��1?�b�Nj�m)D�R��My*E���
:2L��b��c��	-��W���`��VK��s��%���TK[f�>}ÙIk���m{P��eZ@��YAF�����<T:4�&�Y��3�?��S�1`�L	gT��d���6�O�%� �����U�
�,�!q��	|�4�.�q�AZl��@j::]�{�r�H���b�$ɐ��Ea�R����v�jυU��'?�����?x�������L��<��ED{�������������O�ԯ�ʯ,,�b1�DꪂԌI��ؖy��gg�1$�\������M�`1����J0�\l'�w���	�Z�<N�X�W(䨡93Y�D6�
 ��G>�����?�����゙IpLG����I��3K��g>�O�ӿ����b���I��q���\.�Y��|�H��o�;פ�sM��Ioq�!�aF�>Nwb��ņЕDso��v�ȆgJ�+�MGh�� aW9լ�D��hBk0"g$��P��#\h��z�:;�.ݿo����-3476Y�"<�H�*��q����w��7�?&圚�Fifs%u�tW�Gt_o�gv�}nwX'��Q�����!���b�Q"lu����`6��'b��@g��^�mL����qFl���Lf�ߊxt{�BJ|㱈��8~o*q���`�֮\���G�/xh ;#��0+PQ��[T+7�P�_����P��#����Tuu:b�N��,���󴳳���]^�E��ő��v�@=���p>��.���E�Kb���1���viT��D8��7/�M$�\΋����:�0f8V�'���1ظ��	�v�&y9s����롓h�1�����	�d�z%5)�C���y293���������& �ℊ�> G��X�!>�L�1�bN�(֔P��3�̆$��k\�L�H��f:��ŵJ72�ϭ�@�Y檒��֞ӭLb=aNX"��o�V"8=����LuE�3qWZ�HU)9�g��~I�f@W���H�����b?�D��q鐽S;qℤ@MMu:�p�'��6a޾$cu�R5F{�����2���>3�����Hb^�E������)���6��r3澸^�T�a"i�&�JW�<�x�',�7�ѧ�a�<��yԢ}&u�X����ڗ�<z�(��a�'�&2)m��1`Ɍ���k��D9�8�\k2�<�RЮ����Eːg���ֵQ����P�a*�Dwx�j����)cL�{�@���O,~�Q�|Ĝ!�c�#A���U�����a��e(��}:����p8��^߼�����Y�Qȃ:��e���[�B�ML��K�cp).Sb��3�)�VKq���Ͻ��O|�S�z�p�����I'�@�u$f%~��S
�j�Wϟ�x�"LG@�����(3�Үi���v��MF$�@�Yp�E��밆5W�U"b�oX=0Z�eM�M�Ž0�خ�c."A*]��1�����į�گa�_���h�iJ8�����C����P�_��;��;����1K�������l%��� C���ҖW#���u칦}7���]���\/n6zs��\�Đh�&��t+��Q������NY�K�P�1�(�){/�F�=���0>��[[@	?
�,H�F�l�1�y`�!�AځD8<�����ȭ��	�ۖK�^WM�� bk
I�����;49��8d}9������B��r����!ܻ�Ukkk�CУ��b��#x l�+W�`4�8��)�!���n�k��J`�QJ�V���}J��F�����7���I��Z���$���3�s@����Z����/T����}gϿ���_-��xY.^��/k����Ѐv<7&X�t./qeBø��߫o���_�77}��٥�����r��q���8^�������j;�>���� w��G�幧������v�%�Zmj�_2���eR�Aw^ϕ�ž��F�.��T[gQ��ci�. �	��R�8>�a��?�#*�����׿��'�������ݼ��
�!Y[�����B>�]���Ϟ=���~����'¹�׮\[^>����z��뻎_�]a��F��?��J�DY.(U�%ȭ�^�{��o�;��2y���L�ߕ����/�[��4�%j��8S����9ǝ8�����5漂[�(t�iInXq�/j
B��v8I��A'
����
��f�Ժ��\�9�g����N�ϹN?�&���V�W._�&����~c�Jb1sݴ�v���ӧ��|��?���{�\��Ƨ����Ɏ�"G�n�^Lw��m�Hٛ;��z��vq�i�N=�ŝ�͍\^py+<����{?8��+�4�m��-/�ɺ-�72Qط:����ٮ�P^	�X�LK�N�!MK�S	�j���E�Ui����c*t$ghj���+a�/��f���9]\8B�Q��oO�˜!�+8UY!��%ʡ"��&L�#C\07�qCX�b�������-�8�_�j$!>,��� bR73������x0	̡ᑤ���mtAQН@�H����]����|�i钘����A�?����祛sN��iI�à�������#͌h�P�'��'��r���M>8���g	��Ʌg.�t��2ρR�Z�NbY*f�/�5�[s���۫�j1i�H!��DIB�B�lWdfݟ9;c?��?�O��o�&@��S����s����j��/vu�'������{����>��O������t��ӘuQ;�	̥_�3O���������[Վ�ÆaĜ���,�n��1!≴�=��15���k�������̗��%��ȑ#Lζ�fDbq��`�������_����-�4�Q�a�<#�v{H��jI�+�9c���<�6rg�����t]�	��	�"N��5lp�+]�RE��7ҿ<3\��0c�e���$�(9���{�����z�T.9֤�e���aG�W�O�e���g"Y0l6��ӑ�Pv��!Q�L������oǸT�E�P�
�0D�T6�H�J�Ӆv���X�V(�����5�h^��'1u�����f/8x��ڵ�7n܀}��j�c��4��� lb2��
yVu�a����٤��w�e��:sZ�8u�W0|	O�ܬ$�nl�`NU�lә�x��g���bi��V�d���;�yr���� ���I��K=�Khr�_{B2ڷ7�h��ăv�1����&��������_��ҩ�%Inu��KϽ���R��
��,���ܑ���y4�\a�w�L��2��29{�/_����q�M%��R5	I+9��.�Z���B
��ej�؄�#��y	ݨ��P�:��%�J����Ɲy�#Ţ��׬�z���1�������	��֊���� ���ū/��ҁ�I��O��>�A��逵��/�8�K�ӫl�bZܩI�Ҡ/&��Kb�w%cir��v��C�~Ф3I���r +q���^�}��˩,n�~��	�%l��۪7�}_d�A��|������:	ڝ��l��{�ĉ3��K������ثN��YX��0p��\9���A ��{����cQ��|0u�O�4��RD���,%SU$X�:6A�c���V.	I�f7�(h��x�l�B�-҉Z���$Sp�yJ��?�3G�u�I���&���'>�c�4:i�Z2L,�S�͕����%��3S&R�Cc�0�'=�e'
+K�a) #e���j��tj0�IO�aP��2����#�+7i�4����&ʓP��8�����/s����YT��c!EP�U믢o�d��e��$�. ԭ[��^qb6 kZl�����!a��i#c���bJr^�i�C�ϑ0�:ﲣ��x��Uq�6%�P�nH�̓'��<���?��?���o��藥G��懱H�~!;?�b������?���?�����ϼ�}t��緶d��yJ��-��brp��� ��Y(zpФ�̦�9�3�%�,�Ń��؁$���î���J��3���
G(��ǫ���g1����̐��$��G�TR�̥�TR�^�}��_}�y�(����=�1\�"i�V�ᛘ M���S�)�4zq�Q�a�g`# ��d�S�/׺�,z��R�yi�W�jbqa�pM1��U��ؔUd�eX�����u��m�,\S�0|9�+3/f�#�i�0n���l�($6$���&�D�S��K�����[���K d0��ˢ�Qxz��l�v/l��,6X���+s��E����S%<GF>��z&�b��d�t�����Ƃ�R)�D|�R��h�(��9�4Mp����ay�|)>5�~
%kgG�L��-��dű�ٹY�-�׋ǎ�"oM�͵�D���ϵ�dR��8�Fd�c�%�v���w��ݧ�|�܉�Wwn���A�`����X�H�{Q����;�dG\ݬ�85睥0w��N�ݬoM��b>�@^N6AE��(���}�H:y݂�"�{q�Fq�+D���B��6H? �z!.�f7+�
� ��$ȱ������nuz�XÕ���"��{{H���Y�]��2�s��L.u�W��^��7?Y���-�%����t㶜�r+m4�����ۭ�3�AE<mP��R�f���a�Z?��X��8=��kV'�� �e{йa�[�F��T�	������O�kwvw�����9UVLv[�n��
^sx�,qR:,4C�b�;�������ݗ�rdVbv�8o�Y�:����Z9v�g>�3����K�
��i�h�٣Ǡ6ު�u76�q��3���������\&����v����e,-ao��sGo�c�=V>:��w�����w��ڭ�f/����٩��v��H���{k08��ُ�����?|]� ��1H��xn�L��sO�@o8���]��v}`�r@�`N�}-�t�%�	�>�������.���A�F�LN�{��
�����D�Ol�� F@�L`�՘�M7]G���"�4�yOs�i�P�ě������ZmH�K�VVrqx�!@fq�%Y����\bh`�M��@�!jk�x���xd|H�~�pY��h	�[����|F晥��e�[㎳��8/^Ĭ����Eb�Q
L^�<&6`��Vꑸ�b���E����b�wjb�MYN��� $�cx�z��-'��>҂zǴ��g�"\Y�B8�,u@Ɨ5��'\�Z.�,!u*�/����Б�|��g�y��0��s|"������\�v����69�Vڝ(�o|�]��ƙ����w�?�����sۚ�R� E͙d0&N�M˻k�)�p�g�3*���ݹ�|'I�DVl�A���`��OG�rq嵵G���_��W_}�ĸ���g�35#�?����h=`�������oal�~��Ԉ1��O��@+��HS)�:̆ң:t���$%i�)��ec Z&~�qyt��3���i��?��`j�i�#mIyY�1I�#��1~Te#/{�t�}����tS�MOO�T�k����Y�d��8>�pxа|��H>�"R)�J]�.����{���g����	�����O�8�c3�#��'O����f��Q�Iێ���߸8a�����c�Z魙����Y�ig��1Ņ%����v;b��5��4�v!�K ���p�_~��#2��y�C����{�p�d	S��f�SodW�Z�a��djׯ�%I�,�e*:�$��w �W$�n�dݎ�g���T6Z�iW{���^~�;���M�|���h"d_k2b������5;-y%��OŁ�I$��t{���/��~J�C �߇Tu�Pp@�R%��Fx/�S�*�2J�(��y7�������+r0��g�}v��8��&D:_~��83.(g�'��ؐ���?�?�����6�J�|w��ڽ>3�;B-�:�w��iuAKU�E���E���x��֔F%g�|��:|���߸��o1����767_z�%��Ǐ;�Z����Zj.E�����5���䓅1gv�����ƝUAW��ՑG>��p������w.bզB�:hK����x��\	��G��X��>����uZ!��9�=�d���n-;���:��Z�/A�9^t���f0�:�sD���P�+�;��r��G�`��9�LP�	fW�
�s��Q��0`�3��c(W�1����	U��B9V��]p�&�5�ɝ�Z�:g��v��)�	]ԁv0$z`�#+5y�9��q6�������Ǐ4�92�]b=S��Rsb#�9�Ed���	�HbT�����%ڝFA[����$��F��&0UG�B�����(����R�Շ���J GPK�Ġ$?����j�����$b[⾑2�R1�Ύ�s<,� �*��ᦤ	���R��j
+hk9��XD��j���>P��a�1�]�N�y����l!f��:$��+�qL7�G�K1��2��nczI�EL{��}�3��2PI�H�B�'&��:u
P�E��Q�Rm��b�7�7^|�E������)*�Ї�z�)��h�E�������2s�a_mbQ ��9�9��c_#F�I�� N�5������W܋��T��	a� g0�z聟�������m�5>�"a��$���aw�)I2==M��21���uk*7��c{衇~��^�A��J�:��͡2��f2���=�K�Er`�y�D�B�:��/�P�{85����~�mU���j4J���[7�l��f�$� +54��mf�,2¸���'%0����o����ì;�q�J�soDD��Vi��!�"S>,%:-�Ủ��3¯��۝=���� "��aQ�����2�}�"��g>ʝ<~bw�����w���w������ ��D�T��A��ǫ��`k� ��Í0V�ҁ���3�ޞ���ͽ}l�J����-���֮7������S�
b6��6%N�9s&iv;������wz�ۛwp.�ܽp�Y<{f+qjw�Vo
f�s[��4� P�ݣ�Y�sH����/"�Q������~dqv�F%iRZ�T��>��C���s�@�p�嫕N�NL��+��\�获�b�������ߞ\_�����_��_;�-H�c�"(�ܼ)�����G�C�~N��8��_�x!���lB:���S'��v�%�\�~p�ҥ�;��{�>��:�s����c'1���]���������N4f������-�O��������O�Y�qE�-�oU�F^&��\���}u�ד�����Jb����q���9��X�n��)j⥍�������,>s��Z���;��}}1�D�
`�t�}����&<���ռ�tGV!0=Q�3�<S�=�yOvp���*�ؗ�;�3�5b��4a����֭��x@�ݳﻱ����nHrUVkA�$Yo�qkrb�R�mך~Xܛ:2^(\���vr���Ν�mm^q/��[�w&��P�7�Z\���l6�gPߨ���X�����ZZ�F��9//��W/`��������#؍7�٤�_o�����Q!�*Q9Z��L!��&���qr���nyj>K��Xy���0�<����,J��Q.��V(��,���@��n`�T	��"�]&�[�< �D�;��=���#XJ�F�I9L'��t�	�"�EĘY]��ɥW�x!F�]���LT�w����"��_���ic���,!F!��4+�:���� �u���1�EOاߕ���فV22F騹̺Ha��H1)�{s�p�5LK���gʭRC%��27V��P��6�����Z����(�� >a'�CVCF�<Ƥ���q�N�W�6ئ7��HO�J�f�ݑN��&-��[��f�J�b�i����r���e��>61���].��	(lG��4i���ߖ���;�B9�����R��[�;�0���|����?��� ���-���d��h��a�\�h�/��qV�I�Hiv�3��Y����f��}����`O>�$L8���:ubgG��<�c
�G=��m�&P[H��2���c���u]B -�Ő �ӭ���A����~闰���� �΂��x�,� 1	22�����i��_��d��|�Y��R�V��D��[#.d%�q5ѭ4����G}�X*?�tFqm��<O�&�%�����ί��Ӽ1�&�P�k����j4i��2D�gQ�4I}C6���|:�T#,
qp~K<wZ�"7R�0�>x��d�C��Na*y�&4IW��@L�⩧�����LyMj^~�ߢ)�_a������ �$�/yj_9hF�'�8�q?��a����ޖ�:n��<�tRvR*Z��i��|Z�+�$0��MD���ڵk�o�Ơa&�Kˇ>�U�aڇ���!K��c�|ǥ�iĒr�O��N�e�Q�x�0��2"m�~��YH=[3E�G��о腺�}X-��.�*�n��QjJ�`�S��ԙ��)`����ׯ�����,%���U��1��y��دӋ��b���8�����s3�4��h2�\���]����b�I��tRI��v6������?���ެNO;�f}u���(.,�@h*j�BIU��ښ��w�����]��7���V*ela�kq#u������όUw^~���cΏ�:=���j�������)�U!<+�1�����.E��2�mym�!*�6=q |([4I�Jmy��L�$�%���H�jy�*�x}����T��\�Ѣ��\�Z-s�P9M��ƆYY9)����f�H�����xv I�gWVV`��.�bkD��b�|&��$���ŋ�|�����]aљ���ؘ�K�5����d��W��<)�vaaI'��T4������3���n�����9	�4���Ea3~�;��z�yW����Ք��p�'��7�,1@YX7^�d��,b��T0�#O;�����H�����$T�`đ4�0r)��jk:�R�<d����a���mC��Pٳ�� =�MZ
�o���V������6Æ5���a�;wS��b���5��S̎��?]kr�@��n~"3:�虠>���5�VTrz)��#�%�dd���y�)f�?���m��g
���?��®,;�ژ��]�N�����4���;�ۍ9�A[���>�6��a�F����۶}?��5=n���-NM[��U`��1��Y.�:V��A:�q�l�~����_��W��՟����I�հH?����̗�|������z/�c��o�JW�[z��A�a	�NXAd���x9>��$�a�x��Mz6�%���2t�a�lB^}�ӟƥ�������.���9`b�E殦r�pՆV/[�1G�R�����ea��j� ��fi��>#�)�9bÏj�<C�ϗ*�G�g������$-��,���d����O:�q��8�oR����|�z�+8����(�.�=}�)Fj:,��y�O�)V�n-��=s̬��4����ʷ0��^��{nB�X�/���E��v�kج��鬧��Xw=P��t�ƶ�z�nf�=9�$�"�6�l�EE)��.Ř��<	H
�pБU��I��� �̲�Q���i�I�oG�hs�K�����~c�X��v�΍+�q,�<����J���c���~}i���Q1߮��NkC!Z��8ٮVe���n��I�N�gs�I��R��N���M�|1W*u�4�;�{�4� �L�z�T�	�>�����{aIr��| ��Bnl|u� ��b�4ӫ���>����	��D6I�~���na�����~
�<$o˛L���=�Ϭg)3�n߹���(��������w9z�����ר5��^�����CF�w������V����K��#����B����ְ��1y��wnKM�� U�u��)t*��pO��r���jX��ǎ3CYf����s"����v(Y�X>Ipl��a�� N�0mb��l�+�W_}�ʕK�3�S�Ǐf�`���^�w��`_}�_���s����N� �����\�B�޾	���t���f�u���ٙ�����8ބ����Z ��	}���ڵ�����cC^�zE�g���4���
��m0f��eo�0�0Q�O�F0������!�Y����z�I"6,}����I*  ��a��cL*���W���nzl�^�3�jJe���ia�C������H�hO+�(әw��7�|ǴT����T~��%����lk&�C�h�l�p�kk{�.�ywm�?ٌV��
A�n*G�Yt90m�w�Z#�F�wvgbX\}H�c
?�����J��Ԑ�{��31�&${����+R������Hdf��&;��Du�5��|��l�ŨC��,��F��*����T�:B�Ҟ��<{�%����$MZ���!4��|�~ҟ��"#����ey����r�S�Z/*ZIV�@	���:謭��>}zb���O|ⳟ��o��oI8��Id#{;�g�.��ב���ʖP��ÚY܅Ŷxi��#cO������T�y�։���d0�}C�x.OMb�E��||���4��9>>��O|������/���^�p�I(��l,\߼��nO:�[F�ɜK�B�Y���2�ε�����a6�Hp��5 �E0��6�v����#��x˾�2Ð���c�z���a��� ��z1������������v}�`��\/��2C����������`�fa8��F���崁C�����v������)htQ�?�_�1�>�:ǎͬ���r劤�h� ށn�krZ����o��,���%$�$PB-H_�r4Ũ�D{9��#�f�,//�a�4�5����/���"CdA^�z��58�"�4z{��ׅ�"vab�$=I؅�?z�Ro��f�-�X7oJ�N}S2rh�j�)>f���OeV$��Ŭ<Q7��:~�x`����pD�pI��A��w
g,�A�����Vv�N��V���x���$G��J�n1	k����06q�����2x��|�7*D��b�Kx������K.�*�S��_<�oۣt�b`*)��(%�U�DQ#��U�f$�%���*n�JUR�ݔ�#�WG��a�G�5�/��"�?y�k�pGHU�T�T��xШ�$�u0?���� IToZ2F��F�*!���W=���,a3��;����`y]Ɔxgjr������-,�K�|O��pr&q�'�3Ş�?3z�9�f���\o�i\2�V.�X��t�%|q51T7�(�h�B��/���ź��  ��P���+�ANN����Ԕ���W9&�
d�K��*���,Y�&��y���8�f�Tb�=��X��m�60(�^�g,
�>����M��"k�?ւ�"t;Y���ˌU�K1�
��Y��bW���'O��i�9d�yf)=��/M�f�T��d��Q��A�t��glX(����s��k�:ҕKQƞTT�떖=V��[����9Tf����tr�a��7��E���	��ss��H�qN�ޡC�N�ܾ���qZ�g	���/c�f����w��a��T���Yʺm��0�],�=7 L�s���/���������C��I|���S� �sKtB�j�t����-�טm��u�r�|��S�P\z��Z�.����z�eM�nr�����؂X��/L��%��x�c�?�؃>�{��{����!�'���ɐiZ��%�k��tYV��=�/bc���ZO��f �C�[�#3����:���G=g^g�E!���4���y�����O�K�]1pL�$g�%��|d�f;8�+F[���n�Q8e�������3�.�&�q2C��0�e�6w�)h��q�7ŤÒX���	R{nB����}x��(%1���蘭Y[�og�5��:�>]V����Ge9�;l�Y"@ B�S�3����>�,uzr�{��K�q������/�$�B��~^���[0�Z�D�y!����a�MV'{b���w�iӞ+���	wTyqp��@{����F��U����"���������|�Mh��>xS^��Ji|v&�r��~yA�P��ގ���{8QQ.���J�����s3�J���������+�6v�Y� ӫV �1���^�9>�(b>_,_oܨ���d?*Lx��ڍ�~X�<@XNZ��E;�;����+ЂnȒ7Vo��18	ݽ~?RU]��_o�����P�ҡe�#��7)��8�j����!�˼���l�Q��~G
��"$����Ʌ���͍IfR	�q� i��!t_��n]� Aj�R,���� (�
ve�䢡���W�^����y�<�r��5�N,M�;�^ws{��W�/,�M��6���n����ͅ��ТDՅTb��G����*�A1O�GpaQ�V_�41QVn��MZ���,���ՕgR�>h��q���5�"6������byL�Y�ĳ2�hޘ��܀ӱ�#	C
"ͫlh~t��E_�������I�̉'��S�(h�BA�p�H(�*��ݒ�)`	��D��Cz��>�fX� F�V��B�D��3+{�pF��_���`сP�t��)�x�Mj�,�9�P�5���&�/6��Jk������3$�bJ�u!P2R�kEi��jSz�1����&�Vr���Ta	*�W1��0Lll����	p�����aV��L
\��S��� B��$1}��t�jg<" �7Z&�0�ʉ%��:��'��Ů��I�#��&�0)��t�~����~��T/�t�a!'˽�Wk�7��6P�EA4l1U��/
v��&&��� ���ؤ����ܯ/��9�߁G���x瓏o�oMN�w:�J�������������7߼ YgVN{�o�Z1����C�'36���IO��.[f��l�L�'�j6���igR�Qr���E��Bߴ*JMB�cy���ϴ?bM͑h�}���bj����_��C����\�@��֙ad ?mj���-p� S�mh��	�l��k�-J#��3��7ky#/y|ɊJ	�9R�r���<�9H�~�+��#g��v`z6�<���7 ���TH*c���y4����W��	����S1��ץQ��D�J�uKnƎj�f#�"<r�yܽf�-�r�]���o��\���	�b���⇨TN�:t��/@RcB�Y����LA��J.Nݭ��^<v�X1/�PF�����b�|��u	k��8|����$�ة$��h|[�jj�*���C6;=+��A�{5��ˈgVt*��(71/�p�y�ZY�x�z���ox��\�^_�SQ3���
��u�9������������LS�Е%"c�Ĥ�ax�Ä-Z�T�� D0K�×.]"f�S�J�n]���Z=�N�V+,��Γ$�D��|��'�f����y�(��P����Y�'i@�.5%#T�ҝ�R!�إ� ~sk p���!!��Z�8%���ƣA$aA�I�#�=�&'�%�)M)�[�6�	fik������U�aK���3�LOO2�����W���}�cB>s��m�����a||lbjlwW����ڽ6Lv �ӧOW���e2vj��QL�o�I����C,���Mf���X�P#R�R�cE�.\� �M4@*HV���I�N6v��˗/K@��=@
�)�Q�7�I�z3�A�h�TB>�K;��yֈ��q�g��Ƌ��@:�T�W�E���m�2SC��U�m���7�k�'�P��e��B��W*N|L6�
8(�Tx�� �_$�n�X2���	���d%�%�BǠ�̕��
�?tl� vaaþr�
�/�Ε�yeBJ&N��KC'V�y�W"$N"/1�\A�^�7�	��6�L��]1�ŃD�xL�;['YuN=G��5�w�>�ɌT�*�CQnD�����H7��5FTu����8����1�! �R�+�-��ΰ����w�O��`�|��v������dP[��)�� �i��n����~�C?��o��o��o���/��2�m?b_j�F(8����R�x&�iee���/_ß�=�Ms�ڍ���P�=�;���JD����4�	ce��1���b��ܹs����/����"@�*dN����������ZG�r��Y�7W6�q"3Q�xq��+��F mGλXPŹ%�#^q�kz9&��i�d7�cR�|Ө�5�Έi�5HoN<l	�wyˆ�Gw�/�z��{�xL9�Ǔ�NS�I��f#�;G�?�Yhx�]����A��˲�6-�HJ��(�};j���Eg�֏g�0�������j�n/6��pd���v���:VA�IN���]�'��׌4L�Mtu5��`r��~��|];{N">��E'r��0h
�-B)�P}��k���������f���vS'[8,���.?),�� m�v;m�"D�s�ܠٸ�n�sQ?���\i�R����=\��x9�I��P�ÂJ`���^W�]�B���Q� ^�T�셥
�Y�c�۝�\��+� l�%��pc_4Pe�X*U���N�1=%�	�V�ixi�& GȸR���q~��b0�m�����L��X��~�]���Lw�R��ƽF��h\_[�.-,��` fQH*F�N��A@H�8v�V�������9i�|�������<��+g�T8M�´7��eEK� De�f���P��9M[i�Z�fSh���%����#[��k���W��92���d.~�qc��W~F��(��Ƨ�F�X�DI���ON��U�Cb��v���*]�y��KW�0h��xH��i�M�AGy�B9�	��:3���mp薀̘���L�_X��ޑ*����NK��{��M����'O�X+��Ju�h^�Xp��K����d3s�W�_��O[Q�1��ZV �����F�Z���Ȟ`�z��?C%�W�a�dv�4�Y��'0���5V8r�<��O�)�ބ�+` �9?��J#&�L>�,�,�K�!��l�4�ID��ӛ�͆�;s��%5�(E������7o2��)��Y�߂�6bMz܁����a����.f����S��2��z�\z1�ja0�Q��@l�`=1�sVЖ���=��#"-jA!I^_Ǌ�<N�:�L��5��E��!]����ZZ�G=a� �Ը�"�:kx!?5[r��\�N��؆�w0E���4�^;NT��C���x�������d���3+�<�̑�G�w����$(�h@�ƃRՂ�l$�"5��\���� 2�
��� ��܌!u"]� 9�L�!�5�{1=N\����3��i
����+�1��������?���}0T���tfڡ�Y01��-����hk��:�����T�P�"[���CS,آE�j��8��x(6�b��� �{��Ӓ$��Q�[S� ������OgXq����gѪ�ܓ'Gqa�������n(věE�iq��Jڹ��7��.YW='��EoQ��%��m7�����y�~8��ۮ�������/��!��>�����3g�f��h'��F������.~�8|�0nt��zc�i��#���d�r�3	��E	�XI*�q����Fx��)|�1LK���ζ8�P��ȫ_��2��, 4և�E���b{N��b������1����OP`�x���Q]��ЄrY���N͊煬t�%0���gV���wB^�~��B��4��g�tZ�m�"����n6D��i \�k��EJe�����ի�$PK���$����6�5V���@ߞMu��1j���O�&�ǁ5�9\�������֏�#L�|Б���o�۔��6L��ɔ4��$�A�K�X*[�Y����꧅�y�Z��|���KO<���+�q-J�T��Vs�Q�$�GX[[�M���N����e�+��88q��"i?��8n�T$��Wv���9~��]5����j�}�{��;��k(�<0�)�Qq�]��C����YU����6��s�T�tC�������%�4��
�T���t'0Z�;�����I%����19�P�E xa{j����j�S�	��̔�?����uH��_�t��-�I`/F����Ďi��⌐&��bm��Y��9$O��+m��Igŕe3�v@3�b>).K/�����ƝԂ||Oy=x�(?�ݪ�F{q)��YO�F-���$*
��͆��9��V�@b�sLtaS�nj.�CX/�_~�-�s|������gC�>���f�i��\�M�o�>5��^�h��h�i����)��za�O��G�6�n3�����������?��?���gz�8���0�n�h��l�@dd��:����sgo޼�턍�3�c��l'_{w2�.:2/P7cJh�X�
ݢ�a�O5_���1z��9-Q(C,��'����|�+��ַ�����c_�9#�u�!�]�c��]���h�t�М�А�`�����ˆ�A\Z��.1g�;�&hZ7'�79��٢�Q��
U�D-X�F2����"����f"�-�e��c�͞�!�-�����3lCw��SjZ��e#3�x�l�wc��u�A2Y>�/b>��v��V�1��A߆�\���m�7��`��������;ϖV1e���6{HS=C�CD�0P7���z$V����'�Q3��s�{"��-�� � )X���A�W�޼O�95gq)���@�g�Ʋ��;h$Y�[���j9nnւ��]%��ƽ@x6�[[5\��Qɏ�x����\�8>>����(���=i.�~��"V���R9f�h���݇�����J��D0bP�Y>%��	>�D!6����S����~$",�&�������e��C�����+-���K��%��X���_�G�֮ ���Zw�oc�1OE���nI4�X*D��ݾ��A#�$�
s۬7&b���1�ܹ����)�;u��II1�v��������>
|�"� �\�&u���\�c
(�����k3u�m����aEs����uy�r�_��){dY�6�:_�XS�Ç���* ҈�ꕫgϞ�����[P�P˻�:����$�C���]_�����v�,�>h�?����?���������R��!���-5���^�u�,� R�v���<�H��/��r�u|�UV����~ 9W�D���-�Ad�݇��w(�� ����`~�ס�_$=X�TQ��Q�bn��!�SF`�>x�ҥkd�`B�L8��K���"�@��ش�=s��E��"���.�JLr���I�Mf�)�k�$�V��Z,����-�3|�O��^O" &�a�����N�@���U���KR��a�x"����cl��1�V?��:�4��P��
ڢ��H�K�LS������x�''^�#��0�4��a�6p�!
�ܰ�U˸��"ʄ�Єz&-�Ȍ8�f��I�>�H�\��c��URB�9��
����z�<��ɓ����d5�U�����r��Ч���(��14�Y�ݭs?su�\���CN�>� [U2)Yh�76 "��K:������o�1@��f�?�S�x�O������?��7�|B�,',��4�/
�b�@�A������+�@a�aJQ�0�#j��:3i�T�-;c[w��I�BH�w��%K0�m�V�z#9d��Tc� �ţaKЧB|��|��g�����������k_c�5#0���e��)����*��a�S,bKHju^�"S*�a=ǐH�7%��00����_�jd&�f!�T���l����ױ3]�oz�Rm�LC+�y׿�JLf�wn��<�!�Z����.�|�\C�#Z�t�X_=X;Jr�B.klJ_�։�C^�ݓֿH?�c�8r‒|SV�s�b@��C*��c>l�a�x�S֐��\ˆ��4���\[[�^��;#5��tqq^�I�p�����郡��J@M��L����� ��~���̦r�U�kr�P��B�Yլ��ˑZ�z�t�4���d5�D���m��a����@�k*n\I�х�Hs�Di" �u4�k뀲�v:����"+j댶,���e�jf~�:3�_��h�@)K�� �h�nmJZ1�H��k;[*�+߼�&$�C\ĬXA7c E�Z�M1��odI��OB?�ܲ,+��M=.%�V'S���bX^��j{���Ns����}�n�ŋo��	(:1���niƺP{��H.2�0�Q#b�~���,W<I��Oɰ�c0$)̼z�M�J�O]�rE}T3���a��B�M�/_� I㉋HK ��ǃ`_c�9s�uX�-��~�'�=?�d�5�th����]M�fǛ�4l���݌��0R��3ی[K�QbÒN����AR��.��uvvN3�żף=�T@��9&�+}���Fb�O
{7�$R+�E�-L��Bc~��۩k� ��4�q�g�E<��tl�ƹ���J�MY�U�ըY�'&==4�e�$�S	�-�����PlL�b���S͎��V��Z�GW&� ��K�l��<���DVc�0T&����-��SM\r�s3S9ѱ�٦���~`�w�c�u4C�L�&��ګ��L1��A3�D԰Q�"<}ޱa� 3v/��؎�.�/�+�Y8	��)�^ZZ�x�f���Z%3��&���:�a��X����D�BU����-���,��+=�����!�?C�=Ű33ӟ��'��w@d������/��{ֳ`Ht��þ�tA�NӋG�u8�V����ީ���F�^Z/��P5�%�"�(�z�7e��"T=Lk&`r$�	7?�K�Դ�B���3��=�z���O?��o}6!3h3Md,h�6���������,�[�5#%�SSt�$����K'����X��;d��|"|q�Q�����u���L3��2��]M�i�<�Q�&i�[60]"GHv<���>B�D{@�֮�M�Qg$��Ih�ȕ��e��FS	yM�Đ�×�Ν,��1IO��"ܱ�'�a��/L<B���;#os�qЮ?�|�2&�b2-�֝ۻ�=l���Jf�*�1͍5;�BaS�b!F�&�G�UJEBw��z���~��W����(c�#�-�P��rb�Kq��T��l�v���b	�a|�"�<[�}0W�8Q�<k�j�O�y�N)<��n b
9ʾl�9��ר'�ΠպoeEP���B/B�M����Kׯ_w=�~���|XJ�;n'۷n)٘�Ms	ήݾ.*������v�^�� ��C���^���isoobbj��S7.^��|��=� �#�y���}�@�v�뷁 :��Y&|�����X��NMgI�J�qk�;��dش��a4!��k�v�|I�e��Mک��OO��q��Y�q��W�l�J�\�>-��؝ %Q��QݺqS=p��Q���W�e@�o�h.�$8��:�YQ�'W\�έ[� ���o]|��eeeEr�����L.����j�
__��B���姦�}d��ظ#d�<M�t���J�I}6�"'�!VGHL:��X�[��kߢ����E�a&��38�.1!#[$1�$�o��p[/��.c#i�dY�&V�<I+�q�8W�q��N��HU��;t�Z��V{_s�f�M�g6c(��+J���~�D���pe����Rr1��z�J=̞�DS2jv��h@�Gy��7LiԔ�6�#���D�ii�ҹ�iIZ�T�ʞ�)��QGl�"�K�@:b8_���E�î�h�}!���|-���2�ӕB?�oHhi��3�F�Q0��C��vXT�y��`y����	1->ch�<���X(��b���'�]��3��cB�?��C4 �DZ�7M��������I�8�M��#�1�$�̜t_�{��nw���<�$��M!��	<wwg{�\
<���ou�X��L�H���#���`�a���� �����7��ͫW����Z6r�#��9�Wb}���M%�]mQ��V_Z;4,�v2%F'�f��\fr̹1lNvf�~��j`f������6�Ѡ�gJ���l�{�ı_��_���?�-1 9��@�Ѝ�ϼ��k�8l�춻���=@���a�5�1@����2�R���;�V�"$z�[y�<���Wr�N:�z����+��{��99�pg�����3=�<CT�ޛg6�.��K~����s`�ɢ#��+7�Q<J^뵲RM�B�3���%6�����:b&���a��Ӫڴ]��d:�}�!�4@���=�43���or"�lXx,]BC���$�*�H�1�/$�:��Q�X�L�e1*t�\S�8�N)�����KA��z`����̐��v�Q��j��%�ͮ��L^�2�	=V,���E���l�Z�S��
���.7n�"��#%)U�n�����%�l�r��������,-��}�+_��'&��SR�����{�S%�&�+��@�m��� ��a#�,R�rg`7x��Y��o�C����:���K:":iݑ�X���zknNx��A�F�x�Z�쑇'-�KxX���v�ѭ�3M��3�ӓi� �tA�r!E��*0{9������߃��^ĸ1=.Xq�!�Gcd���w�D2=3	˛ ��p�qfo��<��
l9�OM��Q�в(a�>�It���U�����8��ҥK�fd�Zu\u;}�ax�nZ��)ӉfX����'��������y>v�> ��f����Lzc�E�EEH�r0�����&��3�v�A���<�� #q?�-��\S��3���C\��'5߱���E�2�@xF"K�"�!̏Ǩ[3�mvNqOR��ޣk�Ur�f���u#�`�а���ȴ��&B[�)��ćb+'ͺ��Щ@%7��X�G�3KO(a�>���l�g�e ؄�����t�)yS���D�I�;��-���s�^(ƚy�1��ݲ���L`�{���BJ$��K(}�A(�o⑹jx�@h�X��_R��~���a e���q�������K��!r����a�ۤ�����ܹs�~��I�}�c{��^;�*Ñ7����}wkg�h��HͲ�`�tF!3M�IZT��6جp�$��tM�a`K�HƵ3�c�l�r6�5e����W�����M��ɋ�t^|���/�|�_�W0Y_�؃�<�i�b_���զ�!fn>)S����Z�5e��k��tȠ��(m��5r��Cj�a_n	y���w՟ڷBX�J���^����(Laډ;��fq�c�2��T�;���������S(�Y2ޝ+E����QҚ�FH�ܑX0aVjH��B��dl�ZY���p�or�G_o�h�a���N��hO�4����5�o�*e�i��3�%���Q8�L�4w� ���XT�!%y�N��-孎�Q�P��P#�C�7�(ɨ�� %�nȦ�.��3ⱈ{�r>�=t{s]�RY��V�ՠgϞD�+�_�0��Bi�r�|�ە:��A��7�U��;� <���A����~�.1�����HC�͍M�.L\/ur^��	=�8~�b��
�f�P*�(/"c �=�i�._��裏�����o����|/M�^kF
�� 9��k�ݸvg���p��+��}I�G�v-�g�A�B� ����6���N;>����1��D#e��p��IZX��dy��I� Y�)ԛ N��w�T=h��7�nH�L��j�r���b�X(K�i�t��5�>��T��*4g���䩆�m�H��Ԙ�[0c&��9<37ͼ�R��;������fV�����}L��Ңv��)�-�23�sx�^ �'	Uc�+�Y�p�~�M!���ƊW����:��I(�|A\ kk���S��K��AH���5��gg%u��b&1M��	���Oi�4���n�g��|�)iUcղ(L�4Gbg�ёNG�J�CZ�d5.��>���_'�h)ė0b|�׆�D��&�$3܋�)�SL��fF5�L`t���T��Iƾi�P���^x�YD4m)ǉ�)(���&S�C�+��ݜt�V� n-4���0��)�c��>ae4�1Q�k]V��X��IR�0��p��rR�p2���Ō�0�M�?�U4�=�{���פ�'���#>��V������8Lfg�>I��­����{��z�C�%�W�Ӯt �4l��1������#$��2�&ʱ"%<�`p}��jSB ����g�!-��T���1�ɩ�b�xu�z�6�7�m0�m�Ǽə��}��?�c$C�{�ʕ/}�K���llZ���K/��_�@��2F�3U�`V3LOO�� � �~�ǔv����у����q��N��f�n"�HL���g�'o%ZB����ǵ�%�� � ˊ�-�0=+5�$��$���0�l��E�<t�3�����.0<���9����qޜi\Ƴ ��SZ_�u�t{��Bg�g��?�^��L���h;��)��)6���3ϐ��p�?�@�z��ҳ��`�؇�$i!��o����(A�E<0�u;Y�������L�;t�ϛ���/D�eq�C4�o�.�Y6R��$Pa�)���؂nB`1�t*��f��n�>��\$�+~ʅM��9����Ը>��$Mw(���u�Xl2C�JU�'qVoHWf�#!逹�B��~�n7;-Q��C�|~�iu���;�)�����d8)i�힤�?.5���0�B'3y�x5��~q��șS(�i��P�*��<r4�qqnvmmס�JB2�Q\��b�i��+i�'۱; ��Ϭ)hF�X�w7��K>>�m>0���E�,��ـ*��4vք�����p�q)�1��N�%�� ^��CYCӸ˜?Z�x����G�簠]ii�1L�9
wC�[�Æt�n	<&w��O�>ل��y�u��[�c�/ެ�5���9�gϻ�/%τ��0��NS
w6 b������{4��3��-�G�x�:-���s�
��_ǺC�a�^~�e|�����$��?t�t��xX�*�ɔ���s����#3yN�|M�R�ΠI����$�Q���c�	����"#h�1lFy��q�M�a鑅z����+6�A���h�Di�b��`5�=�����C,Y�$`��Ot�I��Fd���]7�z�*��0��n��;-�gb`�	����d����NGV3�ʊB�D�-�î��o�S�1�XH��'�a䂟�J ̲8�����d"G�P1{Öw����1Q��(	%9�ta���}�1*��Z�@�=}e�T�t�cG�K'A��/����Ç��L'"��}S'�S�aL)�%5��0����i��8)��R����F��Lw,�χ��I�wi��>5���H��H����ŷ��fO����?��k7�]6�6;J��pǥ��Zm�%��O�������,?EG�+�O�H(����ə���f#Y���e%��i�;�u��u���ġ`�.�Jg�߁{�o�ɑ�����l�$��P 4&�V۳nx�>^�s��q�X�ACӬ�5)�@8������0O)j��m�����.d�f6M�LH�٤EĔ�F����!^Ᏽ���4��f
�C�JmȆ�Lx��#D�'��nH�`G"]����؃;����'ł�=J�\�-��m�3���s�6GZ���7��Hb8��F��ME���ɀ�	V8ka(�����
�8JZ��I�3]T6t�P�DC3QY����d��)Ĉ��>,jc��ٹ�/�*�}1���N���NL���K�m�/����B~�'��#��S���^?>�-�T���qQ�P�͗�z�\��5�G�q綤Y@��n,1����Kc��]�i�UC@؃��s��v��~���R�T�E�T��q�w�쵶��g��1ow%Bqt�H��;U�X��i)���dq��Ӥ9hfn6>!�&�'v��$��;��X��c��������g�Ay}�v�(vm�T�eGT3��=3]�,+;Լ�Ed�5q�o|ڝ���$P�R��;wbL�	� ]mo�
(���),5.D815Io30�R�J�pn�㼳��+�S?{�ǡo`)D9�I�I%G�;��?7�����Ay�� ٝ�M���`��8��Z��P�;���ՙI��v�@���	Rꏹ`�l��w���<���Q$��AO���~���C�p7kw�-�������S>2�A�N�d+�5��I`�����F��E��(�������s�n?�FCE���l��'��ِE]�غt�Xf��u�b�٠���kGS�Y�i�h����<M%���>C�qM�
�DW]U�,�ݰ�Y�4����B���F���,.ap��?*|�1AN&q3��� ���3�������~����� �j�v3"��\<��D0��h������qY��5�L�a��i�H�GH��%�~3�ʰ��0N<,+�ZL&V��\,&Z��f\�	M���O� ���� žVb�R�M��3���%���֓<�XR��YK�(A,|r,Ԣ�u�YM�(dOY�xA�#ut�H�Tʗ��|V�{w�fے�O.7��'��	q��ƫ��A2�gά�����[t�rqw܋�*�W�a!3���a붰45���H��QmJ� o���$���!�G}��w��.�h�i��*�;�E^{�$R9;E#�`������>�o�N��4Dg����~a>3��ࡵn  ��IDAT�LI�$���oq����L�с�;����02��0���1@�LFZ-�� ֺ��a�@���u��2���B7��)���S�q�pbS��ŠʛC7��'�jW��/�ϩ,Mq}/gq$�μ�������Wp�/�1t��
���tla�9}�رc����@�C��p���!Ŷ8���dؗ0������&U�171�� ���d���S-�Ң{��Hp8q5(l�Ԓ6��T�y�-���LLO�0P4H���À�q]�3�_��*��Kn%	a�����k�|���#��=�(��g�'�gl�H���D��	BO�y��8�h�������K�?_o,�Y�����G͒�#K�5ز�cC p T��K*77	I*U�KB�J�Jȗ9$I�p�*���6�lllI�<��9:s��}z��Y���6��;�R��ӽ���a�gM�:z��-�_5?[�l���MdI��ƅ	�c��?�冏*�R�,0�������q3��zp#a�l߾��OO���R5�"F*�d���F�,���,	mf�խ���͛�˪�+�B�/���<8���+:�r�:z*}�����Hu�p\A���@Hv�M7�ڵ��铄��ӳ�_H"��!�L�<E��5�=��Sr��Ý9�����2<y��b�"a��oY{(�B�8o��6-z���$��ڇ,�����D��%%<h�m��S��A�=�)\߰{�3��LS�;��ܹs�a͹���s��ac�θ��t�s��S}&e���]Z)�s�s��h33�F7��߇��zQ��x]t��ѷ��z�� 9�P	�<8cccx�5����h�{�6=�E�c�T*h�4 ��<�E�41�-Q<�R�6��&�V�%�u��tz�>�
�v���b����z�)WpΚh��g$0�����"܉��֒ix���R[s�b�H��x�K�[hS���`�"�I�d]
� 	%6��������C�V�	������8�\@-4ݷ��2Z�~*-��ۺ�Z���-[�ݗAp\ãxVc`Gq#M��<v�X��c^͐:�܂�T�<�V��
��A#���ŵi�&}L���~�r�X l�/ԃ�lP�I����'w������7*)έ���cz� A��e��'
��J�z
z���"� \�����ϲ�Ȥ���ϟ���ρ�^m�)طx1q�`��u�UB�ZD<��:"� �K8�cyD+Ѕ��{/b��c���I*�������J؈�b
�t �|�Dn�v��Ţg!���
	sI(P�B+�B��fǢp` ��drd"���0Z���ƛ����V�d��u3�z��%Mۅ4�P}�m.�d�J��`�W�7��Wغ�,���kҨ�
���~m�4�4��VҼ|�R.ߺq��eˇ��کS'`U�l��UW�L\���������''g�\����o�Kc��ي{���|�����Z�v��,�#��ܻ)l)���e�����8`\���N)	i��[��x�}i`0_*�"�|�q�I��X�Z��z����YCui��-U:]kU�X���h��2��FҚ���ӽ�&>J�t`�<��؍�?�sb�g֢Z�V����z��՗�&.�5/��vG��[��0�Ԗ��K����V�Y}��ĳFd[���ūf���Ej��^4ަro�LeNo�j�hu��Wiλ��.^�����Xo,�)�bA������
33�g>z(���H�MLO��B�ZO�@���������de��M-Je���)j˦�FR[\�j�u�������B�x�������)���������X.-֪���.�f�
"��FBߵZ�޽�(d�/	�T�����U�����@���3�9��ׯ���ϵ�r-�%���^�0At��eJ=��Z��[9�B��Ա�##�C�2_�3v��n�<�iS�Ǭ�\G:f	� {��1�y�$��ӳ������Z�S��u��%�얷�� Ե����T]e��뗯�F�L�^sE���IҖ޹���3�Zeݺ��AF���|��jMLL�m���vǭ���_�Iپ}��ӪLf�\mL�5��Aƒ�+,��I,�FU�::S	Cst�;v��J˰t���3ƴ�<�y�;�iA=@���K�В�eP>	&�_5!&Y��=Ap�
�T�<t3K��!��'qM��,C?	�k��p��t'�h�RY��_ Bi�Q$T`�׹�-������HjD�L�.'�LP�g����;�� �zͮ -	rZ��r�r8���s��#l��	蓑���34NƦ���h��՝5[��S?v�����t��:�m��bq��wff~�ϙ2j@�����V-[9�Y���e��\�����)-����O�H&���R�������{��_k�Yu��ng�˖��ճF��.�T��N��� V��U?��iq��y_���������e6�ny���x:eL�P�'	[u�L
V�`�\^pp,�12<l}i��"��X��')����n�ͼ���:��ޜ,��"�;c/�:�z��^T^�ɽJ�)_�U4&fh�h;67Wq�e8��\Z�n�!�$�U�]��f-��f=k�}5Ή������^e�s�8k�#0�B@�
%4#K�\OB/�R�+��h�ig1(�ay*�$����n��ԓ纑$�UH����;tɺ�n�0�ט�]^ߍ���L:�����$tHB{uϨ^Іw?z����������q�h��T;νn�5k��6��^����[�j�����P,�J�
 ��S嬡f�����c��ginMC@��LR1HAm9m�^���ͧ]+	�y��D�3S{7޸w�+�\7�̡�ԯ�ff��x$շ��BO>PVb8B�O���<XΛ��nH���#EI-ID@��\,��������Ӭ$��l x�2���$�D& ��	b��N�u>L��X=˹s�*�y	��Q6����0�1�K6�R��A���ܼy3�&��'N���C�M��A�s����/#�;2ra�� 0ř�܏�O�I��_))my7=Mˉ�?I�G'���n�@�M��!yFM�}�=Dm��0�j�u�����G�/F�O~�����_�J=a�ދ@A�|��N����RҲ4K������ȕ� n�i�y��G�j%�J�`J�����O��OsK��nol��@�'�Q'GW���nq�M�N��.KGZ6D�$�R����xkJ��ۍ7n\��E�<-�ԙ���q���98�^����v���Lm��_�߇^�x�4{O��=�FEkE�HJg��%��m�x����$5Pf1T�e���[�l��r����g ��*C�b��j©��-� 9��bg��j�F�u����]q�'|O:&:vF�2�:��[X�Fhˈπ_	�J�A8��P�n@^,j��1
�W�M[��Bv��3�:�s\��H6r�3��| ,��J�JV!���,�A\D�`�vJ:��4���联,��@NU��J|�(� �.�.zG��4��D�%5�$��l��+N�G#r��Ãbanw�i�:2�-�ܲw���:.u���+
S��Pk)Ӌx7�`�'2 =���O���1�X���P/�a�O��)�HB��0�<��s��R�.��+�İ�L<�c��V���
l�b���B�^�%W�Ӊ�I!��!CGO�L�+��IfL���?��S�:�d��u���h`34���+E YȁKCa����r9�e�_,9	A���k���)�/S���=���/�X6����&q�IH<j������+r�[�Y|��?K;M���-��0�$���0R����|�&#���ή�
Բu���"g�؃�Z�s��n9PiSO�����C�}��t	�Ȧ��ѿ��Q
�)���q�Z,WW��]�Uϐ�#��*��`&TuM��t���a�w�Bf�4o�E�)2Ή9�����曁�pL���ٳG��3� ����� �Jyc7#�:�e��, (׽�<���=eM�����jf1@؂�Ox��/5���!6e3P#"��z
��f�v��v��a)Z�06���ӧO�նm�677O��~��aM�E�G-%\��(�ሒm�)Gq�<::,h�Х4ccc��0
n'��9y/X�"S��3����"����&�]��:�Ār��]+%���h �.]���ܞ=�����n�J�
;mZg<2)��ǿ��Lh�Y�2���c�4�ݻwg��w��0�jǎ�?����\�)�l븥^V�DӐ`.���IN E�V�7r�Zٿ���� ."O��PT��y14#����WBid��=�H�v|ǳ#�è1�h�{:�o5lcC���䄒��C��Hm���5aj w��Zc�����	��@��O�`1�K�-�@Ū /��M�̺�lĴ}�zE����x
���oi����ú�8'桙�(fx.6Fu#�g��Ԛ���:e د�Q�����QE�����|���s=P��B"�͆�B�P��ug����B�z���>�s��d4��:v;�P��p⢌�����Pl��H3�J��	��Ҭ�v-J�JK�v���=���v�i!\���v$0'��[9V�@~��nb�@S�
|fI�^�/�9��:c,��$�a�m�c���7^���f(MB�V��N�XL����|��{^{?����T���I����6r�0@-�8F?��iG�[��r��P��NЪd5�k����Vk.d�g-#|hs�:��6|���]S�K�%�
��r9��Lڭ�:?\��Z��t��� �?�d8�`X�j�
���7��馛x�J����|�>�4��l8�$�;�=��@�	i�Mo)�:fP�ժ�s*S򮿭-F�K�1�tR�\��8$�BE�+��H̞��Ի�j��'�o��)�\ο��t3lI�� X��D@tA�>���!�r)x$�,	uF�u9W8�c�cpIֹ�zȏD� ��K�Ŭ�q�U=��2��t�*F����K՛z��F'�S��^���Z�m�s��Y}�V-���u�rkO�G����/����{ot���h��>}V'"�.�:=2Ht=�k5K���XȦh��ҥ�$�ڼy�fC@�C}��-��8p� �.e����Xޛp�3D����[9O�A�A4k���$�D7���NTQ�?<<�m�G�?�$e�Ka&�=�@��m�ɣ"�֮-[6��={�^ck���R�;p��hB�D�@üs��������[����(:�b)�2$"�h����ҡ�qrd�n���z�KfW���aq��nb���Qy#dSϮ���͸�5`6@<AQ�qk���
���R�H�&�N8z4��j��:+W�..֟{�9M��D[�.��CNx��+���V�@���5�k���J�*Xʵl��������<�P&�FGIW`�z����N�_t����Dw|���13,.�ѳ\J����'G���ǥʳ����V��J�oKz�k'��Q{�-�z�
�7�,����jd��(�1�=|��P����ʝ��Fx"YMvl34J_"�)�����9�	��*�3�wV����e!+�`��F ��X�>L܇�vd��2������tn�6�N)�vw�q�c����TŘ�G��h���{���GDC�vQ��曹К����Y�uK�g�_/;��d�Q�^���Y���eEE�e.�0�}�,{/���qCD-����]�Ʃ�
��E�u�6!�~���k�j�"Zg����h�w@�CGW���[o��gtY��������>�uՕ��
�,.V �ԕ��.�Wv����+�k��K�n�@k�wפ�7�p��Ʌ��nw���Z�%��:[��A">qKa����y6�n��/��4���L�B���-��O�:��nݺU��Ō�g=&�ԋ^Q����dq�;��\�y _[Z� �Ơ�����'	j�f�>95�94ҩz��v�j$���yͥXe���s�t:Y�B_a+��2G²��A �1��mz�n�Z�m)�&�0J���L�E��m"���=#!
L��L�3��xӦM֞ovV(M��<y�Ur����LyR�%g .u������G�zqs[���3��!n<\#�0�ƍ74B�5ON�ld"�dG�I=a_��V��wL0	0p:��շ4�: zs˖M��U`= ��Y���o#��XvngP2�����׌.�9�p��Kv�ęH8ζ�W=L��c_q��<�,UU�,NM��U��׵kF��i�>"w�i��\m~�'�n�d������(k��}b���&�4�	(!$�N�&��:�C��ӆG�=��Ah��%���L��x-�I�hxn�O�	���t�E����#�����!k���!�~p*�U\k�
p��O"=�ș�,�y�j��d��E�L;�ʕ+`� �3.������:]��FL8��q��&@
�)x�4C�]�iB�UO����.�� �,"CM�:�G��}��H,���C�o�
�q�⣍��D�����
�=�q���#}Yȝ���6MC{���� �x��L��A�.G�p��h��K�lD6�(��P+
\ �E�w��W�@6�l�5�$��(5 밋x2���񏽪�Ry�Q�+�2�����_#��Yr|�zB0�kb��Ww���cE,^-	SP�~���ʢ6&�F�Ukxx�Q���N�'�=	O�S?|��x�����S��1Zk�kǌ&�
t[)�	������d%�${1�k~�JV�8}ď���g�ꝁz;�A����璗��z���i!CO~�)�v1x���Y�.�Ĕb7;�$i�$hb��nܸqǎBE'N��0�$=�B"+��o{�z��-�T#�c�@�^�7��aǏ��
I�ڵ� aM*A�-h,x
]X� Y!��5�dinOUl�� '�ڜF��l֖���ˍ&3�dw"s5N��8�6ϭ:\n��&�NG�*������p��׼��v�wh��Ҝ��"�f�������bi�_z�%Β~���-�8u���8Q��o7>E|�������.����A��$Kwll慣GO=z���fK�S�ιs�N,N����z�f���4
�b f��i��7�|��j���8Nz�Ѳ�$��xq�ý����.Rkb����@DU��kT���P��D�CK"@�>��=P�Z��@�g�*������n���ݎ�F����w_,R���˹���� [��[�G�f��c�Lq�㓸�ٺ %s�6ϋї��f���tUrR/wŰ�u8�4�q��lb�
��A��$M"�ǽ��/�H=�f����yL�X����3��$-܇hw@���Ę�#�bm)j��ʐ�Qѩ��F[����*N_/O�Th�R� �`�[��'�҅f�T�q���]K�£X��7�kx��G�ud٠�A��Q�,�����(M��X����:!��6��'{ @	��AȄ3��j��NKo7DB�7���@��es���M"0b+4,��Ɛ�I�n%�:�
�7���	K���-��f��ĶG�p�:�D]��	,PR���?�W�4��( �
%�f���#do�Fx�w\/�5N8��B��\(5ͅJR0z�9xҘۄ8�����̳h�B�%Oʂ�IՁ��)#O3�7y�mB�4P�D�	��!?u��zQ�^lNB(��z��������B������%����Ŋ�����ְ�&g@`�C�����@�홠�����䩰�Q$zG���ɓ �n$�!��2��c=N$�ׂ�;���/�j� ˵�	�8���	�ht/�Til����-�n��68�8o��ލDBv���CC�B*��n����,;=`�+���[cd���3��.B�Mפ�^�N������I#�;V��7H�ưl�Վ���}��'���j � ���,u^������z!S�8f�k�� �A'����p�Z�LK�~��e�Lwj����^����yy��ܜE��Vt��C��I\�2�.��a�a�'�;��cc�/_1�r�J��}��=B��ӧ%;|�0�D#��p��g!�f������2��-��=�q�VY�S��E*a�kf4N<�5o����^m���.Y��3���:�c�^�@ycLʆ�Lk������E�� A�ȑ#��2/隞��/��f�$��f`{�H��5�:$��ʼ�Sޓ���h58V���{Z���-̤���4T#Io�y�W�^��\�:�]&{�BL�D�V����(�l�,��iHm����9�w�\��7�I<;ls�Z!� /B�l��V����o�����8�Q$�μ7.�q ^��Bh��%�6B����i� A���]["斀N��DB�������X�\�$��`4[]%��\OWw�[^ry�����z��y��w�{Е]-ZV�����j��ڤ��8JE�E�$�zB�@v�:oEs�pe!��5�#�Sa�X�+nm]l�&SA���q x�Hy�!q'�ׁ��h@�#�� x�\�/e��P�]D	�uD	@%��9`PV�D:��Y�Mڬ�����0��hcD���*i:�8kײ�pi͸�N$�5��Ɍ����\�scЌw,��3��!y�ɉ��|(�n$�b��¡����ۉ�����xta�ZL��3Y�����V�E���3El.,�K��ۻW�6é��FV�FT+k�qa�H��JB#Q�v�`sƜ�5�۪��Gh����{�͋*ӗ��M����!g��[��j�{݀�:Z�i�kZ�X�()y�_cx>�8�Ӏh��*	D�4�Y�l<I|������Q$��s�,a�2l6��>M�ĕ�$�,yo`s�w���#�bu)3=�TΆ��hBϞ����aB��!D�o���48lB��0,y�8�o��ǈb�Drv׮]@�-[��:��Ν;�I.^�ژ:)=�C=��Ck!$���W�t._���S��u���@zG3��Әɂ��t�.�zr�n�m���V���z:]����5�a��tM]灾566v��1A���64iaR���E	����"DP-�d� ��4ƈ=����G����-_�����T��(�3��5k�N�I`���^L.�qV*�`��Hz�~��v�0�@s��+��ܹ�;v�>�"|���H�Ю�5�xZb�Ƈr��n�k�-{�П��SӐ�'@vaP�+�N�?TRd���K�'�q�m]*Uo��VB��:|�]��;D��VZ�w�޴�F*Q<Td?%g{�`(�'�A��6�8#��<�6�>��/}��_��>��׼����/��[�nmzr!����2	��ģ��-��6=��R��� ���~�հ�^�G67�F�F�w5W	��$%�	Պ�Ɨy�(;���p��s� :1�S�h '��T�9NjT�W��Vh}D=ȔՐ���.QsЙ��)8��s����1�E�+��� Sw���X����\{0:W�uj�7��G���V�ZcpL��t��u��Q�gږڴ�<ji�9�"� ��z"��h�
0�AqBw����FJ���Fk�|��r������$���C�� X�`�\�C�ŭ����F'�|����٥�G2�U)�>#
!,�
iOYH�g��p$.j��	*�(��J|�: �@�祁9,���6C��d!g���CÔ85��1���k��V}�=I�t�3���B
A>���C�����OCGK*�e)t���2F8e1+�'e�͎D�VG����&��Dh�ht��,�3YG9H���IS�p��U":�/��j-��=���~�]{�|a������??&Y+5�Y\�Һ�5�j:'�����]��L\_�|elolQ��馧3����[n2:����1\�C�n���Z[`�e3����D�!%\�?}�t���v%�)�W���xA%!Β��h�Ĝ,��{N����JR�?��?���B��^C�+������i%tA�38���c�2�*OF��%A�3������y�q2^��~���_��__z�%�}-��!F��$(�y�>����i��g�$�9}N�+��д;׮i/��n�l�h�����ܩS��9���A6�}���(r�uR��Y�`�ԍ��<]WӃ��┤�J㒚�1{"s��'��o�"���o��m���۶m���'�B/�?Y8�������v��~��K�9rX�Jh����[���^�r��e�O}��E]M�L�Ь��3g���-4�y�	��Ve�w�]w	y(��~������4��s	#	�h�4��m�j��ǿ�]'��k���,i�-Q�u����qvb�S��=�	��]�w�������wP'�����R0��_���n�d�kT
����ַj��Z6lX���,C��C�p���YB,��o����֭3@�sdd�����o���$�ڷ��-Mc�J9}�N7����ԧ����-,,��_�,iZ�s4Z�,m�r������46�A�]0��IxF igH|m�no6
�5n?][�;�ܤ�F�c	�C�>j��
3�9�|�N�H}N�#ţw��Ǧܥ8�P����S��5�L]3�)��$�Vߢ�-/GF�j���e�qFe�& �U�=�|���s�/^�|��7IyM_��gk��'�j��]*�BPd��? ��u�ȓ����%�I�<��!�����!���������M�6�W*�V�<\�_@kj9�%��!	��^��'��=3Jg,V�fͪVH��n��M-��ɿ9�"�1aPw���րc�*� eq��P`N�J>���ab�����:~)P��D��4�ݵ�axވ��tP��ݽ� ���Z] E��/`�۲��&�>������z�L�;�(z�(�D�j�r�ek5�2=�龊N,��LB5UA`�f�l#t�G���?�4�������j˩]��a���0	e���$�ٜ1��خg�W�K&��I�(��\�r��|1P�1��nqv���VӋ�I3˳Vc�1���.�����X����n��Q[݁/�F�=\y��UjG��/�7Jk��� �/�.+<C�H�Y)�s�I�*$�
�K.�<��O��9u��!e��v����%��1�┰zhy�@�����V&}mwk��&S^��Ò������#�<����>��'�S��/>��z����d�.��׾�����-�'��>o}��xQ3z�G�$����������HnoH)�YJ�Cx۔����/~�.���vۻ���[n١"�h9gM[N��;v Y�@d�}6��!����?�S���8��ݒ/H,F�D �7�mB[o޼�����CSGe���=R$�@}��N+v��Kꁣ������I
50Έas��:y����|}��5��A�S�����	g�����g>�9�V����<�Uk�4É}�[����J���3�y�Ʉ�4xͧ^k�+M�5r���G�*���g�M���ݦd�{𽺸��ۄ9}4BA4�n�^��u)ya?��F��w�$��Ha�G	�������}M�^�ӧZ������Q8'.8=!C�`��~�iC{����5f��@4ȵ5�A�m�3��G���p���Z�~�&M#�Ї>���~����2u��؇��ͅaTE�����������]�nYᜢT�j�H��n �*YэH��V��d��y-9��;:CC���3/�7(�%T�y�n(E,�0`_��1���!#ˊ('~hr��Q�2��^m ʼl�h�0A5�ALf��Wp�-9�#fx.�p�ʡ_�o$띪i�al�4lf�D����b5<b����b�d���O��Զ=Ȝs*�n��n���B�B�}�Z5�kצ�MLL�8r�8�-���Yx%��(��>bc�BN������!�Ρ�4���)���ܓ/蚥����!c|����t��"M���;6��%0��"DTѿE`'�N��v�yp+RE��fܷ� �b�299�C٩���	N1�����w�{�:� P-Ą0���q_ Y���#b�L��FD��j����9��[�Ip��j�W�E�c�}��0e�nrB�x��]k)��S��1�"�v�4ʁ�ǒM��vf�,=_�4�~AR���f	�K��\�?K:<vI�����g�S��ڷ��a:'ԩC1h
��|�yn8R�^fL4ގ�.�a���Ry8�׊V���l�����L��!��]k�F����-�Xu�l�T��9����H�T���e�"?A|��%�z��[�:~Y�G�I#�����o��I0��}�qf�G?�`�+_��{�������1��B��M/����	�)�w��G?��o~�СCT䂣��]�CF��;9|��+��=���%�����y󆅅��[��5���!%SS�}�S�z����~��lfy��6=��d#s08Vػw�}��jui��^�s�-�hqz�!�W�m�:1q�Z]��A�ann��0�y3�#<k��Z�����F�卺��R������vK�#�˻�� ���JJ����ԭ��Zs�	=�?�ik��~�'ڛ)�;��3z�cc\=\۲e�D�$�f��Dw�5�������c�r��$�T�w�p������	j0��}��;�\�v��AB�j �h-4�#Q+�1hJ	ءe�~;�9��tu���'��y�9��x�g��Dц�B�R�B6��x$W8�����Y�J3��C9[5���d�b)��E~[�DZz�v����?n��֭���)��/�v��f�T��g�$I��/O�?���%M낚�Xc�����x�� MP	x���l�j.���h�QP1��@?xC_��US"�UJ�QQ4"!-2���$UT��P%G��$M�7�r������/�{�Y�{���ѣ��\Dm�B�D.Eu9�Zӂ�m�6���R�R��$����%�/�%x+f�Xv����*�U���Q��������@��,m�>Uu��	l���EX���-xL[G�@�G&�B�>���T���Hr���~�> 8����!��D,��Q� ����,���W[c��-B����K��.4H��d���~�o).�]!�����wN7��2�i�8ƴ\�6p>��7�X�ﭐ����0�P1�\֑���s!�;	�Q�����7�Y�E� ���p��z�Q8�R�?>ÈS�s��d��aIX_������#c۳�c��i�4�t{�u}�z�ت�����5$�
�\����}�Xޑ&�B��p�W��:|c6����\�>_�۫����d�bn���E�%7��`���H��Et`|⊶/^.0�Q�y=i��8�-��Y�� ��A�x�E�~~ɲo�FV�J�R���h�ׯ_�ӫ�nذAp�駟��W�J��$���M����H�$�'�]{��Gu�7��dM��8&0�s�����nAXP���֜���� ��Wف�@�'�n��Yy������|�m��f���R	؄/-z'tU��]�ĉ����VQϒ�||��be橖ڜ7��f��vv�� ��#<��#z4�~�W~E_��w�������s	F.�t���׌��"�5E^}3�ZOꓤ�I��1f��An��\ %��Bccc�z5�={�"Fuw�=h`O=�ԇ?�a�Y"���~�� s	��bm'A-��#Gn��v�/|�/���V�zC�?��e�KM-A��[(�:^�g�5W�>��s���\kq���Q3P�q�����Z��.F$�.ugl!��	z�g���7�8����Mch#�T/hE#b�#�:���|D�y��^�u�Vr�)��� ����(<w��l��`��o���~�im�����4m�T���Τ�4���~�ONΐ]N{%��xtpf���_5^��� � ��t�I@'�SuӦM�&�,�,l*t0BE�	}�����#�G���-�������i�@v���'&���*�d_�b��i�βJF__�^Y�"�� ��$��F���^���1vc.Ԡ���w.�Y�������љ�];Q_�y�C�{��|�'�	vZژp2���50����U{@�Z�QR9ee�-�炵����ر�^�(p��a�ٗn+��m�g�=�uG���[F�X����O�L�ָxkN	Y�*Z"����իWa	p��D�* &�4$�G����l�T�@�VMB�4�!:����W�@��$TrΒ@���!���l�X�φ��z���i�4�Fvl<\YEE�e14�u�z1�X�g)\h�d�l�b�rI%�)��$!��-�ud��l��Ef�̇����X/,A!I&~�������4� �h����8 �z�uB���s�u>j�P����b����f+�-�'�B�M_��<#��\�ͥ�ǌ�JFBop^�9����Ņy�\Ê1�q�Ϝ<z�Dm#� ��$1���0�7l�a߾=VX�v�|ŀ�^��mГ�˿��P˾��R��I���#��Zv�9�|=���2v5�~����k�j0�"QQ���`N�:EZ=T5;/B�$8��#1��=a�z���3g>���	��ٟ��k_{��c�tk�ײ�Jyc�z��XZ�e/��|f�8�wAe��*kGa
hq7���.�]�=�������&��7#�������� ú��:nWw�D�Z���vҫ���\��r��aLHHw۴i��������WYI&�O&�6Ѵ�;w�K�w�ܗ��a]�w�RѬmڼY����y,>���H:D}*�ٳ/#q(�Q�Y��?��0M|�H�c�,֌�8E6��$�p�������{��C��Ǐ߼y3IQ֝ͥ!E�C܄�!u��[ږ�@$�GML�8�f���ai<����\s>dG_��B��~���������Dn��A����b�^I�e˄,x.��K��Z\�!+QR(R��pYr�~�╥�5��m�n����R�Gee�]�8��}�����3�E�����JM-I�ҏ$�k�t�81)8�lZ��C,����Dpe4�FJP�����>���v���a�%6q��Iu!ħ�K-.ZM����_}@S��GC|7�C�7$p�m�.'( ��ģ��%L�96��jc��H,�N��̙3�gӷr�����w�A�X��V�4: �;3V��,�f[/X)�֥dMU��i͂e	�sޔZ]�V���c�dy��S@�K����QԊ�t´s��3��5R���8J�(%+��P��]�}��#��r<��|(J�vuY��}q��i~)0�Ĕ�4P��:b�Y`?I��(�i�N�j��=@|�E��#J �VɅvf�F�@���,H�ӉE �^D�N�X|޴���U�Tk���,�\H�O:r�X���b| ���k�8����F�h%s�rY�S��6Vn<_gw�\��9NB��0]0[��Y��������>��ޞb��%*�0&[�vu�A+�<H�����%^�y�eQO�ϒKZ�}����`F��k���ښڦ7n�=�X�J!MNO'�f�R!~�|�ਇ.r�tt}�/�<9qM�����P����ɓ�������nz��w�eJJ�@���<��'>�O��O���Ka�����1@��7m��
�g���G?��7��;�C�(��IA�7x6<��׿^�ᓟ����E4%:%z�Z�	���yC�3
~���y��Yt��s�ќ�2B!}�G� ���ĉ4��\� �]o���.���P�F���9@s�3X��Ξ�J~�k^�����j=z�/7O���"�Y��;ê�k�?�Î/s;�*\{��i-�r���ͥ�Uܶm[�2�'�Y�%�fC��I6��ZJ�MX��O?��,Q�Yr'[����޽g�ܹstbe�	)�|�͉{(��/���>��:������K�r����*�����g>�]����{� 2�w�l�B�z�v`���롄�8 ��muE$K��F�� �LH1A%D=��~�b@?N�<�裏����֜�ؤ= ��sO����!�B�z���~�<ڱi��舼�q��(r�$���M�������!^8��HI�X�Z/f�(9�5�w
�CI�{���)��d!�Q1�4�'�_�x�u��Zh���ߘ�B�=�B�M4
(-�\�L�z?�IV�Y"8ެ�'��B@.��� 0s�I���8�����+��hY�|ň*{(:���ئΒ\¨�`P�T��'����ú��ϕ��Ŕ>��*x�*OA�v ��4 �wo�a�>��eXl~�������avcc멻�y�6ʒ��KM	QB2q�9�Jk�Q����v��Z�$EH'f	{����H::T�<�Љ(�$DBSO&J�nUr�0>4s�d���V�x���Y��-�{�wѕQT��_���9�Yw�q~#s"��N�2"�kvTD$�� i�E�æ�6��
N8t��L������_0)�������k�.#Gƛ�+�����k z����}���|H׻���I�%�q��HCqn�O�~���m4�����0)ܓ�[1��P.Q�S�g]�UH)4��0��&8�?J��E>7c���/6�ys�z���$��B ^-\Y�fՍ7�Xp�s��r�L����}�]��������LO�ZJ)�Z�#�Pl2H���n8�T�_a�O�gz���;v�8v����*����~���K_�]����iE�̰��ŋS�l>x�������%�t5I�7��[�lْ���W(��s�\hמx��>�������^o�y��� ʥ�$�t���������*u"8.�,�`�U��}h�Də3�EV�2RY
� M�������x}�(���g+p��eU��sA��2K%og��K����7�
�ge������s�z�%��5qf�Bz�_�I"�`� ������ײ�����={��"�Miu���;1>��{�@E�	��%/}՛�qa|��_�� �<��pH��U¯��c��C#��.QQ�(������6e�-�p��:�!��+���P�s!|����M]���ba΄GM����b�6�+0���৬�����7�y�֭z
� +�׍��uMj>��Ęt_:>���a�Q��{�n�[��P%ʷ�3(`�Vu'1!�G�
E���gSv�;d�@TA�FRh5ތ)ᐫ��b��3\�1����}$��#|�p�l->�n�б�P��y1r�I͕�r4�EZ�ݻ؄hu�-�'�&$G����m��cm���t�b��nv�̤D���;�Y����]�јx��,�qR_��$�[��PN�` �4�� D��`L���/L�f�3)>c�����k�B��1,��$��fҸ�KdDE��R�00��gH1Ah&�R]Y>0{�_���6�Mx�[m����w�Y^���t�X$"�:c"�y�Ύj��|&*�,��Q���~��%N5B��y`i�G�Ta��z�_�5� ����o���R.4��+G̐��/���sZhw}51U��N�.�'��P'�5�I���&�7)m�`�].�wܤJOW��~�!�ވ��0�Y�� �����$�h�����mFԂ\��ӑ�%L�|��I��$ڦ͛a-��)�Ug���a�$~Ot /�.�ҥ����hG��x���+v��eت���OKN�!�#������,�]�~�c{��'���u#?��$��l��j�^��Y0#`,ˤ�u�)`]DX��3�W�>��SB5�+1��)������ʠQa= A��铲��+1�Vh9�W$������ʕKҝx˫�%ݶ����G�d
G7�~�B7eD)4-��}��Hz��o���|�#��X�I0s�j�n�4&�s�M7YϾ�rbj�צ�d2�;o�eW�NhY�ctۣGG�X���x��i�&�=�R��
<�o\?11�'�'����!}8	���$*Mj>s��������{����am��	A����~��_�ʊ�+�Hɩ�f��5	�v�ڳgR��F�̕��W�<t��3�<�ַ�E�
��9��6[��J�?�ˤ<��	^��ѳ[���N�h�- ������׺KdP���R�4p�C4ж��������0�[�tg�yx�+L+������Q:T+�c��V�=����6|��g�|˖��s�"�����&�z�ka&�/1��������<�o\�+W�^���l��X��)�v�ܩ��nѪ�lj߾}M�,�:�)��,�@�}��8�Q�:����!���	��4��74�狱J��d]-��%��@�4$�q��-���a쁥�F�$�#�:�%�P�6�P��Drvo��8#���׮[ժ�)��^��^��{�b7�'����%�1v��)O����
�|3��B^�^����^
�׶Bu?2w�K��2����IT5�S�ҴK&��7nӳ�>}���6m����ax��X�;צ5R퓨\5��!�0</οVh��u�@������ϔ*�B�ۅK����(ɛLBnbT�D�8b&J��L;w���O�q6۞n� �+c��˨8hF�=k�%�P�`�h��Q�X����		�4ë���.����4omZV�zcd�V:����^��Pz�Ɂ5e�0�b�,����Ľ�nZ���PZ�3���9,Tt�eI3�@������Y���f���[��ry�����,VMdԛ���R�K��������l����������������̷ݲ�I�穕�/��.,hv�[W�^�=���._�w��W�.j�]]�S�N�H�9wt��X���R�&���n`rzvan��k��V�3��gғ��b���K��ʹ.����/?��c���o�����ӊKuj�s�3��CC��x�;��Z�
����y/�{*nl5]v�Φ��s�~�����w����o6:u�N�v���ɓ�4����G�$����H�����_4A���7��~��9����ݪ:�����
B�׌fL/�5����.<pD������^ڥY]F�￼F"�s��jt�ܿ��v�]w	Xhj��,騛��%� ��Hr^S�`mY)�:j��ARw�̟;w�_��»�ф����>|���+jh���Л����J��~5o�r��eb���SP@��_��_���{�\]ٮ����g>_��j��*��зh�==�];z��%��;.�Hx⩧��r'!�"�8<2BM�x����_��<������қ����q�F#S��a�k�&�-�~"kX����HR�P��@I��"�Ƅ�Q���з������r���I������׾V�I(��ג��4��^���7����[q@����	�W�Y��q�ĉ]��h�\)z�ִu^���_5D�z�����\���c���'\�k�ܼ�y������/�$K-=�v�Vm�ڌ�����&\c[Z�L&rD`&��,u|]��"�>l#�t͹�6L{��%�?����׽�A��'��A�WiQt�n��͘&
��N.�������y-_3�dU�����qm|�
N�-���z�B]]�row����h��zcՊe��d� �zIx��bŲV�)���ۗKҹ+E\�ˣ�#��ս���5�/�-�K�׬]i��nޒ�YҐ���KZ��̴��Z�ohļ��%��J}��t�@��u9�2u4?���z�V�J�Q?�Sj��335��Ҟ��}{^�LA���?zBϮ�37k�}z�����n�7S��������tZ�Ds�J�ث�t�Y���H�Ѻx�֖z{�%�t�Je�X�~��lb��z����Z���Q��jŵ(dR�֦/����Κ�/�l����_�F.��VƯ^[�f������	�ށ��+��=ܟ����R_[qL,���zz����i}��>Y���<ߎ  U��V�9�!��[�F���_[2F~iI�rY�ɔS���D����r�e������֬�%>�X�m�a�c��Ӗ�9(�.cCK�p$=Zk���A0���X5'�A�.f�[�G�n��XʅJ�z�-�ىG7��,�c�R��݈��d	��44W����!Q�\���{�,bk�{����
c��`�f �͇j�,�s�ng����xՐ����=�i�̛�R@J�@i͎���Z�hٗ��=�Չq�Y��I�\�����&!���(��^�Ibkb��:����@�O*n��QR��[G�n�YA+����\����}u)���e˵H��$�%7�y&�v���֬ş����FY9ծ��:���D?gI]�.2��H�R�| ��Ќ�HK]��o��>@:?O�3?�3_���?���Ռ$�2��"������K��%��14C�!4�>����_��w��4�z4��O<!��G�G���g�4��`�h)b��͢7��#�V��7
@�.3gI�6T=���b�
x����w�����������Xw?��k��Q�$����Wu'�5Yw�K/�D���^j��.l9Y��E�x�A��B�"���E6��!gxd��kW�h�D�=��w�.r�c��G~��i�>6��i`���8�t��n�i||��}4Z��������>��~SL�� f������?�A�3���������#Gy����#Ew���]�!]������D>x�`��c��E�`��-�u�p'��������x
�.¨ʅ���'��.@���ګV-�ti��/|��tЅNu1� ʣ%�"
�oڴI������/X����~z�k�f��޽{`������O�<��טWt�B�Z���̺��^xᅉ�)�>|��C�A{��Z �9�~���A��i�C8Fg�4]Ք�֘p��Z?:�
,�<ZN��I�C�B�X��י�,_F�^�9fY5�4!c�g-Va$AP�'�������1X���X�ի��U�\CB�ѽ�Ȇ!���Y��@b>JKs�p�d�����	��M��4�	J�Hx�zC!q|(���Ax��<w�B̃ly��-z5��<�j�Gޑ����6��N3�!xK��$A��b�x�����O:\c�7�;HG�uP _�E�Z�`��a,y����qF�`-�FCMW���/|�h�)��&A��B�S׆y\J��@��q?]���o�MM����IA��u'3Z�j�����Ya�����{z۞u��*�A���2Ϧ��\��x�Zitt���"%2Y���g@x����ӳ:�ڨ RG�]e���Ξ�H)�+W��J����lΰ�j.���%wi���B�^1d5BkR'��c���N�g�К)�$��r�[�_�{f��D�j3���R+T$D�U.���{��Y@�������dA��`k4�e��������Nb��~���t�C�>���lެ���� �vFչ@uh�� �H��%�Y0��ssY@Z���BS��>\	��k�WJFB��O�"|�����IF�
)�dcD5ëVvk�~�Hk��ŉ�<���o��o*i���c\h@z]R擟����1��5p	��Ƕm��zj�m=�w��W^y��cUHUA鋿����k��k�x!]��������������=-���U��O��lH;�ЁD���KP�.��_xn�jn�9+k�jI=��ۻI��n
� lv�C��}�C��Ǟ���[!k�M`6��/��G�������:G����g���\-:�zG�,���5�"�zg(���Qю�_��Jr�s���}�S���9<lK.8i!��v����ǵ�$d�
��'8���g~�����ׄf|�;zT�{������T�c��2�|���>W�`�D��a_��`�5�;vh���'�K�yuA0�%�֭ł�^A�ܹs�����F.�M%�?����S`?��o4��s�Ia��_~�{��^̼���Eڮ���Ù��ݔ�]i(ߦ/�sg��� ڙ������#���1x,c�,l�=l!��n��8�l�� �D,F��][;���9PEgp�fÛ�̓M��ApG�B�T-��M���d��zN�jX(P7�G5�wiԖ�G A���.V�L�>���lfd��IǪh��ٳ�^��~��)���h∅�����U�sse`Zy��Q�=&�<]`t���k����ri��@ 7I���4�vYc���l�K�#��a�z�z+����$��>tTs88ػlt�A���r��>#Lf	�inh`���&V�^)���;z��M�i�P��I~/��(q秡��p���/�Ԝ�,�"��u�t'ƍtF벮�n�2듦'"���9��j��/��v�6(�w��3�j����D�6ή2�1X��'��*l�4�c�4��Q��:m�B�@%
�����w��H�b�`T,�O���t���`t��[��\�t��RY��Y�Z�Q�5��3R�%�P 3�-�W�6!���R��jn�&'%	��p�-���<$�]k���"Fo#^�:�!�PЉ��=Lr1�������,��eyf�~�x���,pDI���3�\ɫ"D�yW��K�J�]q�z�.(Â�?�ܺ��߳8+1�X�O��\oX^�F�V��[�©�#Dމ.N�����!<����.gȼ��{oo7͌׮]�������~�z��o�.����������M<H�n������;����W5�ee�_y���<�ɓ'7n�g�>s����}�k�_y%N)��-����~��9u�4-P8*[�l�����~���$mMg������#8~��氯w ��Gؿ?
����y!���-�ؽ{w����6�nݺu�|�;�⥗^Z͕���2)��27�)�[o���9sZ)Y��9zF��� �P�F����D[j�zL،0��4���k����N�J&��,�G.�x=���0�7C�R[tMR���/ٙw�y�97��$���������4���o���?_
���T��ȵ3�S��hY\�+QZ]������p@��iӍ��sg�v���(χԹ���>\��������}�����e#��n)p�♐t�}��ӭ��ӆ��G��?��w�Z�Dt)����}��Do�!#����nﳉW�l�gIBm�t�.0�H!%$M<[�=L������W�:-W����-�o��d\�'Vh0Ϋ��b�4v�'�'��I+#/G_єjThw+o�X}Xj[sB�7/�1��1�4�˄56 ��5��hg$	Fz��2*cc릦��y
�C>����c�U�F�]�M��?���\Tg���1rB����&Y�Jb4C�u����N�ǜ�n8���b�k�t��]D�M'��i[)	Yы�B.���(w�>�<B=�����Y��fEjl��[�W���"��* �Je[���G���&	���.x�.�,Tq�j���~��B��6G�';P�LAtꔥ��Z�bq�����7�e�LiV��ɽCv��ۙ����$h�`�v��~I���IЃ�3��� ו+�'�p��r����5LUT$��a�m�8�/���`�,��H���F��]M9�g�\�{�0e.�h�!��#Q��#��0(#)��M���l�
o|�5N�j�z�a-�d �Ia��T��dӛ7�t�]�n	��j;�����m�OQX(�4�bf��m��n�m�D�3=�+`�1:Ĺ@�˚ioZkX���n6��{���C��(�/�Y����,��+\�dDV���Wh,��'Ig}]�EKHW�v�[���8���e\YpJ��^z���O�.^���y���FLv�{�������w����(y-c���äp���z|�>|R�8p��q-ۼCFz�Ps.)����o��Z�D�.��3s_@G�=r�0J���N�>�U?8W��w����Z��Z=u�u�zv��kt9�TK�k��H�o��z�;�_I�^�f	����#����xB�;w�QI�����"�1�����	Y��]�v���R7F�^O�6�S'�h6�P��{����S��^~�e����η��m{��-x]X.4��V��=%�7�O�/7����OhD�y���o��>����>��m���,����{�s��O?�������v��<��SLl.$�F�k�a������6�f���g�E?���S�6�@���N.\�M~�J�ӨschŅ��FkҼ�֭_��͞3��s�\�:.#X;gb|�����lٴ�};\���*���c3kؒ�ڃ��?_ַ$R8�˴���:J�����sz�<-"u�9�	�THc�6U���z�P!G3�Z��4���L5O��_Q��@ �I1i�s�׽4��¨ȧ����о��0�r=e�s�Y�kºGhþ8_�p�<�:����:��1�	��&ןt�uw�*��Vݚ$I<�pmݨ���6�Č��2FzzJ�F)V c�)����D�0��hb�Po�F:Q�ۂ1�Q'�k���PY�V�����0׽#���H�s}���R��B�'�EG�G6n�0�x�Z�m�y�ױ������>h�Tزe���,����Kʜ׆�)�E�����`fC��6��%�G�R�F:#��E��8)(�b�d!��G&��$ݍ!��2!z�����u���=�\���a$g��ek<�dF//�ws��>����R���-�սX����������V]����R�K�4�rk6�a�������vmu��F��b�S*ՎY ��N,6����Bw��%b
�+z�yd� �gi���l=�#�<:�tDB#ڋq��8iȱ�"�Д=B��M�T���"�Y/��@�1��y�4�8������B��u<�gƴ�'��3���f�g���'����(ķߦ>�C�e�VD��c�yC�vI�9���"�ޚw)��Ǒ �� ys�(��GF��z�!MR��� �~��������s�=��]G3=}��#���C}�+_Yrw�Kj��=���e��}K'�h��� }y= �Y�ԯy�k~�~AB�!��9��}�+��5�h���^��+B�R�����j�v��r�G�+���*D�g����w��7����p����K 2�J�����pN�A��#<1k�6ha]aq%�H�G��.`k���k˖�(�ś�z70-���t��F��Q�}�v��ᇿ���F�n��7�d��0�$hv�ޭv���k!S@��c����� p��O<�,@�`S������y��B��ׂ-�&&��cI���L��W�u!� ��K����Xs�)b�n��رCD�|��5�`��˖-[6o�|�r�1���/h��S�8m�cq@w�j��}x�ΚHeC_�pՅ���ڨO<��s�=�)s� Iw�ݟz�{�onԩ����� ��Mh��f���5J�y<\͞,!-~��ɋ��oǤ��x4�
@ΰ��X)�z��AȀTt|Z��FEt0,�;b�Q"����*M ��u�X<��M�\�_	���F�^]l�LƓ�#���N��`����;VozbI�9�)T�#�(�@� ƻ��GL���A�ELsZ7lX77�sq["�1��\�Ǆ�@�Qث���A�5��ڈo��;3SY�j٬S^��s `��GZ	�N��H+	F �B���o����W�ƯN9,���ͦ�s��aH_��n��/_&�b:xi��3�,l?��I�M����4����W�U��X����&:)�!��^m9|R�+V����9
���\梸���h�9�?�6i�:bbe-Uk��OήML��8�>s�,�s<�z}�}��s�]:.ss�h���{�F�E��u0�-\���y>"��u���p:55�6����qJ��'�Pq\%��8 ���1i�@�@����_*rM��|G��6�*����?�!���M�Z.P�����\mѢy��i�c��SsiB�� +sHn	��x�f�7ŭ�A�Z4�%+�9c�p/�Ay�+�7��,Vk��2��fK�������	�k�^�|E")u�NiHe`���FA��zmb�V-���/[�WI"�N�����&iR$IW�_%�,�sv���vs�%��x���5��z�y��E;X��t�?����T2���۷O����$�����7���Rݔ��G�x��֮]G��^�/^�I`����fV��6��U�v�ۊ�2X�m�&�J���x�ᇧ&'+.���sy��7ܰ�رc���hww[v�؅�^H~��������'}��*uKl�@���r�CwIt������u�����Ns"э��l�,�w6,/�i�T�����eO����cZ�����)�=�7���������M<� � ����a	Պ�+Ã���h��p [��k���^W��}�����7iY5`-+�^ T
5�=����B:u���7��,�}}�9��ENR��i�ða�B�w�CK����Q���~�gV���Y2x߾�ڟRu�o�y� �ǹ����0�b�����f`lCٓ�e����G����,��;���f�y�u�͓ q�1d!��%W��6��6Yb���,8��p�ސ�]Q9����,Ff���B�c"���
�1�h4]����J�+��%9��'�ŅEҒpab��,��ig�?I�-�m�R�~z�p���i�4�vp<�������@*����d�3��
�rZQ�'EN������4 <"�u��xbr�{^g���'��=�u�
���i>笁CZ�B�(��j��j��@�/�3�:z�i�r���W�"���]�T_2����W�nۆ�0�4�Y,NM���cvz;jk�����d"Z�`�M��������7MNΚ��'������9p�a�|��f[�X7&���n\�f%f	|��$�*����U�NM�JW&�*�Ar�B���R<�x8 �p#'өfX������hzS
L,*�	ģ�1�j�7R��P++�.������+#MH�P6cB"\�X���_��s��7������s�֠�����V�}N�$Ի��1)��fg+ў�<F'	:c����$0���G�]��E�Qt���v0�$�fȨ.��}{�����;	}���+����Nw��YG���mX���b�:>T������3z������}!�m�0>��z㐺�=�,EWkL�5&�������16�,oi)$#���ʠ2׬^K�!�v�`���.88�?ޝi2M3u=h���"S�� �&�D�<��S��Qov��p���i~�׭[�[`�2/�Jo�6Ӟffp���i�q�&��K�J믺�>���|�^��\A7P̂���cP��uN���f����龻w��2��%*0Z�E�c�ƍ�̵��������+�������ַjN��v��ɀ��:��kH�������)�ܺu�����d�5�����i(#��� �ć�4��
0Wye�"uĽS\�ȑ#~��&jj�ٶ�5=�K�h����ԝwZ�U#��>@���	�li�\�5�fmZ_����v�{�o~�k"	���E���ܺ�K/�$ ��O�s�=���D,��"�	(�x+@�V·"�r��Q}^�D�T���	�i��xH�ծ�}�ނ��TB��J]�T�A;���N�����-�
ڴ��;vܢ���ԣ<
�ϼ&Y��2�;PO����;�q�v���~�Bi�Y���"������V�JH`�|Ŏl��HX���$��!�1�a�__�#��� �
��{Yf�N�Jȑ�H4մd���4�x�4ϱ�E�������k�d��Ҷ-�%�<�IҠ�괫"��1��dHm
o��p��̶m7MLL�w2��3aFJ|�p����Cm��3�'��ζ���BA��	�}0R�N7�vҧ+	I�`�c��K5UL �ן}�Y�M�v.v\������{��U���k�v����I�@H	-��Ҥ�f,8^�%�2��9�k.�ol|��JQAE�"M!��H'@zrROo������f'��/���g����繟v?NEi�挽� k���]�m�n=�������t+�܎�Xk���v���
z@��N���]!3�C{�	�qH�>�|����@H�E�h�%�$s�-/^�H��[�l��V"Tb�=BƱ�i�:�W]u�������;w}+*V�5¤�'�N��,��U%?�裉�5~r���imi�s�!J�%R˶t+9�eh��Ӑt�5��b�ֳf'}ꩧ���@�W�̭2Hndh��}�k�~�I�Ms�|��.��Ƒ���B�a�;�_"N\��k�9�3"�h�E^w�zWPK1��Ș�P.q�$�gݙ3�;7gl��ՊO�"���!�LsL�^�3Kć�6JF�u�ʲ�� �|\��Z[[��h���4�w��5O�+�_�qvF|�(VKe.��M�+�{K1tg!��C"�
ѧ�QCl:N�l�f�Y߯/�9��&P��M!u�C=��	�_����u�o�Z��ILӰ��O<�rG��a�a��B �h���Bީ�(5q�#{ԑ>v�q��+����g�z:���왳4�ڬ�<�7�i��m�+��H.T��S� �������/ﰰ��/͗�n�R$�E�L�3i�n��_tS	���Fa�V4�����I��:���qI�H,��׿�ee@g�����+�p�%�\uՕ�F��>��1_����eּ�j4{Hd�y�g�(-�`۷o[��Y8Ne�T���d����A)Z����1�����.�s����zFiL�*�4ig���8�6u�:R_ ��:ytL���a�f��f��o;n�+��z(-�7��M���W���T�9�'g�u�ʕ+#KM@�b�ډ�;:ƌ��r�	��F"�4y�$[����۷H�  �Vl)�d�Bͳ�����w4��NQ!r5�|]���4��8�A��M��Y'E�#�@�>�hu�����X�� ������:��;�,kr����3��oN뾹s�	T�L��
�5�|d�@��lQ�+�[��AK���LmT��2����#�Z��{��!��Z|�ӟ���8;�Å�W�gәb��*�+�=�v���j4zT[KS�Ӹ�H����t)}�u ��6,]�>nٱ�yd۔�\�٫��D0gI�n��B��t}��Rs�Yo,�i+���t�<G�t&K*zdu�:��["�Y�O��#]��T`�֚�X��{� �Ǧ�oH��g�T~���6���h��@�>'=����B�@��� A^��M)�F��j�ƍ�\�$`��t�[n�v���I�^�h��Y���,��|��wJ�tp�g�F��p������N�.,^���?0 +������Nx��k�(U����s*�w�U�^�,�cFj?��X����P���+����U�
!C��KV޻���+�Mƅf�擈^��2ǋ�`V���
���u�HgdB5���	�kxa�j�P�������o�q����K@j�����/�Xzl���X"nQ�B]%fK���uTm�X�������^�LΙ}�;��k�y��C#��;d���z{m۲u�NI����W\qEGG�XJW�E�fL��=�T�g�U���H��SH��؁1#_x΂�s<Ӟ��;j��#K�6]�@T��5�5��%�s����aO $����I���}v���,Uh��z�h�H�G![h��R�
y6  ���������v�=~R�D�JV�PNxu%#�nߋ�$c-r5��~���)�Iښ&��C����D�3�*�㪹Ʌo�'�u|�`�Q6['�@<(4�љ�(!?4e�� Gs���'(��\ ���vX�4�d���&C)�=�ܣ�?�O��M�慖�����SN9EO���Kkozb��������$\�!I�
`m���N^ʷ��X�D��k_���t�g�:��D���%{W���w�Ko�}��d�	��|��Қ�wB��O(�������'kX��tw�74,Y�D�o�v�F�_�J�W����a|�<s��Ri6F��e�@�9їO:�$=��6�Oj�(G�,�O��G0����I���k:�Nь��F�bh�Ǝ��]4Hh����u>���ix�V�Bo��K%(׵Rد�/�A�>H]�����;Q��.p��
���g�Z[�u�i�z����&׊*K!W=^(mB��fX���_�����K1�yѵ�����,1�0��6�cC
�ҥ1d���L�QP��z]���!���G�Ep�Xv9�:����#�Ɛ��p�u��M��jrd��EY=���s���N��|�J������a��P�3eǎN�����D��U�m��7�vBH��!�5o���{ H������RN7��+֑դ�`�F�Ϊ����@:U �BR<�z�oԟ�6�f�jBN28"��P���v����:/~����,�lUo�<�^	���T��2�C`���]a �<�y��*[dk���L�O(����������m��&+NZӦM��n�tG3^��N����yA
x+K��.B]ǘ�Uߥ��ZG.��YŮ���5B?qM�S��}�fL��V3u��p��#�H#S�1GV-tFB<J�&A3_�TL/�;��n�����0�i�J��^�[��a�����1a�	�6�o��s�9����@'0���\y揑��w�+��u�]k֬��c���=��|����$)�\��nx��ާ�������n��v��3���7�!���/|A��Z����W
�9���̜�?� �S���!`W��!ȩ�j^����-� my�����`�k�.aI>Cɷve�|�u�j:�W}-B�f�kr�U�9>R�4����_�Ύ`�l��]Q�	%���4�fp=��}��DM�e�Y�����`κ1�����LV�;^�H�Ϲ�d	Y6+�9�V*W�]Z�+��;Z���폪1�����r�2d�/������˷N�DRO�n��pe�c)�|��G�lvA.��m[�n����ҙ���F@����{�WuѢE���GGRQ,�#)��C�q��XkCv��2�G�Ԧ��u��&CO���7h��+V���p��lL������7o�̙35 	8�}T�pM��;n�q�;��,~�wo�ԩSJ�®];^xa��q�$Y�c�U��L]:�Z 	}A[]G�L��Ԗ-[4{���͛��3!w��!���K�H�j��5=��� ��� i�zqJ����م�Hr��L#s%�D�Ћ.¨�ܠ��}��va�2������}�{�����酧]O��)�"K�&��/x�]�v��u�D�*رe����0[�QK�U����!^�t8Ęv�ڥ��fP�)Ezӄ��0�A@c��2i��	D�%����Ղ������А�5�ppJqf�o3ѥ��x�]�(�˦���1�k6\���y�N�0a"u��#VM2��EӸ�ŕk׬F�w�Q�Z$ʴن���D2M���_�hl�>D^����Ac<N__� �����M��v-1Z[i��Fl�$d�>����)4�x˨�=�����!�	 N0��-4>:�;��w����ty�f���D��ґ�%�A���E�o2�ڸ�t��W ^��.!�����5 �$�e���
���f�(��"�^\�^�BACم�g9H�c��c��U�z뭷~�_�0~B��nim���f҉��+I���d�}C*cv����B��F��,�{odP &�|�98���Ј�!��~> ��	�iR��tУ�?>��Q�w$Jf�4z�[�m��%����������
ƉOXcpp8��#�r�Wm�⥡A����6���� ��f�NwŴ8 �p_N���n٨�!��ʓ�3�m�nWJU�x&P %hjr�<�̊+�{v��5k����뮻NW�3g���s+WH�koK�s��g?��olnmy��y�b8z�O�_u�S���#8�@lO�W�}��f�}$4��R5�]�sjp�����H�H��Q�'�z.�,�n�x�8J��0�..�db�?W��y�1���w�̨T�޹Lw5ak	�`9i!Ԣ'"a�GA�`b�������b��5A��X�Lid�}z�N�<�����}���1;�k�'�e��Ld���/I=iҔ��'�q��q.�c�l߾S�q����4Zv���d?���gϞ�茬�E��CI��ب�6=�w���w��]����&L�x��g)��'m�1@+;�|d|��Τn�����8A:���q����E�#_�Ε��.�@O!��ց�c����d���BK_#��%&���5��������.���%��?�At�+�sa__�8u���w�X
��u�|�R� ]�4Ϻ��-n���?Æ�G�ԳK�z�Z��^��	g�����u��}ibMT�Z���#�A��%���k�tAHY݆6�]w�+�CN.��&m�������h4x���B�yc��l�y�(q��[�c�j
����BT-�v��jժ������~.�(�v?a�D�	���? �+j��+tM�`������ L2ֆH��ӟ��ۓ��N����s��Kb�T9d��F��܆'��_�1ZU��^Z�����o��Ma�j���~������rY8䨧�;��{s�vuҤ�}'��˖-�H4�$�N��;�V�Y?yQ��m9�9})4b�@T��0Hn�x��ѵ�#2�#6=ͤ<�����R�����0"v���,�L����
����'w,'Hǂ�x\?'������'j!_�!�V���)�C���l=?P!��"��rNp^daYș)?��54!�@#�1c(�;��{��65F-%��J�pp�+S�0tz��< �Ω���72�;����(��ea�F>���~@��m�8S��\��]������p�7����c�0ׯ��o~s���[s�n,YԚa8��jC#�Q�$���
�YW����e�+�	&�H���N󥵱�Di���1,^���K/�4u��X\KM+
֦u(0imU�@����C��q���ԧH���׿�u�v��M�0$�/��2=��E��|��R��$L��_��W�Ȯ���Sf���&oA-���S
Oap*��]��g2co����A˾�)���Iv�V\P����y�T�	����]��Ȧ��}�!E��y�q���5�XTܺ�JRn��fM	��}�:��k��>c���?0�Ҭ�E�s�r�-�B��(��>�6�Gc����ȫ7�Rƪ#@���6�bssk�
�a�Z���IS5w�!�D�T �/X�w�D�K
)R/�U]D�.粃ꛄ6�Y�ܦ�������T�'����w�}���_]I_�#����h�ܹ�GW���$8��%HN�K՞�Cc��i��+W��Lx���jD4�Ve�͞}���^���b�j����/k�Z�ɓ'-_��D	�(Rގ+���	��/̘1͹"��Y��ƕ:+��Ӏ�_�h�x1���&���]�r�����o~���"���̃}�)��:B۱�K�:S�E�D��h�)����տ�W��`[�Ns���u�&)M��ٴiӧ?�i}M[���#�����׿.t����dwf���C��/�Wt/ЇZt��#q(_�d��O��F�Ѧ��`�=���VG���>��m�2�	c˖�*�"`-����q���v��&U?�+�PT�9�h�]A
Qڬ[��K���m6����w\3+�<����(�5`}gΜ٫V������R��ii��g ��h�tkks���hA)flmuԆz
���Ɔ��āG��~x��'��=�����"m�A�|h�:��<4��cˠ�X����wD�2{h ��z&�r�V�N|�����݄����]q5ֈ�C�-�"@r�S�crf��2s��n��w�I:A�Y�f@֨����(ĕ	[�� .�̶:���C� 2���-�x�@��*?"��Xa��9Avb؇y�A�L�*B���)�����˗��ߦ�k�;n
�1�.^,8�]�4S4J��dG�5�S�J�0���z��߼J�t[T�X�k@�f%��G���+�1賴繭�_AO�>3'(��O�
*��X��-���^��G�=�$����M;������ߖfH8�B�H���Ґ����$I���}O�����v��j��d�Β8�y&��N5c�H&m�����V��b��}�:2��1d�:߿��՞w���;��ܥC�o}k򴩃#Û^�����;���4	ZY)�����SO���e;	�-]�To���/}�#��}o���+��������O������:A���1K��}�LM���L�&` �V���̆���(�[K�k��QMp��	hp����{��0�����ʘ+�ٟgllt����!�n\��T��Y���A��n�Q��xr7���d�G��Āq�V�dF�0�t��аc[)���&����3flپ��p0,]ۜO�rE��1e��x�[��AO!"�'�tR��{�-�O�'���k��#�v��Q�q��%!q��ȈruI�:}_ot*��u����?�����i+'!�L�	���O~��ӟ����gԡ,)�ohpi(�֭����_bj�O�P%�H
iht�_g7��]&[�Mq�����/�t�����S&9��	&��ZߧO��ч�;4H͉)�,�m۶������K}�h�r ��mTH�k��~�y�Gt,%��La�F��7&<k1�N8A�r���y�t��ε1֔� �(&SZ��H����~�4n۶����6tq]���ჶ�Q��v�1c�b94_*��p�?��?P�Ox�Y��ĕR�B�����ʘ��+�l��	���S�6m�r�y�i҄�5<G��F(h�-�q�F���09`2ôdS	�hrH�������F�d��"����FBD�ֱ�u�K.���R��1��$�0p;��g#D�D -�(V,d[]�^}}�$n�����e�c�G?�� �n���;��d2�f��CQb�n��?�d8��� ju/��rP*L�oq�G#8�$0�T
�2fa�ρ`t5G�`kA��=I�ćU+�&E{�X<g���W��H��ݤA�\n�&;�ل&� ���	�E�'G��'����|@梦�|��s�QƎ#-xj�C�*���>#�k!�[��<�ی��J5��<����I���=�Q�~��t��a!��̰�R�@)�����ña�U�6��BET�.��y�����R���dWk�b�/|{�n�J"GȮ|�S��u�׊���M��o|㦛nBh-OH�c �0nf��/j����
��ӘR�����h��G�P�3�>`��^~�eC~m==}xv)�v%��.�TV��w����W_-��ʥ��@ۼ��p�J��6�Ǿ���կ~������?x�UW�p�v�=��_|!����� q|�/�<9V,Y�c��'P!�c�w#�Ü�$��&$x�D=a���,zfZ�e�顡���j:��<l��0���zK2DJ_�����aR,O9�ɨ��-�5̣���GG��|l�t�V�ŲK�:x��PWK�h��\���PǬ����(/r~�Hj��僻d2[��pK�������^�u����V�n�;J=�i�:�WG���zH�	���mpS=�.�7H&#�q�������}37-�P �z�9ЙF�`"�[�(�B�UK�_Iuiؠ�5���v	�e��3gΤ	��J���7��j��+��%ܯ��zj����nJ_[��4�Ri�UBE���k���0�q}�Qr���Q5
Z����P�r�)�g�o��{�'�������AFD�a�Ė�,`�aТ�HB7ԸO���� �f�����.�,\�� ��֐�Ӳk�#�p�]wI��I���]y��ɟ����O=����23|l���!�?AC ���o��|ٲe+W�c�h��T�4;l᪋/��@T42�"�.�e�����4.ZԦ�����)�Ν�E��b��ݥ���њBZ�=����:ڿ��]�>܈��%tyDDX�/J����;;j$���O '�6��f%� �S�����_�_�v�y�,�&�RO�[�Y�`�Em~=���E�w�+����+W�_c@
<�N�e3ĎD9�+y�9��bK�F��!T�-.XЌ$%�)� 5���(�{�.��󎤒4 ������Ό1�P'�s�{ۅ��菾 �
���q��	X������:@�F��pL\ZL<��QJ���GE� �^�Q�1��ɬ��S�L&�������k�R:�@s�*4�/�8U9�`=��e'I*ew(�)��su(?Rq}m��4�S0^U��&훂�}��_�M��d�Ȁ��A5�P�1u�W��ER�)9���/ٓ�/���M�?�����뮙=s��B*�#���s��F�8�$\{��7����O2�jD2II ��QYF�#������������ p��+[�&j�x~}�W������}�C�uj�V�[:PI�~�Cן{�/��� ��������׍.���n��Ļ��.x��ʐ#4LuH�|BH��?zŗF�֠%C�#Mz<Z&�ϫ����}ޙ���S�\k�YTkx�⚔�J�\[�O�S�9����>&�����\F#P���-(�Շ=��ȇK��5o��B�b�&�ւ373��U'S�qP]L4�Y�y�����#73W@2m��l]�qIm�u��i�%��U�p�L�ݻ)x�M9�$����X0�j���VzZJ���u)�����{�V+V-��P�p�_q�����wZ�U�$�EɻBL��ׯ���>w��g/]����N�Mu}�ў����Es�xj+��iǻ'�O-Y�D�����=d�m���Hp>����9m���1а�����Y����>_�v�t-�]3)HD���o�u;:��ܳ>p;�2 ��w�iY]�S������A+w=�N����Oqk���
.e����4�w���V[12L�$=�yF��&G?���'�8U`z9��>=[�+tqH55��^{MK�}u̱ӵ�_����!v�2u��YO�я~t���ZSaJ�y�yo��#�x&d������"�E�~u��A*.ѻ`�Ȫ.H�f���4o\�Z٦TȒ;�ɚ�۽�������2i�)�H��j/�a�N����(~�h�F}G���ө� ӆp� �9����R(�	Ο���;�֬Y4�~Ն,��G�{e�t<2G��y/�62 �Up��s��$���G�@���GM��E���Y�*�E^�^�$�c1c�͛w�������'�n?�z	�!��x��2\VST�=�`=�4~`	̀�	\J��LAn�+�Yٺ���7ݺuΞk���W��֥���ij6��I�p{�N"UI'ł'D�K�� ��[T�&�*Q��u3�t�'^��T�'[	8��(<��{��p��⭤� �i+�!a���n�	�!a4����������=늘�`YUf!ѝ��kL�d}GE}��]�C;h��J	���i��q[��Eψ����9C�6�'!��@'�j�ysga����$mm����Fh@��s�Y�x�uk��T�	��¡px�������y���w�������~X��<��w� p)������/�Q��eV5H�f-�J_�ͯ��t����5?���o��6]�4!30�	�	�邤�ԥ�<�)n�;�̂�*>�ì��N;��a�c�pa�Z������� ����<�l$~�>�<�,aJ �@J��n�|���� �8�!.�<)O���;���|�HQ��õg�N�Q��.�=��]�p-0��a@��N�zp�F��٬���g�����s#�b�ޞ񓦗�őj1�(��VJ#ã;�������l׹4�l}ݞ���\�M������?y��R�V���������)/Ks�P~x���\*�b�
萞��@S�Y��⚗]�bh�6n��Qm.�<਌Bg'}_�Fo_�v��-�ܒ��L674�XC'���Z��v��1����׿��{�[�O����P���DQ�w�������ؾm��͘5��Q�Z7n�X�
q������޿������w�RNgb����k;��<%�n�i�_�}�=���|䓟��E���Ҧ�ޓ�*q�	|�����7���q[���3�<s�j�Z��/���q���"��W2��j兕+��ٻ)_��	�oڗA�@.;��#�;��5k� �5g�u	�S�L��4�G������#ǚC�Nf�.(�&%z���t~ ��V(�r��T��¥z���e�Fi��F��T�V�F���,]z�7�{饗��H���d5�ġ��L�E40�4P����̙��\��H;��$CB�9���>p�	'8��3���NX�r��Q��l��,ɑ���?�ޞ�c�=���O�����eҩ��]��I��(�;n�v�%�W��ƦEj���*�ʢ0Wt�����;n�>������Kg�F*;i��ڟ���u�������1t�׮Y?w�܉�k��cA1��o��$js]�Eqc5*�+z���^��'d� �k�>��s�k�X�0q"Z��m��j�O?}�ְ���J��9K�X )=jTK���L��
���r�3���k��C���EG��m��Ŵ��%��S��Z'�O���-��0���­����A �_	;�o���dZ&�d���������L]���頱��x�;M/m��@*[(��u1~�Q_�[%�9g�&�ر��Dx������`���q]]ݨ:`V���"��Lxʧ657���^����^	�1���W�"�W�N&g��]R*V(6�Uud����ŒA�j�*K��γ^�M��L�X)�X%m])U*�K�R.����թF�y�q.$�_�r�1��\Og�z�I�J�7�6��F+��b&]*�SE�xd��mߙ�k��������Ns��~���#�>)Y�,�
.s�X?qK��T���E?��O��Qg�gY��x0�M"T�Þ$���O���pֻC1U�uA�|C��dQ��{���|�P(V�H���@��iSu-	��k�����k��Fg�оM���N��mm5u�4L�$�}du��c���t�TN����N?s�8����/��7�|s���\U0:��4�\�7=,OHᢎ�/�\v�xʵ@##�BրJ�mmSF.��A���PvJx�gQ��US�}:ĳ�_ӾNĥ�_��Ef�i	C�����@Y]���ۼq���Q�����EyG�W+�j�*U2�̕(.U���J&�V�ja���F�7،��W�$�7�v��r���B'�Gb�����v�Hd֨�m.ʅ� �j��j�&�0##R]��Xպ¾����x��M��H��$ʷn�*5�!� =!0���Q0�r�c�:~��\��{�><��b��c�㛠�b*��p�c������}�g���okTK�,ѽ�-4Y���mcHS�Ξ5k������nƔhll����� �����J%u���_��U�T��^�H�`��)�^���/�L�:=]O�c'��� ��~���^��w߾�{c����M,�8m5_��)z
���Bx�e��:,���g�q��,͡�п�8kڗ�p+U`���^k4�?4i�$M�>׼i��-[B�a_�E�E{`��q��5Q�=��C=T��_�<z�}{�\x�E���	�J���K�e�L����cX�h��E!Bi#�O����?�Qی��(%]�-.�M��Wډ��v:�F����I���ڍ�7=���l��l-�6����'��+�vE@��j�*�B�YK�������Jz(�)4Z=#�é����#dV(��d|s|	���&�������F���v;"I�����d͇��!�hhp��SN�a 1�8tZ��I'�*��%v)��HF��+��əB@"E5�N�+%[��/�L=~��m�V�ŽXSЌ�!����]���Ǌ#�q]�Z�%�˰%�����&�^��cdH��g�i�7͏�Er�nD�M��h�&��~�@�뒇ˇ�j����\�?�5�g(?�$�\��!>�5�	���e!��d#xYQ"�W�Z�+x�R5��o�Ty�|���w�����j,;jHG���z_HHn~�#Y�2N�|����;O���#XD�82��$tn���t�b���iV,��W���m��Ep׿�7n<q��S��N2I>ܹ{ϊ+4T�:��y��#��%�F�z�����mo{�I���~�?�)~���1�\r��4�ǎ�X�t�]w�%�K�b�Z�O����#^�i��$T@i<B�ػR>��{@�k79�[�tmX�v��T�|�B@��O�#�V�l�)�˷���4�|��L#q�'���W��^M�΋	*�觧�Ql���ƾ,�٫�.�Q�i�|D7���7�'#2	�%R��J��ZMQo_т���Y��,�����x�;�L2��$�޸}�/�eERp���JbΛ7O7]�~=�}��E���l�^!��uh$	8=�QҎ������i���-���}�[n��`��;��w�:]X��I"UPIZS���N;��i7�J=���0�*�������X�3Z����)��)�裏J
�ؖ��X&٘��MU8��ު�]r��u~�y�O璬��«4�����w�4�F�?�)c�55�r�B�\�W�����ݐ0��y�%ڳ{�/��kt��K�]��h��S`�`�c�Њ���<����e)~mMf��( �Rol�o�tޖm[�@]=ݚ��}�;�#C�Ǎ'�����|�t¼y�|�'-Z���+4���H��"5e�W_n�o�����`^�7�67;�����9���׌X�MO;���\����0�v|cS#v���s�z�x�}t~_�`{{�v�1��v�_?h�nm��,���9f��P3���W�W�v'�Xl���Z����X6��ٳ)���c����_c��k��o߮�0�J�����:��5S��+(D I]~�I'	�雒��>�L�(jI*p>rk��g��aw�������@��`�K[.ױ�k )��"4��򷷿W�t.@{FzLQ+�ݒ󤲤�i��������F��8��]��$�.�g�2C�R�TL�݋deQ�5zt����@��D�=7,[8Mz-ed,zZV���4��-=�f��z_�ß@N�S�	��$#'���.�_����Ç(���w�"ڇlLt��I��+�̥�F��TZr$
��$.yd�T�bC��	��[^oD`���'�7㋪y�2&��0� :ˇ����$]#C��}g~��; TQ�H�0�U����>�[k�O;�!�~H��Y��*��(D����[n	�t�.������ZK��C��Z0�VM��:�?��t���~�͠]z�)�^z饹����}R���\ʡU]���9�O���7~�f��R��ޢ�������J�%�a�?�9� #s�U�\ٿ�j�]��l �jMt5�	&��Q�r�(�F�mT%5�����:��!�"c�u)�U��"���;wk^ᓀ8�<�>���	HVE]�c��t�+mV�?���}�E'��(�&1��5P�����u�֒��� }S
i���дi��y��A�ծ�Km@g��Q�P��I�<h��i{�u"t�b'�p�g?�ُ��Z}�p�̩#����?_JB��y�T?��\�eȵ��1HOD���m�.�w���*&��}�{���o�V���	 �lt�p�����htt,�;�Q]Ш���D��?�g�&s����|��p�y��;� ֫>�O�6�����8����/Y�d����7�9��M�R�$0��)u�p��)S&���W�������P�
.�K�t�>ٶm�&���q���޳{l�X*m�W��i���{�s�9��$S���?G�̔�����8�4Z}S��
j�4�7n��0���n�b���!�q�1ҩ4��+�NXm�ܹ��dL���aqHwx�}�=��BQ(�fL�@�@��6���k5 �2�����sIL�GN�8u�5k�U��0X��--��l\�D_��c���k�/k���궩���s �a��6�3C|3��~�u�x�	A�G
���sι����hzT��c����і}��E]�#c��
���2��!9d�(2���T�"���*|�`k�J8��?lN]���`�=$�;��H ������i�鴲4�yW�O�[<�m�ӑ�/X|'�S6���q�WV&�wħ[|)Z�]���Ȼ�{�?an�R���5Cr�������!$D��˖���l@As�����}��_qM{�r�Z��_�hG�EeN��lYD��h�Z�|yg�I�Z�U����I���}l����l=��S����:0�"�!Ro��KsU�6R)Dwu&3����>�������	�h8�i���ˣ9���X���Ǵk�i����87��pW�+c�w	�R�=m��Л��\��i�:"�7��!;-���ב���}M�g,���ԑ�J�:�\Q�i�Q�#�7b-2�u6�����&�G�٤�z�jb�)ϋV�L�LR��61��_����{��g)�{�����r�+^�������'�5k%��zG�Z(9`5f�k��ب%o&g�Z�F儒LĴc����/�����ߚk#��Yێ�qHRH ���M���q�e+krp}�`m����@�4dewq A��IЮ��L�8#N$��/_s�5O=�䶭[#ߟ��!���d���п�]w��"b�����c��uUO���O9唎�q��l�N-Z�o���?����+d�9�Bέh�\8.y��C��$]�t{����j�j�d���Y�ܴ�Ǒ�d5ne_������H=��U_`EPOK:u��8�<[\y啗]vYss��m�4���!�h�!�C�'�Ms�Zw�����]���-�Rv$ �_2᝝�����\q=1*��*����Q()�1v���r�ղ�����8��t}pRWo�.��D����H�Z�f�b֦�:aA5W�o�X�l���������$�2�+r�w���oy�9k׮�aÕ�N�4�q�!��x#�Q�N��\�����g���N�2qt���Ν;� --MD$�����uڱ�k�G�z��|�+z��*� J���
�((G���h��0���h\�=���=Vy���}���%^I�Ր�fs�'�����K/	d����}*:���G�]غh-��П��#�q��AW�R�S�Y�.ב�H@�&S_�w�ǲ���%���d�y9�1͛�ǹ~J��w/$6*�B69�ke+�����1�A��ᎏMg�9�����������T2��
hw�YO���ݚ(M�>�\���\+<)�Br�B��U`�Q�ĸ�딜G>9 �;[\����4ᧄ��E ?3�qY��U���J�)�ZV�������(�(�R�>~��Qh��o�����;��Z�Hx�*V+����{��.O����ZEφ���3n\Ƕm;���&M��l,}'�t���M��m��z,�����|�#���)ɋǿ�b��ǎ���)�x�b	:�$6�?4�K ���%���:6t;О����z҉'I�[��s76�by���Nr�9;��0�4 =a�ej=O�n��/��2�r��/�9`�U�����"CE�*���I_�E�+8�Q����>��0"2�j!�����|2��V�YC������
6�#F(8�:��>�Lp%��3i�O�s�9ʽĹ�]W*���~H���ntJ�<A��,�^ZH��qcQa�~���8f�V2�,z�����^�ijl�*�8�*C(�*2��
gXhg��K���L����DEi��#Nґt��-X�;�;�Ԇ4�n����������?����y�06&i�{�X�筋�~.9K�j�B�z�k�.g��� شi���(��ͯ�}M�G�G��ַ�U�ׇO>���b��"��q$�n��e�w�����%�\����cU��Ġ5#��^7�$-KʎOT��I�tN�BC��-`�� �xLNEl�<�?�xɘrHt��0"�Y� ��QQ��^;�qj·��7ndl©������[`N�S�6c�t������w�ygѨ����������B$������Zħ�z�s<�I��=�YY�%c�����/I����`f�}��u�֍��?�=�G����-[�@��c�a���C��iD�.Zk-(<R~8�bK4$�D�T�S,�u`X�C�jJ�͛��TD���C�.��2a8;h�?m��8Dt^H�s\z�����R�'&V�Q29N>����!�G�7 0������K���A���L���Z����*���r@`�#z��4g�U������1�<[�PZ<�!4�X�Z���K���A�RH/��S�c�8���Rq�gd���,(��7�F���`s�$�a:3�J���A�c�`ф�B���2 ��Q��B{��E0cA=�ڄ)��=�~d:�aL���4f���Oڵk7��<�X��T�Ei���=�RVO��3]�P�G5�ܠ<j_^+�xz��]_������M�d�s���BZ�Oq�:/Drq��
�	���2 #��U�-���?��#Te��?��:�,}�2ө�2�7�"���)2��(D��o��5rr/�S��4E}���C]3&��t�R؏�V��w��ݥ����>��s�
z
g�8�=k��r��#00
�c��RG�f�O�����ȷ��!l?r����$g9�J(Z��P#	��u�2�)=��RַԴ=�|9��7nE�/��/D�~Ȑvݫ{]VI[�Sm[��
o�~U�K�>B�b-~=�~���j^	>˦�C��jd�&֠c���F�q5r��R�Pj��	�h�J�m߲Յ�sV�HnuI�#��G
[��H������C�^�Yr7�}4�z~�=6�˨C
��+�E������)�3:4C��jڽ��.T��/�[��փ>�f��b���ƦF����|T����n��F]���\h�e�tS�T~��]�Omb�9�&+W��nq����~x�?���k��G�`�]!<�lٳ8!����u'E��:��{Y�}>�;x|�G,�3��[�Z�+:�-��-f��	5JV�5������&D Wv��t�F��V��g��y�y���~�?A����)�Nf̘!a��h�OYp��Ŧ�M�m߾Cc��;:;�ĩ��&AwW��/�Tc�����K�,A����E�Iʾp��'�Ѽ��˴�z��"��@�Q\�L�����~�����g��AGm'm.�
~������:w�L�g�}V+�V�ʍ�8��i�l�rڷ��^��D��w�4��c/{�a�xP_���H�kN����J(����u@�+�_��
�����j$�Ms�n۷�B���'�~�z�!B�B��.U����/����G�P������;�d��\�������v�t�?�c�+ʑb1��(�xάN�%/b
�B
�!�6�Xj�`Xi�=��CKuI%kK�/�AuQH.�a)�UcySC����p}�~5\b̞f	~~�;����)
��Ll��5NJ.��i�����l(��.!�P�%!�a��,x#�{ǌ���:ڤUq.,��r3c3u��6�K�!��R��Bٛ
B��`���Fi��5��o��K��Ο�+*�b���}�o��z��\}Օ:�����Y��$���L�$��]��x֕Ij��ᩣ����vOg�� "�P|��kC>���o��"}g���--'P��&���ݵ}�iS-8��!�R���'?I\��Y"��mv�}�տ����k�E�]ݜ R�z{���,y�Oȱ�n�	�#d}��׉�"��FIe���B�OO=�x4ӾhB&8��'�6Ɍ�®�\����i�q���Z����\�~�N�u9�VDCnjnn��l�*f�\���C���G6�� ů�ai*�U���"{��/	uN��Q��H_p�o���/�%(+F�5�~4�@�O�Z}S��8[�d�D�Vmw�?-�D0�E�hs&Z|jHTP��!_�+� �H��A��K�HH��(7�D[�
A.\��#��@�ƍT�;�a�zꩋ/�X kx(�A�Ƌս0-?�y�֭��Oܰa$�R<۶m�_W�Zu����Cڻw�C=T��'��r�^X��8 ]�O�$+�#E����/:Z��[��A�kJ��H
�Lr��3�&��K&����L��z=���.����Ϲ���d7QCC�^�4����֨�����/�T;�d�!�T�v��h�ʹ�3����ONaֻP����t��w>��ڷ�vK澋ˌ'�n�1S׮�(����5���^��N�a�K%����I��Yаd-�4$R�PC�� ���~. �+��|}��Q��^�Of���g��h{̘1mϞ��������F��LbN3�]Y���a�����������IH�mQC!�\z���q���j}�����0�u�V�^]��P�4�����|�]��l������n$dD�g����M���і��gR>����+��Fg�'hlZb-
P�pC�}%��ON��Ì� )#e�w�?�����X�S)�(�)���OGN��)*���)A[�}4´�d��8���s�ω'��Չ�wA����9��e���z��j�d���"�� �)�I�D��B�;~|G�8^TE�W=�D�`�����V�����`�n_{MBɽb���g���98;i#��w�9����ۤe�'/>2��D�����U��2;��/.�+����%ϩ^��§�֌�[��^�T�#�(x۷�Ԅ����fӗ]v�}��'��V�������x�0�
���Z�5�M6<��K�s��+N?A��E�����Z��ti}}�;�`����X-�!O���=�A�XpI� و�՝�(!�EnDf��ʞ�"� �D �b���L���Î��u��l62'��Y���Z�-�����+��\-u���-��oQP�RB#�6h����6����`*2C������1�2w=	˅p�/� �'d=FGµ���$�ɸ*k��ɾu�;w�?��I��R����u��M�8�h�y0�$B	�����i�P�ᑏ�ⓧNӒWʃP0h7�::ڥ�s�d��B�F��ߋ�o&xN�#�K�(Թ)޾c�����H~H���6@KH�l(!UZ�~�ԩSo��Fڊ��j��`�ش��=�=��FI�:-��y�0���q��K/�D�]M����J��8q�^(������mh�����J_��w��g?�م-�u\�4���,�];v�^��>�}�߽�re��%���i��B����t�	3��=���[,Y�D�����Z�vm�7�&(ZԘ�P�� p�A^t�E�!m;��.����
w�y�֑���Ңa��`�X"?F��}p��d�5�g�9g���#[*R��|�����'��N��56��&M��Od�2�_����\����.�������sqL��p�4`�������� ����>�SkC
`I0���"Z�p���pZ��Q��D��С�b1i.Y�jbI�^xA�^+^(��A�������	�
s�ڴ]�_8jO���i6���W\�x�b\GZ}�Q�)}��cF �,_�ܨze5�K�ڌG�>��d��T`T���<��y:?��Od�#ژ"62[V���GѰ�\�Y ��`�F>=K��'��:�lŭ+^xA(�6iʔ���jB/٘��?�ٍ�:����2R���֦"���px��e`��R�c�A���2�,�T�����t��a�Z.i�uI���uS]y����1��?83�vb��x*	Fy/�O�Bk���꫱u=m��V�e�iu��M����'��Õ3�'B��6mŉD��p������ӪkΘ1��������>��b�Eٗ�WyCFW56�Z�4��uG�qK�F�+���g	r%(��V�砯u@2���l@�iw|0�I����Q5P�����
�לH��y��߭����� ����[��i�6�-:]�Es귪Q�7�XY���'</��M�!1h��m��~�����7o��ak����q��ϝ#咎�o�Y;��'	����d�joh�XI�@W�P���5k��ږ���1���7�wd薜H4�_{�J'�8�	g�I��T}*=�60�F59m��P���?']_+AT�=9-�CB^��Zf���,�c.<p����R�>)��C�p>�c׮��ǻJ��Ya$?�k�����e�Պ��(��&���P�������#6>��N�S12ɩj��@O���(���nۡ��4e�����q�Gt@�ᇵ��B���fI:�JJ]J"��B���#���-�҄Q���-���D�֒�E��FY��q�ƒE���P\
�B�����իɷ@�#�Xc���|mza�3�8��~�ӆO�llt�-=�	�*n�����������$�i@�۝}���]w��>�9)BW f�8Y�ց�Ћ�,�D�B�s{�h�׍kC���cC���Y�O��LB�DIh}�ۡW�������Դ]�e�'=C,�K- '@IX�b[8?���<�L��JӞP�
p'�	Ʀ����t7\.}��A���O��?�Ӯ�;IE��6�6>��/�r���@t>=�瞫i��w���2F1O�_M�6���ԅ�/s<�^����SO=`�X�FI���{�p���xPw,Y���G�44�	�lZe�|�n�<�9s�T���O�����K�I�v���8�,ڜ����O��@ ֚=	\=ˊ+���hd#1B]Y;����^��Z.AsJC������O]}��e�V��VD7���zd�Q��ʪ.�q�é��,��T�^�N_[�b��3~�����|п��P�6X�M)�䃊�(�J7$X�P���s�QT~ [��"$�� M�6���^��N5zv:�Ι3G�,[KKC�T|�x��J�@W��;]f�&P�BW�N�/8P4�q�]���l0sH��H&�TY��{C7%��Ym�
9����
y����a�ư(�ruG�Ea�6w� �^IM��O�#���Q�T�pt���s�n[�,���JY�@��q����l�n�K�7>�E��K���������1��3���2o�'|+�9�0�]z�R<���E���	y_c��\���p���H�J&]�A��(�v�s�ɵ�'Nү���{�°s�jK�i�ޖ-[XP�UZ��F��b��vN1�����*�	1�DÖ�I���L�1I
�0��#�H��[s"CR߻�:C��k8����~	C�|'R�X(�zO�����a�f7H��U��Vq���%O���th�#�ݪ	e��2��7�R1�ݿC��K{�v��7��<b[F��G��gg�vF���N`�8�/��64U�#�����p��娪�:mʤ��zZO�.=�5�"ԭ�z�������ȷ�� p:5��F�}�]����V6�Nx���V��uVH�M:Ѽ�!Z'�W�M���*����mߡ�s�h��4�'�|r֬Y.]F�o�~A�1c:dv<�|y�w�����-�'�>i�)B���W�C],P;����?~lww��	g��Nl�x�ɹt����:�N�WFJ?�	^�Tl������k�����hB�6��+�>�J'-n褫]�W�W*�)�{^/�:�cǡe�y��υ�~��!�q�s���>t�W�.[
��N�>��xժUO<�8�E^����	�H��vZ&Z3�Ҽy'�#Q�Q�L�<���{��e۶mm4�K�"��V�����i3�N�>e�+��A�n�֭F
^��������)�ϑ|�/cg������~�d��.��y��Z|���Y�@W��GFN�3G��s.������B҄�YZɿt�/��-�@Z�=30�?vl����n���H+,�c��h��'�\��D�}c)�+(%�*���rs��������iK��g��3���ۅ��ɓe!X�g/'V=���?���W�;�<�8�E,���9W�)�n����?q*V0.��O����hN��+���^�,|�k�:�0E��PO��5��DI�
%���>��I?���5ͤ 4<e�fJ"=�(��/1"���ۇN߁�OW`������i����� a�����������3�NPe+w�G�ըB�C���uQ!�P��^xHJ��W��Hޱc���:�Q�R����f%v�g����cE|���d|#���E����6�,�D(��汨���y�BΙ���Y����|����K.�@K�73U� w��"�� �S[<��$� b���[_�T�phoo#�����1G|EPu��'Lp��S�L��e����S�+�,����H%��Q��O�C��t��:�L�������C��K�?�|����>�1|��_}�[���1�@����<��J�:���J�.ohX�)�"J��J�c��⿈�@�&7]��N�-W�� �dc!���|�E׃�0�+�ܰ��߀��:\�v@����P�)Q�	slTS��En�y�ݱAf2�tҙ����d�s�̊N�s�fk�srG�S�Ք��@��b��U�� }& ��矹X��-����h�����O?F
l�A緗�E� �!q�ZJH	��)iji%���;��`�ޞ>���������
�k� ��뎤�СM�6I�v�/6M!7l�P6�ܮ.��#��~:��S!Q��E�S����e��u8*���q
w7��XzjQB	���-�q��݇��B��ʕ+�ϟ�qj����&ʨ@Z}j~pn	�k��Nme�=�bW�۶m����/Uq�e�I�_�^x��ٚ��{\��@t�c���� Q���Ki55]$��[�9s��礱Gq�PI��d����H	i𤷓g��@v�X�Y�N�.1���W\q�+k�Z����/�|�w����׎�������r�c�u�r:M&�Dƫi��	:�k�6��C���O\}�պ��m�
��R�g�B�8���dZ\x���&Vs�-��ҿZ�Gy��3�{�!�^�ٵ:���g̞/���m�7���*�k���5��F,j��(�F��rdm�"�D
:�j|���Q���∪�H��Ij�ܱ#�%��T�VAR[��u�֘�����@AK�P�Έ8��{k������y�є�[�Z��>њj���zv��*e�i��P����c�d$ZQ���MY��66�� ?}�Z�4SI
���(���>�
�w��E��P�
�!����#�%ի��.D���#4H r�huMm�1cF����I:9A¯T�A�P�PZ�7��~��,S]�D��	C6�� ���2�^������n�7�-�VT1�m&�#|Fx1��c�Nu��?��ē�Uu��ϐ��X�̯�/k�4�.#8�4�!{2,\H�ږ�����iѫ�� �kEß�������ޕ�a/$|��wd�]]��1�L_�n�O2�`�nnv���uѢE=���}������pbC�5S��[f;Y��<���_�[�N��}�����[_{]ߔ��h��.���&j�
=��i��8��4�+\���v��{~�?�Yz��&+W�QH�8��	��w�J;
�����2'��ºcx�s�Jh* �la�@E�@��rĞY#pD3�ϚAMhp�Vj�pK�V�ݕ�5(����o���4��r��V�2�Fvl�O�fkֺ�_T���g2�TLg3�����ܙ*��z�]biT���nhj��}���p�9]�cr��An�E[�S��DI����iPӹwO5J(I�[������Jh؄rrF�@�f��>hR�߷@�Gk#���`_Yú����o~󛅄�@���Ʀ�������۴��]��7��IK�,ѯ$��5=}��$
�����$݋�-}(u.�p�}�����6hh.�g����WA=����v���R�{��Ӈ�R�G7�x���g��s�3��`@ ����C,�ի_tq�	u�G\zӭ��j�t�v2�!J�J���4JCp��{�� <�zO�D�[�78rP�īoj$dM�}ς�b����N4s̢V�=ɴ�fL�3�j�8W]ɭ�6�K�iׅPBdd`�'��ܳ/�,PV_��ey�j�� M\�8�gi@��`�%�\r�צ}�&<�m)D LWç�q�F�YGn��;�5�qΥF|�LT��F_֖�V���0�1cڴ�H$���&D0�Ja�����sJa�����o���h� K����� $��4��C�aժU�]�f�:���;[E>��4b[�5�\s챂G.F�ƣͩ�''��� O����੢�:|�Dx���%�
I1qR�7-`����ܳ��.�1@}c�����՟tʰё�E1yS5����S���ҰR� h�)����i�"���iR�]jY034�h|*�vs޻�K�I��X�HU��x
-�ޓ@F�*���We����mB,��Q�hb%�tM�,��w�I����V�B��Y��D�+�����Ir�1ʴ��V=uQ�L	���F���75!\���i�7p�;��?:)@��ꪾ$K��Ik頑�����ɦer\�l���>�b5[�:���2N粙\�Bu��7�=U���NqXBi�U�IpI�A��it����m�vh�W��`$;�, ���_����r�%�y�:��1S�q��8�e�ٮ��}S@�ٸ�ګ���?���[Ǐ�����_�җ����4��Q����k.����@��S&�F>��~���{L��&d�7�ؽ��&L_�;�V&�%BR�o�o�5e���R.�M��q��~�X�D3kcY՚����It#����½��j��1#��]���]�� �3'l ��;LN���v�i�L�'U�ے�/�H��Wc�Ԗ����p���;%�OS	�����AX� IW���I:�ʑF�8�SN���3�"M�5�c'N��o���ܹ��:��2�ue	#�ө�Mk�1��%�;I� �
J%�UذaÔIX�O<Q�KBQ��wZ�ju�������@�`��)�F��f�Y*{����p_��h�X�p����mw��W�K�2~<_4�_i�::��L�L�����O�3._����$��vp�*ܖ�Jt���I�m~UKp�EKeՑCC�;���(a�����5{�zE�fI�)M�5��$WԄ�.880�1.:�fΜ)�Ay�&PE�w�vĴo�U6��=u�anW_5������s����|���V2k5����Y�儶�����X_�7�Hps:ϐjc����T�?{�⫮�
.������L��=<Xd縝�ߏ��>���J���+]���O[S����"�#�?�D�Y$�NI�a!���d�  R	����R��	u��,]�T����E���5�~N�|�5����e_�y�晎��R�?��Niј���B,��:���5$r} �����Ie8�N V����$'ݍ蹉u.�(�l�e<�W���p;ؕ��O	O��݅��4'K�Y�^ӫ+h�2�<�2������ tm^�C��{s��@<���}�u�O840�ڶm�.;w�\8�����?Kz:G�k�v�JV�	}�.�3K�/�VH���@�74�b��E�ѯ j֛Dc0�O;�x���:�3fL�'BS�i�K-q͠(����\c�f4E�0��X�6NT�o�d�D��R��Bj$���3�<S?�Y��fϞ-�,�WB�֚V�2�1�-]]m�lY4o$W;�v˹H<�5)�؀;uA-�Ќ��5�\%��=�F���G/�믚��/�x���d��-��|����
�0�Q��f�����E��v�	s�/J��Gu��?��(�l���>��o|]�02�V����>�6'߫Z�4�����	��Y6o�|���|��������=}	^�L> G>2g?�DM�7�.�O�(�}C�>�5�����eù#6B�&���P�����P�.H��RvLy��0�֯��|!�U};��΂�³���FU�<���Xl��Z�Z�ʐv�|���ŐCm��\}6��׹WS�6j��Ē��\�={fSSú��k'LpQ$Rt�M�X^:Lq�w��Q�ǒ����I����,b�����\ס�R�é[,[�Lcnn��E�/� ��n&t�[L�hC�\�R�32T�߮_�^���ho��ګ:r�<���
�%�Nd��F�[*DU�K��v~DW�PoL��Q.RPd��5vi�S�{�9�in�A������ϟ/A� ��`��ه�Y��$�v��N����k����vl ZC��ڇ�;��N�d߁��\f͚E��9m/X΋��K�����S���Nߔ�i�
VM���^��U�	�`�Z�&��NYKu=���[��V�P=}x����M�����#�U�u��/c���mm�Qc��\f<�]p�;_��H�#J�	�h���#�<���%P;��D�)�ܼ`���̙�Ie/-�G[�ۑ_
y�j5��x����1ܿ����X����A>�@+I��JRTh�+�5nug"��^�Y�60���q�%�;�S�0 ��'�����BH4Pb*ఐ�q�/�B�Ց�p����F5V�j0C�j��B���s1l�2����$��,�	0��6cM���z
'il@,PE%$vH��]�=�0�Z�Z�诮r��p|R��i
�gLsHq���5�h}�s�&]U�l�8E$Z�D���T���	@�:�$n`���M�8�Y����J�ʄrt/vu����ӐYA��=�� �|�'yu�4(E(���O����y����AX�x�����9$aҒ3N¤�rst�����ߪ9=*K�-$���j�3��.�v��\z饎8Ө%���M���z��z��`�n��xP��r;��!�&��8 U<eL�?N4�&������+W-\x��ؗ���ڱ6�Qph��-�;�|�:+_�èZa)��o����T� ��C�=G��!e��[o���/lkk��s�KÝ��$�[7�tӽ��;q��}��׿��\z��g�uFd���PWWq���~��_v8(;���颋���ڮ��]����QoH TADoL 4�l�c�k��S|{��1��{��yd�8/7.�㌑���%1`�L3��&$$����N�g����ק� �����{�2������_���®��K�k*U�Y�j[�_2&=�VX�!�/�ʑ��3.1Bj�����E�Q��ڐ�����v�Gׂ�"�e���(�4`tA�
Q5W��=N�ΟeŋQ���L�^�l�vK������}7��W�.��S��\2�$�&�[��*�%�n�,FqFT�a�}�)�i�4����f�KW�R��[�Ks0U��]�[5�)����m�ok��P�$4/q���7����/�h�6Bk*5����RY-���C��q"�Q?\T�������$tӒ'&��������u�8���^�ՓX�k5x�dժeǏ�x#�	FϢJK�D�Dl�5������
$[��}��󛧞��������sY�K[#�ujfZ�J:f,uOz�vD��D��)��I����?"�3ݖ4j�/AI��+����.I}��^�E��w�;�Z�x㍋��J&�b�k�kK��6Bw0������Mh
Y�<1�⊫�R�l�#`V��W���kZ�f�����w��X��,�^|1�18�xe8� �S��m�n'�L���Q#'��Qu,��e	H_u�UR9y�1착�	��Ԏ{��M��J����oMaY凶2N>Eij �x���a=����k�u�i��,뼋$tC�y*�3���FO\�l�Ν���H���q����^o��W'�vn���?���k���&B/�����n������~�^�y�d�Ɔ�D�"�[n�`-�ވ&��hH�K*_/����|���L2C��($p��\룉�)�g��n�_��E�c��/�}���<��y���<2�I�բy�~��2U�k��Y�-�ae��ޗ�zZ��0��f Q�yP���#�&c(cP>im�:�aj�ė5r⒔����ɒ�ʡ����V9�ch{5+����֊��=���g?��OP��߶����\y��;
�F?P".���̶����͛��\�5G�vt�_}�կ����kkk^K�&aNfɒ�1�n�җ�t�؀�JZBkK�)��Ë}Q�Z܌8w�D���B�z:�#ݵk׿�ۿy��e:�hZjщY� �B4Y��{�L���A�]�r�N�����C���v����w����},�Jo�r���	-���hIE3������z����Ȑ'=�Q��2�81�s:=a�ei{���V���WPc�o�y�~�_D�$ń�����7�b4�Xn�Y���2q�n��0c����=�Lw�g6�SŸ�i6,���X�Q�`�b�J\�\���Aь}f'�Hj�d�s�5��Ѥ�RRXu[K'��X�T�w���*U�|��4Ǭ�j-Y�R���t�-1[+V��Ks�|:�o<�H7�+����L~ve�ё���Nh��V���[(yf]�z�q������՗^7������X���ti�l�m���ڪ�@_EP0�d�'j�2ɨzbh^)e@�aݦ���8q�Z�,^�h�������������=_*�eCu�u$�������Ç�j̅y㕭��=zLp�g��3E����ji�6�����O�FBT�xtt|zz��Z7Wlinӯt��I]$bӎh�+�ʊ+�]؟-�p���E:����T4�;�cX##C���`֛�	C/�.��Ri��>��X�qOG�X�t�Љ��|���w�H��Y�+�!"�Z6�m�ֵk��'ZU�D:�����#��G��N�=ydΒ��H��L�zK��}��t��W�����^'c�K&���A[�J�.m�pW�(�՝�w��orrJ�?�Ȥ��MdiK�A*�u૥L"Y��ϥ�%�!+�Q.��^*�TR�$ZZZM�hi�xڻw�s�=�!�{��~5��_�3��Э$�K$�/���J����SS.44�bQ|�.��p�;�����#G� 70.����DWo� i����HxA���X���;ċ�^��#���h}}�8���ۿ����'?���B,�W�����
Y��i��1�0t�N�k��n��H��T�$�(���O~��;��S��@��tiT�!��]w�E-����#�3<OO30s�ȑ�7=:��|.�i��){�Ś�z�=�7�p�'-	��F��.�Ft=��c!��p�%�В�F#�G��e�xp�5oqS~zn6�ܔ�׋f��x�t��F,�vfjZ�i1�-���~`���Ė���� r��6:�ZzxdXL�`����(55=�r��CV5_����lF
�edg�͙t�Z�+X����l�Ţ��-�ӳ3]VW(���q�wc勨h�,��.�<��6"������c��e�q�ŋ��K/�r��-Om���/�ʋg�4�gyG@�!��z"��CD��r�X�:Vg�pHg0|������>q�W���~=�����)w�髏=��ҥ_}�#���^�6Bj��>�xԽ����/��~�С�����&�hq�9�~��`�&ڢGq2;N ���{�����������o�Ú�׊��aD<]]9�p�ʕ� 󎜢�MLNf8}&�5X�v�m�}�o��o�.�3�Ѿ�%K[������1��h`�e%"� �˭�]��Q�+�5���w��k眻���������v638tb��e��������}�{�w�sOO������n�Ȁ�.1h���߻�v�����*z;�2Q�ɦ3!a�T(&�DK6��ܚJ��&�K�P���"�Go��":��OL�������c,�����	�8��k�"W<-�M:Δs�O�аqI���[uv�����B�[�ƃ�f[){�n���Z����V���Z@����n�}�����Q��72�ݻd�G��63%c�M:0RT����9��U�q�O���j�)П���ꪤ�t��C	1��Δ�a�f�|s�P�,�>��-d�-.��2(�\N<B+%��p�bR�=Ν��ٺu+���7��\��W�e���n�֭s�`-��ρ	��4��'��z�zI��BȦ�!�K��ؓ䮖�ĉ!b��jh^����k��@;v��a<-���M���̉���%���!�*#�#�IB�ꀽ�"%�q�=����O?���t˖-t?w->��2��F�W_s����V���!��\�SX����L��e�]v�?����h�����/���XeMn�W��c�ZJ��w���1�Ej�Ъ�5��Z����h_�{�}�PBN����+�H���رC:rm�\\�ʼt��Au�E�B�wWw���h��e��d��R
'k�s` ��_�SfB���ҧ�yf̃���Kd\x���N�!q@m�l��<���"~�Y��<~\��z�9245���7��B�-����nX��Gʉ��.�n���GM�~�",&]<K]�"��E6F�'�I˖-y��祜Q���B�����!M\K�aÆU�V��cx���?�i�!�0�5�ё��K�H���\ʀD�~4e��$�k���(��dXP/���J����UF��o�.)�ը45�I����h����dPR��	j��$c�_�9��XԂS�Id�:��[�gw�,8���=E�v���p�ꂱi�1��xe�q�غ�<!4Kv��kH��8�<�IKH�+��۷�#�@���RL�%�((9�Z݁F�4Y�25Z}�~�:=qH*���2퐊|�tD�䘋Nd��'�x}u��q�:�7�|�� ]�Ja�!��x�W�N�ErޣEu7�E��V���k<ڋ�~���3"*�_�U�;Izq�(͈J^�6y����7J#���݇�K��0S���=��7ɸ�4W%���THme>���"*�!�� k���zg\�R���o}�[:�6�XD>�����z�߲��=�&��sy�4�A2�d�HC%p�x�B�M��J뒠���=�=��Wiz^��W@����5��	dVʛ��8��C�i�pƓ!���&��զ����I���HZ��?	�X5��>�:N
F�7ׄ2!�?���u�l�{�Eq]B��mb����/H�Z#��Xf�8���1fOI�ٽ���H���]J5DH�e@k����埦�W<$Z����q���,�����N�@�<�9��c��͒��d2ܵ�O�&ћ�-�\2�5fk>o�Ӯ��w��&Ӟ�X eNs��צ���K�kv��N�F��a��F�H���$���$�P���9�d������5k������	br�d�^W��o
J� �X���g�5�^O/0: "�E��E��P����jq_X}�`A����=V4J.��%������UFb�����=�+b�G��_�~�fJ�
n�7��<�H�׎���ftb˗�ܰ~Ӊ���	�¡�=�5r�'�|�I��R(Ҟ�p�%!�	!�k�Ȇ�oI��e��Dq�B�ͷ�ҡR�N�~�a���k��_�v�g�����X�}�۶�t�w���[o�M���W��@����ݩ���d�6,�\�ʕ��0�,y�����׳���#����)ɸu8����q��Ŷ�#Z�� _y��b���� ���{��zW�Ն���I��8~^�¹FG�Hm�@c�(F�ѣE�L�[��;�`�2ѧVΨ�~��/v��N?}���п�˿������	�I�}�<��Z����W_ݭ��z�][[�={����;�OY�C'NH9��ѕ�����!�*�"����8_0S�[��dvt#LK�_�X��[-�>��y�9?���+Ec#�T0�NP�HG=B1"��	ۭ}�"C���Ydv��!
Ƶ�<<X�4q��WC?� u�L�Tw)�;�h��J�Z�Ě�jjbh�}�=^��
YRԉ��D<��`&M�"�PK���CC��ED !T�7�����.&r�v�R�$##�t����ёI�"�^z�[��n'��T��(�)Z�v�\��i`3�u-�HzU��c%Q�dAr'0�AF/;:�&�-�&&��+t������7 u��9,&�9���ӧĘjq�C9n��Ʀg�����o�yH�`ڗ�L
�"$CÆO�Dy���`��v��I4�:D��OZ��M�*5�sLM�m��z�hD�>PHS����i��3�JW[�Z'G'À<�g��r d�'�m��&�N�&�Td3Q�T(�Z�����`�J:>�xJ��Lj���Ҭ0ҭفT#����i׌��m#w0`�+�|갞�b����[0�Y=ٱ�WcH4W�"a�i.G�d�Dq�T���fӹsY�$^W�K0!-�/;?���z�D<�11��a����7h� ) ��������1�ʃ����ij$��2���9Q�Z����Ȩ�#. �݊
�y�? g��0t&u�n�ᡇ��_�'L��q�L[�^�.�H�)� ���5����xIt����j��z�G�ꢋ.�p��"��~>�dL���"�(5�0P��[ԇ2Ia����/�=�����x�$$��	t'k�4N(�e+uRo�j钰 얯\���W8	21z�Xƴ�O0{n`���\��/�n�\}�Ĺ�J���;�Dr�I�z
�v��r�-W_�R7%��|��ZC�1�J��}��\@�2�<gݤ{���w�]w�رcÆRى^�5z�[��c�!�4�
]2�ڶ�T����O��Pn��ƈ�L����}�j�
i�ZI�P��J�R�D���t��z�E;-E»*�	�B���:6��bu�2�y�֭E�Ҙ�n��֭�z�Z��X���C_��WEQ�c�����Zka\W��m�v��J���-1;;��o|Cc��nu��ɤft��7�V�s2<t���=9$�ŉ&Ij�9���c�a�͸Ot��7�� @_I�Zɥ�7ɰb7���z�r�19�yWF�.FD轶@v�Ī��{h䔎��M�����B��\Ѽ/���-[r��`�y��B�OB�zO>��u���C��f�Y�/;�O��$K��F]M�j�'�\�O
�P=uq�8�bh"6Y_b����Ӟ2�4�@c������<VO�lܸ�A�� �k�z�>���jn$ړ\�jh���㶕Q���wT��%ϲqo�\>���ƾ}���|���͙N�MT1�0�����S�A�mD��ʋ	���?�я~D��w��9E?{G�'8H�aP	Ts8tF�����;�i�;�d����]��,����ܹB�<зZL�*o����KrR�S$e�u�l=��� Z���O�P�>,VF����h{͚��Z�w0F�FG���'�C��ڌ��<�Ũ�iW�8&��W�;�: =-x[�u�S��Y�L�O��6N���ޠ]Eq.u���+ƃ���@�Fβ�z��d�A�Ϫ1�Y�⠴U+q�����;ԅ����S����e�Zu7��3˕�����'�e�ؐ�k�e��dT^=�H�{F��G7j:��O:�r��6&��j�Z�,��MCe\�tE����Т;�J�%{����vT�5�Z���֒LD��b".�K��R-�#P�[�EBN����֭C�A��*�H\��� ��[C:�sV�\��ۗ��
�B�Rz��/�&&Ɵ}�=�D~G�|av��,�ܱ�SG�����<�&�O���挠���B2����͛u�t���i3-�-��!j>�i����� ��$�|�^SqI��/Z�ώ�N�J���d����pOWWٱ1��g���a5��mXW^y�U�p	T]j��ү�y����h���24����K.��h�t��\�all��v�j4Ҁ��q�� m�q�	J���)���?����ɩ	ݙ�mu�_���z�V��o�`hA�p.��O2Ig<���J��d���E4��*���q="����Fp�K��2�%�Ө�_��Hb�����#�<����Ķ��w�����֯hW_�F*�4Nqd��e˖�CCnD��3 ��F��u���aA�����KR�ID�}��'�2�����FH84{"YG��oz�f���|D���I�A�j������?�#7�kSݩˤjF�`j����H�!]&���_}�ղ�c�q�p-���=o�2�cC-z�]s���>{�3N���	jj`�"�y|<r��Y��P[s��
�3�To�饎��T�=!�T\��y�F��c���$0�N��=�r��?���=��1�9�Y�Y�`���hjfzxt������W_�����n��#�����Ɲ���i���N���u?@HZ�+_��u�^XȉMג�i���krj<d[��G$��C�X����������ƹe:Mc�Y-�nsq�(.1�/��Sv�;����qmǲeK���6$b&�"�L�B�N�f�������~��2T�߿a�F�w���r���8��x(9���$2��^x��D"]l��M���zO�P���� �/������+��r��g����}������n��Z��i�����~�J�\?��3:��GX���"a1}3œcc�.��ȁ��d��f|`hW�X�����T�-�u��#��d���#.K��� ��z�T\�Q�c��I�p��q乕�,���d�p���8I�P��+�6�C;�h��j���ꕕ�T���X=��V�� �zQ�0��U,'Aʁ�������j�I%���)� a��&3����'(�/n�'�u�3I�Z\�d5��@�qvf���XE�������Lើ^:��]�Gp(f�L�	M���KzҡC#�����~���F��$�	�2��ԏ������hן �Gnsk
�tCo~}��nX�j 0HMP_��g?3�9�����D.ܒ�h��T}�k�.ћD8��������N6�~�y�t�c������]w\��[��
|���ն�n����nXwhF�ׯ�����Y���U��<��$������f�;�Q�T�H&B��((�J<��_|Q﫞A��o�}Gg��%%O�$X�;��KRGk(�@k(酠��ѧŶ"�N�+��ԾJ��j������5���}[\[��%��̹�t(����缾O�Ӻ�����GH�J፫�,��R���XW�����|�A񡬃��wt� 
��lڴ馛nz��4f���g�mۨ� �_�#Z�m�2:"W��%�%e�l8�)�<��0�o����"*�/Y��X	�)ӿ��bʐ�����}�]CCcz"8�W\q�n��o|���To�j"���vS荧i.�����Շ�Rq�0�,js�V�Y�i�z���mƛ�� d�S�i�����o�d5 Ԃ��h0�!�;Wo/X���%��j� �<e^�\�$xi��4D���x�,&08���T6�6�?�u
����a�C�ӴnFTK���zG����HD+橴�a�aFQ���vٲ���V����2Y��ګ1�J�7�O1��ζt��pG{���z��k��F�!&��;=f�AKk�$8!���ZChIO_�x�H�_��_�����+����U�o飚�7��DF�Jn��Q|O�ӗ��e*��1x}��2 z�W�3
�b2��?-�%���%ɸ�x��hTd%"���;���y��ub��(����~�!�2�F���h�ّ�*���c�]r��M٩)kKM ۄ�\����i\
*�%����9��Z�]4�s(XXZI��r�@�×�E-��w�d}ww�� ���:�a��?z�'�V�� !Hx>e.(����Q���KW}+�Y���g:���'h�Q�/��ȑ/�w� ��9�#�����D�T�U4]<��t��	%Ṭ!��/\ #�����´᜜F<1�L�0wbpxxhrfz�X�$Sl���C-q
����kP��qEQ�{Pv��h]�lq>��w�:�cn޼H��4#�B�*�wɒ%�"G)+}�j�������Η4��zܺ\�^,�+�D
�VA�>��K���?�ɏ����jIR�e�9�n��G?z��:�(��3fv饗��N�Y�됓JZ�R@ʐM�{��������p�t�	����o~���w��7�d�	ZC��6�Hz�n���i�婔�%sTxr��+�֖�*0=3��׽����d[[��trrjhhX�����g�^��,��"��jZ(���ٛ=7��霍��k���ȱ'�N 5�u^v�a  	oq$��������* �ocG����G8p@��6������(  ��IDAT��}�=�!�&i)��VkF�"����)�%��K
��r�I=T�G?��4�?��?��"�A�����'%YODG:q�����k��ZIT�]�Vg�4i]�:wB���;;;�U�'Q	���F�^���OW�0�r�~ݿ�2�a
r2P����<��2���;iY��]�l��7�9��hC��#�uֆF}�QC$�3��q#ε����/�,��Z��EE:���Ug�YЩ��H�*��?A��`:x�s�طƳf͚I���� �D���$�G�hD�����녳C.yi+q�U,����T��O
6�u1��Cң��1Z>+S��8��u�����=�չ���Պ���F�X�Ue#MNO�-��${4n>��W�����L��6��Wc���HŹ����׷Ҝ�;I�4�[ �s�q��9`���Yt�$�,�-��U�������ĺu2+� �'�����Ջ@3��6�@����Ita\Ǘ#��6��ǔDg����~\��l��n��������=+1�B��h��� �1`{9n,�o��2�e�._�X�)��x��_M,�\.{�u����?���6�RC�iǓ�-��)_�.
�W���/~!Nx���&�GU|�VY�kn��f+Ւ��e[`��=�3bRCC�V�������b��,3�}
�Y9aU�Y�ȸgw"�l�՛X�#�g���i�Y����K�3�z������-&�/v��3%b��hݗ��,�rݣeݖ$3^�i�JuI1�u������߭���A2I5is��.��ۖT��d|lD���/����x���
h/�VS�s�3%�[欍l����]��y+��#�T,�I������p|���&9Z��B�Bq�wt�gj^�dæMO>��7���9��@�h���h2����"3��i��I���Q$=�N��|H����5bC�9����Cݽ���G>�ͥ\I���
}�����蒋efi	�z�))g��{�]�5��O� X�Q��}��ĕ�i瞳����b�=����UW]�������S��ڷo��>��-[�h
�X����ڷwo�C��1��v_]D���B�=��v�����I?����IJgٻ/�  EM?�������w�4=Q�k�S����a�ؙ{5�A���8?x�]�m�]��>r���^+�̹����vJ?�W�ct+mn6����h@��>�W�$�������&�����[߲p����o��ccg�]{��w_p�۷oh$�k!�i���a)��Z��{�L��wx��Z�q��w���g>#m��,�-���7H9�75�����>�!���P��3G�҂���'��R=�����<����sZ�)���Y�kH�4d�9.C=��ǋ	z��!h0�#@o�o���������<�g�y���	kS�}$;':)���/|��]	��O�((�Rb4��_�_����Z�E:�T4q6��W�/��>qKi��'횈D���z�^���O�(�`ZX��်�ߒ�!����$P:��E|YT!b�y�9�7�ҔW�\��B��D�Ш��bG��n+�
z*�E��jlZ(�����ӖQ;���)on����[x����N��iVC�r�9�2O����؀�j��U3N�x1)��h9��;�f�-m��$��]�v�`���{z:�CdR�NT��8ՈߢOT�'��C"��؋���'R,>�;��0�#�,�����9�,�&K{��9e�h�����Vr��������	�Eq�S�hȖ��V�˼���?*m���^�����ZP�B���Gj½�Ԣ�XKG���{��.xox��j���Ny�q��FF��Fc{z����g�����U�����R[��~��G���� �^1\'(:�홸�9���}EC���V4l7�f����$���S��3g�3q���%��hP�-y}f��ݙ����R�,�w�gX�־RI����M�q{�d�t�d�Zp���E����S���6�˗-Ѭ�J����z�<���a�ۭ�H���Π]���fiK{#1��;����t2ai�X[G���Ds�5���&[�Z�;�K����d*ӿhq[gW�T�кW�C#�Xl	�)@��ÑJfZZ�(�3�"�)h���Řh^.ֆȁ�
 ���ú�2ɦ����q�_�`��Ը�S���R�亖�G?�ᣏ?F�F�jgIČ�<e/�o&c�&�D�eh�M�`�1��%�����|��Ql(�3�`���)?]ո/8=-��z������| r2���<��Ò��D=�r�;Xg<i�2�99 ԏ��/_�r|l�0/�0L�L�s����-��ID�u�Ç���s���g�+�(�F��>ۄĒ�˘ ��X$m4NMV���.��|B�j.C'Fp��?ЎH�������D9o�t���?��s^�O�D�֦���GGǞ~����~���;w�߹�zQ�hLO��v�g����馛}�1�e�h-�r�����<��U��
�h3ӋEC��r�y�{���/k�V`1=Mo1���Ww��g)�_.k�1,c����֖���O�7�~����U�8/��c^s�RCz8&nl*o&��P$�t�;��O��O��Mx�W"xǎ��67��(�G��.��r��d��sF�dc�즗��,��E�֟X��7ވ��(��� �5�����#��yf�F���sM�
���S��(O{�5j����^XĤt����G�N��P�L]���$�4��Y�\�멃#�M+#)x��qҿD{R�+�Gj�N�Oh�t(t�U�ĉ��>,���	r���I�ls���S��*Q�B�*�,��ѫ��=G�Wh)&�JeMk��)�eI�bNiƚ��4 ĩ�Rh}t�c7F��k����WM\vװ�����H1�dAݱ?�6-���"8!�5�nWW�g>��k֜~�����$�ܣ�s�%s������ާ5�U�V{�L�$)`+L~�L��O}�SO��7�PQ�7JqS����q
9 TkiM(c�s�(�-�Xe{"E-x���Bn�H�Z�����9t���>�f!:�֭�����X{x�6��ٓj@����w��ײ̝CΑ��S@ע�C�����H{wm�j�njF��)�A�,�+�s!�K��� �B��[��+6��TD)U�Y�N�bcjP6�#zƃp�Q�T����j�Q�P1�*qf-��t(s���q1�Z�r)�Z00By�u�Y�V?��#������6x�c�-)kn��zP�X:�>#��2��mF����J)8�F����Z���n[�w�1.9aV��������x��!-,�+urff��з�0z�G�;`<�����J��>'-T���r��ҕ�9����Ž��������<.ʊ{�E3����PQ\��l��%�MG4En-���~O�8�4m����?�����3��'#���˼�����Ѧ��Z�	�\��רP��#樇�ojG�F���a�2O��{\�_X���  HD?>�<�D�{�ȧ�?ix<a?�B"�l n�Q��R;}�Sa������ne�8r�<��zܚ5kJ�Q�c�xSճ�0�������}ŊZF�d����3eA�~2�M��:2<ܿ`�����cd ��"酢1�N� 	J��P�t�ֳ�������k�k�B�6q��À�s>�^7y�r4�|��(Uw��$Dqk�Zشw_��S�j"p=d�+���^�C�,q�{�S�UFK(����t�N�1D�zO�]�ȭ�Mt����*m;�<�Mjs�~����O�'����г5����wt\u�U�/��)u9� �`������{L;.�E��w��]�ͪ�m����p"i`�����P�9�@��J�iNP��� H��IQ�	i
s��X"��#Y��U�����᪫.߿�0r�R�^8��6˦M�ۮGht|�
1JU��h�iSw������I͸4Y-��r����"�����5(������f�+�v�����h�����>��Ҙ�rHK��ѽh9ħ>?�=�'���|� #�4�ni�P5��أ�9����z��{G��Q���hA~��mݺ��,944��l޼Y���^ra\Gм4m��DT4ͪ�M�<��7<�����y\õ�<�FGE�*�Dqh"�,�ȱB:����8�-�wmJ� �  ��!D6��G��Q�ߐ�c�L����ީt���d3�z�x:}�����W�HJ���HW �F����f��/#��X�(ӕ���kJ4ĬC)+|�J�r�3��SH���ʎ�A�����ZZ2�eո�2:=�V������uD�n�"U7�}�>�ȷ�"���XF�Ta�~5n�(���\�C:������px��H1U=Y��;a����F�@�6�����%;8`"OF�U�LOY_�Z��/>��'��U�?_�T�ߏL�(��rrjjF�vlr�\����H0A�^"�&4em��Ԕ9�ۈs{ߺQ���34+ڨ��|�ǎ;�7�>��C�����5�9xD�D�C��K_�����O?�N��^×YV"Y�OR���f3(Rh'x��V��y�%�}�# 
عsgGG�������$�8�F"�����<�Lٻ�k���q+��\�RW�8��a����h�{���İ.��2iTz����*�x㍿��od��ڽS�����e�{��a��N�v`n���;�S�}||R�����R�-n��u�OL��P,�\|ǲ��D�9r9����e�T����V)�S�'��� �Z�A�H&C��iD铄�h��#��S�[� �j�8x�H ٠GK��uk��y�0h�L�Plim���%r�犳3�,�VL!а�pУМ���/���;��ӟ�3�܌��e�z�b"n!'2�0�lRCCF+��-��r������D3�&����<�����h��sS�ޞ<D�Ee�͆�%�^�� /���q��a2d�������>
�$�s�%�90D���xt�7�p��}��g%q�P�)���׾���O7yv隒����mE~�P�M8�4�Z���~����u�fCV,���T+EJ'�Dʐ% ^��X�!@h.��t�)"��B$H���o��4`�������\���$p�?i`
�D��<'�'ℨ��'2ګR*K�I�A��J�i��ҿ](6;���K5%�����J�f��oO����On=[��2��V\�χ�~��M:/.��MG4��&�Ap�}[�AU�aI>�a`�r`�g���[�n�چh�b�M�<H̼����K/��{̇�MCԅ�x��f䞳��] X�����7�}�'"��k�b;v\s��j��i�H��#n)�X�������Tpr��oũJ��F❐���^��jG^|������w�,u��Z�%�l�}?�r%�����x�~w�&�joû.c }�E�J���n�W�5�r�>���:]��t�}�_V3暍($�A�;Y��N�2-�y�La9F�;�N���[�v�L-�]U*9aXÆ��ž@Kj��=��%���"5�ٕMxI�!�{��)hq|3�D��� W���52)�����;؂b�
+'>(d!o2�,]w2��R9��8\���&ce����Q����>�� �t%�E��|�9c\�b�	Zsv����x������W9����tYEEa:���cx��U�4?ss��}�y�^h4�h�w�z;�Q�,�'-�$@$�}� 4AGQ�͜�o�x0�*^��� ��}���r�޽������?��z���G��7_k*�Y5Nt�{�6�UPɯ}غu�g?�Yi	�bd��1���袋h����ژ��SN��w��7�Z��$�˿�Ki�Ǝ;�nbUd��<�����կ�=GG̚c�;H��'ɺu��xc?��K��R�]�y��W-�(Vn��INc`Ы��L���++�p�+���h�  �'��f�rꇆ�.o�q�:;)s�?i<�Ɂ8z�u��*�'����mm 1��\�D� -d�'��A�7ox�á��Ց��c�[%ZG��eG�_�h�G1�_
�m�����9��'�L8v}�,�;?��PR���>����Sg�_�{Gf�Y�\z0�pϱȠ�:[�j̽}ݴ��,�BK+RZ�x����e�s�'z3l4T�T�_n �� �e�x�H�eZ�3�<��)�o�� �9m����۷k�C�SS+�&�Z�all��͢"B��k)j���ҥK��!f� �	dS�W�&�S�Q���p�y�'ND�od/Q}WIm������J?Ӱ�hm.%N���K��&�N�Ls��!f��s��<�3D� �vޛ	i��\��J$_�����s�{_�౶���K֬��!�#\�h����bRoB�B��I��3��$x"7�g��XD1���Uţ��V�롇buO*TĤ�d93���� ��Kñ�)s��r���5̨�����!���ZC�}���X������o~�۶mۺ���w���z3YJz��	3�Kh�a\ɒ±i�&- � 郚X{���b��d�Av���~xϞ=7�'I�lˬw�lsU���7:8g�u����RXvʻ��jM�N��ǎ�i��cc�����j��)�v�2Y�z�2Ѱ�1�D�	g-�d��Ņ��g�FqC|�}��8y+đ�{��㤟hA��¥�������Z�4�@"W(q�4[��G���P[� �1�PF2���L֕�z�3�+Ck���Ɵ�q���7yg����Y)@�d<�ֳ0�b�.M�/�'��u��U�t�Ok͗�\��_xF��$�o?Q �[L��Sf�5���s�|SS֩�NiS�8{�)�x���MLO͗�""�0n�l&�F�FeEyRa���f�h���i��P��F:����M����������^-�m�/��(�72�q�W~����~��m�azjVʘ8�u��ד�Y��Oz�ڵ;w�$<J��]���j����E����@g�(�����F��p�l��K.��C��\ �12<&���e)��w��,ļ����)߂�4g���F�����北��/�V�F������ں��KW���b��X�1��%�����;�A�H%3!	 �5��O4r��qO�;�ӊ��;�|�)�����m`�p�A�א$��o�J��-u�-]�\��q7�&���95iO?z��(��3חѪ���ն^��w�~I������{��w롰������.���@�L��f��z��?�aQǕ��|�����܁56�Ù���Swp����$�:hsɷ��z㍽�v�:$�d�4�n(�7C�MQp���#��ms���(D� Ƕ�����^{M��u'��G>�ő���G˚5kt|�\] ��
:Ȥ�P�z�1�P(����V��-ת��8]c���O÷�a��LO�1<%��/�>T���-[�N1�K��¦�D�D��PP*q	�#sqS��Ƹv�o�$�u�*���h��ȥ���H��F�(��Y����k����`�sVi���g��7�6����1����9`<�s��J���,�(De^�BuM�1���!�J�b#Z����}��pd�i��֍^r�C�ҿ��c==]W]u�X�~��1�	�M0wO��Q�h�K�l=IU�������+W.�]�q���L��r�[Ta���e��5H�]h
:�2t�B�:��Sg8n���0����L�6"�J#�)"�!�7��m������t�VgS��?���mįkoF��Nq:�b`U� �P(y�����?��c⍀h�e����$��G-7�~Wb:�J{kA�;�1�'ZEHډJ(�9h����0���%M�x%i�$��M����Yo�'yW�D���Nz��j�G�ɳ��m�]yJbM��k*�8h ���k�9�9ɒɓ���g��]/�5M�vlq@�0/+tvfBT1U*��3SP��07_���i��T�2�+'�*�����'g�@��4|�D���HĹ�E��
�r�����}V�>ML�
�D���3b�HTO{�?5#��=a�=��ޜ~����kݼ�@7�@���z�1;Y�5�đ�t<�ζ�g�}vrj\k�d�?��?�ѽ�����;`�4�Jf ɺ��g�.��������]w.����Pus=�2	�W����/3ݻ�ZmZ^�ԝT
�5@�Ć�c�{_jqW=���C�:"tM�M�����ClW�JA�'#3�s��d���b��Y�x��I���j��k�x��=�\Q̋/��JO�c8gμ�S<�R�m��2'��8La˖-������b%�xF�N.��.�V�و��"JT��@]K/ן��Ygm�[)#U�6���^�T�.��/~q��-���E� �����t��.�(
чZ��I��?x�v�������ۭ7p.'������ߚ��jh=��+�}��"r�-�{�b7n&��a�Q���v��Q���P�ăsXK��}D���;�CʟtQ�J��'�|J��
zs��t��r�Jѡ.�s��aU�n ���n�{_W����[s�V@�$Z���|�3Z+�4��s��"Np�ȀVL*Z��ؔ8Ϻ�tX�Fu�e����z��K6oެ�4��Gy�����Y\�:Ԏ��"K�:;:���բ���{CF�9ې%&�0�F.�E?�����C#� ����HE
N��^}b��Z�u�Z���GSB��ۡ/��Ӻ�4[g���1� L�� ��x�~�o�~�(gicq=R�@\���M��L�����T�K�B��Y�Qܩ�_^ ��KOx����(�f%��x�iߟ��J����k�Pyz%FϏ��
F� r����'��7��׬Y��O~�����p� �er�^c愢�{��Ċy(E�~ #�*�FD/��xGy�╍��j<v��a�!ÿ�D�D����(�(��TO��B���k��d��7$���A��/���wg�C�xڣ�>z��7[��RoA��:\*�>Yd���f*��xm�D֡+a���8�|��#�:���L��Vm@���WW�=�ytt�����7��/�6-�l%�tk�y=S0j�Ƌ5�:_��#2N@6+�ʰ��hF2��ȱj�rY���g�UICؘ�*��L�#�y�j*%S p0U�@�Xm��b ɴ��Ҩ)�@�Q*
��x�Ʊ�@�}����XB[5���5|���Ύ���V�;,�ƥx���EB � �	T��646�a�T���Z��t2�E�O���X�@�û�Q��9����鐥���U1�[o����+_~��^x��Bє�Z�e0+�&����~��ާ߱�Ź�Y d�M�r�B��z(��n[��ٟ�����'�ॗ^���F�Tm�*����>�On۶��/"�FO�V"��\�z�$�޳�z�����tu�HƋ#�c^|�%Zam�d���m���_����3�<szvF렍fBs�%�����ћ!v��;����΋p�p�l���eG�@�%]tY��'���;ɖ�E{��s�t+`�PԦ�f�?3��)���M[d�C�ZO��4��n���u�xSĸO?���	S��l]�ҲQr覃�&��vh��- ����cp�����AG��йO���K����if("Zv�M�z67�0@�©#��[I�1�كY�VfvVG@�=�M�O����$Fɔu5HxKY�S��ꫯ���r
W���;N��Ν;��D�IH����4:c�hY4G�˨� �_;"�S*��E&����W��2����VA ���5ċFP%FY�c�U�fx������7<a�<��x�Й�\�Z�O`�<�"�v�1#�����V��3!_+u��j>�ʀu7Q?���o�~MD%
�����kqYcus˶�(i��DF�p�M���}HsS:��!�Ҍ�{� x鶚2<K H����D��W��a.n�ŦS��Àhc7�}"c�VW������hk�L�_8HI4z
>	6Ej6n�hm6��	������7jfՆt�(��ᘗ�G�;�}��_��4�9As*-K TZ������ȑ�"��V	u+�9x�(�j9Ţ�x�	r[��&�!zd�S��������F�j�ʟxp``�m}�5'̓.�
/�1o�����r�~�6��K���DI��.!�>18�����+.��C��l��L
�ks�Xb"�!�d�� r�$���L���&e�$�$�n�8�Y���M��e�E�~-%��YS��� ��8<�
�a�<�W=��9q�-F��Y!j	ǨĨx���;�n�1lV*�K�d�S����է�d�LN���f���Ĩ�3"����� �~f�G�E�J-EW�
 ��?��K��i�=�ߢ���ũp�~[
Y�H����GG4VI>���>SU�pG���ک�x}S�fAw���.x��a��ܜż�+x���"R
�Jd�����e^j`7�&K���6�044]��А.��)I2&$�@Q��H�5�r<�|�Y��.x�{�{�j����OG�d6�(�[�����yP��9�FH��gow��2�~��_���Pi�<@/L{�I=T���`��3x�
�$Y���O��믿���OĻ;ڻЀ?��o�l��p�p}�vAʁ�e�F���C�L��>��P�W\�Ai$�5/n�\�v2��)'��v����+�>�|H-qF����E�td���h̬��"7��z^��ڪJ���կ~e�o?I�o�r��8��N��J||vƶC�
D�v� �>�O4)#�I:xU/�u�3��O}�S����?��\�R7y�g�]�{�@���؋�;���yYpD�G��ٳG��mbb�#���l9H��NC�ؽ{�;_{�;J��d,��ts�*��{w\]&z&~
h�Pd4�Ԑ���K�[�lѡC�h^�v|&ʁ��@��i��c�����haɡ��s�d6�)�j�޽RL�MZ��Ν1��.�l�;��f����D��C���h'@��s#2F�҃4_ ��}mi4H��3b<���	���#_�/��A��+�2����)Ӭiϥq���v�k4��Gp Ԩ%"i	�Tt�Y�����ask��|̱9T�;���}��ԇėa���g�00x����Ed�g���a�קծy�hzh��lН��5-�/j1E�-�"����+��ki���5�6mz𡇴z4upc�<�!5%H�F5������ I=t�#鳲�t�ugQ�F����?�|z�'tm�a�`�G�	�bq +ɦ �qxA���@f�^��q4<���:)R%���/x�Q8�e�8v&�jҼJ��iR�:;"3�L?Lx����+8�lrBM1r)�$�x���-Y<_(�0���ǙQ>�C��r�*T-F6'�L��	��9�Xd:re2F�H����0�FnK�J?�����V�f�^�������	��qv1]�S#K��6C���p@��5Ua<��D�3)�C���q�!*f"�W�u��q
md˄D^ ���x
¯hM��3t ���}5;=~P��lJR�R�ӱe�������r'ʕj���F�H�3-e�R�+E�ޔϟ�r��Ç&��F��s���+�k)���w�ލl߾7��z5Ď�ÚKy��ZE�s��є�-^!����c�dq:��g�U���#
mUʵ��D���+��%���,���Nv�y�r`��Z�۬z?���+Ԣ��}�����?�m������w��c\+�l�r	61\�6�<��{���2&Zzp�~\5��o�ˎ�/�"n����;m���]]:�]�^z����p뭯'<AX�s��JR���zjѥf�GW�Q���eܪ��~TL/	~�)���W^��אNNБ�uæ��������0���g2�de���i����_�k��3��t̤���؛�]v�v\�Q�!嶎3R�<�J�495.mLwwO�ne5b�7����`I}�a�Pm@b�U)�� �c�RU"fj����-[�\���]1��������J4#��P�T:�Of�\t�ֳ��}zf������R�4�+�I��"�Ԑ���h�ݴ(�z�=s������^�G8~��T&����#��u���OO���Ȏ�[:z�f�z�-|?k�Ž��-�Wv.^��#��3Ϡ��^��J��y۶X�V6�oʢ��<�\L˵u빾ku�?m�X���椧o�f�CT/�JX��jյ�eMz���Z�\�U+	�}S�}�V��e[�/[��G,Tӷ%)��F�Qd RNR��6��܌oo�<�h�į�bi���kP�Ϣ\��5A1�Ҭ�5w�_�:�eVYk	��M���P!�󾓘�Zm�]Z=<�(1U�D?D�O�����>]s)�S�Y,�R�tGW��+�ㅲ��k��������:+�&
d��=����zy�K閖%�-�G�[���"s��-j}���I�8���Uݏ%�x�ّZ�Mg�&&'�����V�"ӢwY�Z\��7�M����K�O��5@Z
��*�i=�|��K�,�4��m1��;h�iw��������&k���t�f������?�������DfJ���>Kբ�(i�%P�R˭����J_?a����OsO���מ={뱞T����y���������d���qٙiK�5�i��g�_'���Vnh�H`=��;��?������E\|����+)[�l��؈��uuv?>X�N��m��s�(���S
��o�'�~�i�8�qv� ��"˷��ϷV��+Q5@qs�Tj$$��ʧ�^)Y%���nr�o�������d�u�='ݼz�T2���M5�)����\w�D�����IG/��/�3|av>����򩠆zR���6=\wҪ�z��w&��#)�)B�T����%]��U��H�[v���l����[��I�ѤP��!� }葄)|̺���L��1��kTXi5IG�H�E/%W�,±������"�����ik���g�=Q�<21�k1Ov�������TJ=�]��Xۜo)�W��;8m�Af�u�w7�7�?S�R��8O��0�9�|P�5�y*qc����#q��!�إ˖S)��:�8��K֒����4+�j-C�X^*�6@� �#��I�Q8��	�*�-��a$�*�b`rƴ��Hʁ+�@�a��r��M7����oSN&�p��IS���Mf���p�aQ��.O\���?D*�ƣߊuJdJ��nr��j�K3��b�dy��I��Uհq�i������_'�EϽ���[u�)g��/��"Q'�
�U���hve�*���'�{��A���7�.z�	.{��hD��Rɏ��GS��qj�۶m�ŉ4Z �$�I��W�Fڛ$�i������߃W2���!��r0��`�����"'��_w�uR�^y�=W�/�Pw���U���u�9�D�4�;��aCE��5��7��z^�'�R��0 �+�$!�aݙD5���y��Aƒ���C���M����Ozw?ݡP(���<x�~B	N�BqC)p��'˗/�a	R�V���G��X,�����?��Ĝ�I�9a:qww#Є��26K1}饗�k�6�� ;n-�F�Dr�ptqZq�iTzo�������Ǩ�y�*�MҎ͡Y�8Q��jedH�,y�@�Y��hW�b1��|����\�'�&R���v��"YY��k�vP�'��Ku��o���T���!���L��,��45��D��}i��~0}+jѐ�E�b�k)�'N�-�Ш�~A6�9r
_�r��nG�oܸQG���"?nɠ�Q��S���'�C�&v�%�V��ID�)ՁC��=R1>���:�BC����ọ&�-a`�3��iZ:"���<��u~@C�Vw&�d�+�2��9#i�=���ԃ�A|�q��n�i�K�Z�n��1�#G���K�M_��oTO���.dO�$���Έ3	-!��eBر���:�A^\��Ic/L$�UxU��l-��SߍHb���ɸ���8o܄�����g�p|"�����TqVb�ؔ�"����:�G:����f��YϷ�6W.g�T,��"�2��J �8o��T����N؁���o�O~�F�۸��� ��Z�^P
����+\�{�QBր��Hږ��[�#::�Zۚ���u[k|�*Ÿ� �P�O���6��Z&=�&�:3o	�=�;vC�Ivx���eKs���Gs�)/�J3��E:��Q ��.�`��G��b�&t=͏ბk�o����S��έN���8qB+C=m9�E�\�y�;����+����a���1��xS��A�ݻW�!�"'b�?��I���&j� 2�����q�2�w���Du�a�׮'���n�� ��p�e�i��A��-[��vGިTؖF(	�{�T:�K���X
:��H�B�֝#������%aIk��v�[�P��p�W@�iR���U<�I��4 15�R)L��F�II��.H>-�_ ]����ts-;R2q����X��	����8��{�$9��4,�����h��� [J�\�e`�s�ޘ���y�b__��$�P>R��f��I�]�vJ�[�j)l��,�Q�CZ-S5B�t������IH |��Α�-�z�[y�2N��d�{ۥ.TR�ጢ�(a��3e��tr*�4���(.L#7�ȣu,���o��2 �.]( ��I;��������w��":���d�PzH� �ςp�t=#N[Lr��F����v�ZF���l:���蜙�*��Ho(�^�"��`K0Btyuؒ�n+��%:�y�:Ъ��<���>NI:r<<�ފ+Q�/���_~��<����H��ј�C�Q�|ŢQE;� �M�ԟD�[Г�
�B9n�hj��0�o���K4a��dC�Š�Eo��`Z4-у>��-BҢ�!�!,f2�-��zsVI���?���:�@P8N�?X�dX�Zt2��8�ײYɠ�۷�t�M�ݬ��E�Q-��GE���q�J�c�E��R.�-8j�����'
�bҐEe-���(��ݼ�j���TCCt�ƪ1H���㩏-�J��5�DCJbkɮ��M&�f^���&a}M=��#u�$�,N�9�I�b�Uck$���FF��D���c�E}���!�c�5ZP5&�d�{s�Z-�Ί}���=RCl��4��b��X(��N��E@jf�G���E\�9�4�*�@DL��F/���O��+Jی;$MY�u(a�
��,c��0g]A��"�J�ZP:Z�V���%'P����f@e#�Cw�oR����/��P%)��0h	�u�֠bj����իGFF��i:���(��RJk�n�:� Mi��{�&{��g������֬ ���9�f�&Ѓ�hz���iHi�r�(�G��]L�R� �tx$(t��B
`λAi�X��E�w��eӋ�y��mz�b�V�Q�رC�H/�-��(O�4mX�R��{����㜆��:{|��惁�C�Փ��M��ڵuSjm��в�w$�Z���R��Vk3@U"���\q�Q���9sf���
O#ր���b-�(��f��bF�d�TY�KO?�Q-��ο��%���xnn�<ߔu�i�U޶c�N���E��W���k0`���[�G�K�BG�a<NnM��V䥻�_����R��)�zY����	p��}�;�#G�Հ��l~S�����	 ;M�'3��ѳ��4n��� ٩�gm9y� �>�Uz�#9H��N�.V��A��R���O�M�����W�b���LMk�t��%զ�1A4��U�*T~�@ՠ�Z:��[t�^�.$���=�M8P´�$�A%O�{㍃���o��������p�Vc�� ����v}+8����(�5��
25W��@Q���5��a�O�l��(��:�Y�Kţ�'���LB�u��P�I%7�Bѿ۶m�f���p�jd�)��8��O���h����8��ѣ��ﾫ�����Ĩ�V��,�1�0�-�2�t5�(Ur5_.:q�/ѓ��#�����/�Z긯ɸ�g9hZ�[$#�g&n\��������uK�-5Y+}�$We��k�aK	<E���T%-	���+q��e���{��~;�ղ>[�YG���b	q`���n��Z&1a��^��&���N�N1\Q��u.ԧa7��)Tr��h2cN�����dJ��7���#���<M��|�F�ń�.E�V�>3��W#�F���09391MO!Fi'�G��v9�sɲ�Z��B�chh���e�����s�&��cϾ������>R��1~��Ç[k�2��rI| �(d�㤡�a��
=�Yc���prrjѢ��'uU���j��\���8�W��b�z�+�I'�U�*A�H`����K�h�qq ��f�}B=XY�0�֞67M���N�X��P����c��Sv��U�$�e�;Л�  �2z#%XT�Xa����P�"uM+���c�v˖-Z���1��H�H߽���aP�qy���OT���v��r1p�h��C�0�v�<���`�5i>�|��u�TP@�\
�O����֨��δ	��om"S^�&E��ތAϴ�gP`K��_Doa@$���
�J����\� a�u�yO�.�F)��"FH{[[M�0Zۚ��yΕ�y�p��� �%I�4��~������`��!��P�V<@�n���h��Pu�����ի1��5�x�%�EpC"�O�B�Y�R�DN�:5O!���Aц(\�&��%� uE����D/�N�/���>!:	���q!��ȭ5�^�4��I|�<�^!�G�E�'!�����:���GY$-�V�a���īZ�����$g
V�B$���>Óiө��g����7��?~�>��
:�	��m���Bu���Y�R��N��=�W!vY�����%�2|�C2
*N���;!�5:]�G��n�0�j����<4<����˘!���%���2�kj6�O��Z=�sD{��_���m�G���z���']AOFW��*�Z58���؞*=����F�Y����7�4�#��7����H���#M|�:�'�4��<('��/�|hAv]�ȹ# �����Sո,7\�n���#·�m�{���	O!<���X��#P&����ql�L �K�XgW�aHKifk�"����Udk�)�fR鑱�l�l�~�r�[6%2]o�d^4S+���H���,9	��͋0j�K��.�N:t(��D�6�y�#�eE��:��(�l�<m��#��1�1[�I>o��7�Y�i�$�Լ�������NyGN��+W�%KC�w~v.����k�A��`��_P4���,J�g\ #`(��ʒ�a�5HRn5A�⤚����k���$3�����muV5����k.���0�Y])�N=�F�0�=MN�2�VԯyrRfʛ�s�zT��%�aI�h����G�#���htO:9�I�~�zil����8&�Ih��y����ի'z�[�X^�G _�E3T��~�(�����FہVy�.?A�CI�94�E��k^�'��<|��M��nі��p�+�:kj�V�t~d��|�	V)ݦu�ɱqԾy�������ܒ�����9�o\ �(�&���ś!�q^-�k�]�F5Y ��)�,c�x�-��Q�H _��"zl8��Ü71�8`g�Y�^^��#À����p���b�Ak���QJ����C:�W0�(�A<�@�h�]t�>g� Q,ZH�ͪ9A��$T�s�����=��<�}�?ʾk+�@�4*����Q:��p�I�蠼��yw:J�򢣓w��4Ҥ���p	hr~Q��h�a�k��1KPˬ�����kH��ڡG�KVI��{�%��Gs���C��$S�*D�2���==]�ã��κukéZ��2��l�k������7���.���>ӝ���fNH!�D�Ye,��D�m�Z[�V׿�k9T�����Ֆ��*�L2(s3IH!	!�Mr���3��󾟳wN����x�������}�wz���_UMŜ�{j�(~38ޑ�hӨ.��!Q�A����rl Q�N�D�%�,s:$�$_L��̹Ʀ��~�w���G>��M�TK�2��M������B�>����k�4�&�ᄈO��u☠�>
���2Qoj�u�֮]+|V��f�:˵�z��98��dʳH��X���y�̀�8��-��ŕ�܈1�VCw!�25��c��Ʉ�8�(�z�h3k�� ���b �$�����ş�l���x�&L�"
K��T)՚V�d	K�_C��A z`~��#g3$z����Bu�Myo=��p�Lkv��r��y^̯I�o���a�R1LcM�M�HmX��ب�
%쫯�r��`���>�$B��2��p�b�b��;!:V��z�4�gD����H�N�"Kc��I�{K�I ������>K���a��VC0f�^�%b����<�t;���������0̀'�ᨓXGKIVң���H���.8R�2��f ,��A�k*Q��55�B<N�<��P��<, 14�RZZlM����_����.H'%�s��|-�w�)Ɲ�l$�	V���D1}RN�Ҍ�ȅ++I���A�$���ܭ�4�*y'G��{��qbQ�+��&�o��Bb�^�=f;p�[�|5�\�BU�K!>pc�K��@Xx�P�Ӣ�G�'��Q�/p���g64x�K��@��{�h�Sҿ�oh�hm+L�������'�c�[�I��ݴi�M�H�'��4Tͼ���_�(Z�W���p��|��wN=�T��(r�����l��l�!����/��0��Qq��陪������$$0H���R��ɘ5u�^��e�c8FD��ӆw�ׯ�h}�Ө��ّ��r$�Y��}��� h��H���/}؈a��*�$a�c=ñ��S�i�+V� +����q BU=���N�0EHywv
�{i�V�FX��c}�W����U~R'zF�tȷ����!���?�%:,"���j_l3�6?�D�^���#��ɽ��m/3��{��y�gvww]y�7�t��͛5$e��oJQ��F�Ī��Q]��u���7qb�/	�~W��Z�Ę��a�o^"p8㝊_����j(	���߾;����/ǻ/	���&!��p�c��-j|�W]u�SO=u�-��4�@ޱ��j����/ڱwR�v�	���>�Y�`nذ�$>� h��8C��CL��B�{�������&�Ep��*�#��3xy@�v�q��`\X*�X6i��N</�LA]�~�esvP`�A8��55��U��LT�&(6	�&�s�g#qd9q�%h�?YNą��E��H�z}:giR�kt�lݓ-�����[�N�:���l:���26l �β/�;x���4�{����c��R�|X#����h��c�II���]�G�<cjf�-�>p�A�I=N�D���b�)4\28�r�ьׁ�$qgp8�����@ɀw�C`I
�+x������
y� �E��.C�A�*@��MI1�1�{@g�ʕ�������R���V�z*�p/a֧��W3@c��u)�w$���^z�b1�c���w���
D!| +<yXt�޽{�XGN�3��Ư	�=���
���SX��М�("!i˖-�:�P�AR�|]�ȑ����
��x
xE]�G~[`�ū�G� ���� �.��.J�Yo
�=`QЊ�1�g�s��
4fxS@�j�ሓ�#͛n�h�L陪+�ұ1g�V�����#Ϛ�<����&��=8�C�.�-*�but������ZJ��E;��^�M���2#�PaA����.BQ�A_��$�ER|��#��Ud�#ڐ[N�h����h����5��fr䫞����1D�N����r��P��45u�W��s��2�4B�E��r���)�9��H���B&�v<���⬡�	�����f�֐ �� ����+{�c1Er1�~D=>�[R��O%J��C�[zv�,��^��H�x�E���]�Z�I�$��"�i�*�Ѡ�K��Fq����*w�'�A/�ίu	��/{�'�b�Gq�l9��Z?���^��?o�\]��
s��@�?P���
��STW���ٖ��*�8��>c	�ar^o���%���xR1i�-W���À	M�E���g�}V2�.��ˈGE�M{G��;�@�
-�gǚR���?|�w���J���1���X����*N�U�'u����/�p��=$i�	�!���^�ޜ�H[�>:٘9YWո�#�� N�a�H�RxȚ������!��$ʃ�mlB��V��⼀�#	�.�i�2�Օ&��T\�_L'�����]�Դ��l�[��H�~ȡ�ơֈ�"�\�O��Z�� ����)Lg��-Z�:]m�U�M��j��d�
Ł'�I�pD���m�H�˫hl�a��0mZoww����2����޴K2^��	%[u�%���n��j\���ېs�J0h5v�4�+{KG�R$��x5��2�hIO�&p�V�U�]5)�YuM�> ёv�5,�]��`���`
����n|��,"1����`=W��S��c�}�(4'�s7h�1��@:�8�P-�9k$��?<1� կ�>�Oϻn�:]�TD�B8�3�.za�"d�k*HE'eG?覚�9ɸ�nN#׍�M�F^�8���\x��ХJ͔��\�S�$E�	*5-�Ɖ+.I��'���t�+ht��7Jg�I�IHLr^�y$��B�=�W��G!������3�S�Ijjh<}�i��C=����%9mj��-�t\Fǌ�m���ޔ��Ёr�4o�l��1E4�ԻH����"���Hu��;_q�C�b��j`4  ��1��IH����?���5`�%���_�"�(K�܁���������Z>��x�O%Mv`/V!���N�s��M��k$��F�p�l�p����zbS+�)B
��$h� y���>W�D�Z�[��7<�أ: �E����y���H�0E����5B���p ǉ6������5Z*3�I
H�G&ҍ��,ӴH
����t�k���1SS���hf~�h"�bU]Dr�s
\&;��K�q�4պ�Q��i�K9�I-��)�+d��d��o��5�!�J_��k�(�1�E��^W+-M�Uw�$�w�+j�IQ%q�
<j��>$�]a���$��	C�������-��?%^����5� �d	��21E�Q%a�
�u/��;��>��]��XV���S�R��h�X �����{��_[�n��@ =qg&�yݿQ��5�[��JO�?_xZ��c�^KҪW�y�i?�xn�t�d�>���_�Tf���X5�p�8��	��*N�İ�d�sq����j�r܍�e�_��C*:o6&�e�lܫ��ӠPuQ&3�V�vuu���Ǵ)&j�����a��\����Кy8�O�Mҩlm��|i۩RNN�%Vm��am�l�9���jCKcm~rAZ#�M##	��jb�!��±A����0X�p��&�d�hh7KZָ�=6����r�$�p�PFD�>�sx�0.�-&p�� D2�5$m}��u�����E�H4!�ǧ�]�0��Rl��W� ���g�� ����$z�7R/��1�I�!^ψM`Wm�U���z
�J��D��"������H<=�;� ΁E�A5nY���I��*�GH�������w-[�L��H���+�iwo�n���@X-�$R�7�*�"����U^u?���0G�9}��Or� �	d�C��@�lhHB"�F�A�b$%��9�WKy�0�F�}J� _4y�%X�� �&�P�H����9���s�_S���)��6l���HM5<I�H�l���C#�U���� h�I�$����z����QZH���!Q<\.��Nc#�b��7o��ZM�Y�-<��!&sƌd�ԡ���Ds@��x���6[��F�^Hl��x
��ռ6��W��֬Y�WL{FAz�<E�EzMj@�d]��������!i;�bzm2�E����<9&�"A@36�T�D�h]�E]�S���+ku`�Ф%MN�1}��$���� �#�>�6��ٖ�f�;VS�G;e���E�����Ƅ�htG#�z��[�j���l�3�$���"w���}}G��1�������k��!�`��oh�y��Edj&�)������e���"���K�&��5Sb��dxIΛE*�����i�;ᓉ_
,��c�Nc^��2!��d9>�=��LD�-����
e,ih����-ॶ�~����o؈����{�����w�#8r�9˙p|c��Ey,QL�"���[X�C����9�ΆcE��N�������^h�LS
Jy��ì8��~�9�	�Z�f�#�#M�)��N{QL<ʱ����ܗ�'�y)k�Kq{n�%�/u��#���Ɠ�G�m켏ZU*��.��I��ho�ی��ڟ�B�);~Y3��  �2��8��J*sr�y�.�����0*��U?�~#���c̼�η����:��;��M���e]�V&&#��'�L#���]�-A�Sp�'��o�~+��f͜)Y&�n�0a5�Ւ��_7��0����G����N[���^����3!Ry��@��d:�(v�U�� �q���òI�S���8�)$]A����"�ܚOB���[P��M�ch��^ZO�!�$pt�z	�'���y�/��S����2�h��W��2JGI<� �����
���<�����_���7�QQ�G�$�]k
1�ބ ��c]��2|r�>�F�x�)�P���lEh�ϊ�"��R-h�4|�V���q���Z�����^9z�������Hטkشi�����*�,t�#���T���[����u��ΣGg�o���J�=�KK�$�k�؇yo��Ж�w��tM�O�ʆ��#�I}[Rlj�A�H��q;�D&SO�U�'�c�|#�4���N�����P�A\ue%,�ъ������	߿�+�۝v�il!�f��{b��L�'���`��M�	Ŕ�q^�
�<���N��퍖¹K^?�c�X�a���q� !�1����䨽�D�����Է>k4��0o�\똙��Զ�jܚCG5�����N;P�X6[��+���C��s��aPu�t��u}]˧�1�=�
�y+����ӵä0��i
�6*�����Sg���S���x��$/���l CuN���oT���;q�҃��6�dT�f�x��t���X 4�&1�v�fFV��nP��T�=1b<p�Ԥw��>f�_,�饗������0���=ڱǬj�x��(Ggꩧ���$�(sMZ��?B*N�bu�q�t��� "V%����b�"�l�'9�8Ғd/̡d	0��ø�d�y�������a%�����`kE�Qܲ)����D`P�3�G^Ι��6����2�_+F�S[�݁����yƌ^2F�==��F�k}ƪ4H�(���m�瑟�������[��-a�0Le�(�Je�}\��/�A5������^��:�XV���;i����R���`RĜm�zΙ3;�d� ��J��-�S�j����s��Q!���Z���	�
�,:e��U�ԑ_��7z!���|��g�������l""����� I
c:,'��-���M&�M��{��F'�\�F7i��9 (�$FjJ�R�]H
���)ѷ��_��n*Jk�t�RJDI��/�󆉯�Ӯ��
�u/�8r��&ëx@n��,��'�l�)E�S�J�<���	�)Xsꩧ��AS �0��`ĥ�`��%&3�J�2���U�d�D�WD��b_� 4�9f��8ٮa��U�ؤ&��;�H����M�uwp-/*�z���w�'ղ'a��(L���aDɉq�ZM�sR�ը�h]@��ȹ�K����DJ8�<��UG�%�<�q}��@��VE��b�qJ�p#�ʐ���|��;�@bkun�y���,��'��D�]SSAH�D�	���pp�N����8����+�#�ci��U�-�t~5{�z"Z3� BR����B�${��-�@� um���
:�"��V�̋���1Ź���5mc�[�첡������tG%�$9���ۄk	r�	q�Q��d���{O�>��?|�U������5�L��N�Gf�19s�`��.�*��h�<g���%���gv⽎g�}C?YX�s�wX�z�2���%X�P�3��:�/����^wg7֚��y��.����l�%<'�����'��>�T�=�?�Ru�̭�l͚5�W�^�p!&���g��uf*f��L�z<�ў$(xN-��<�Y�����F�2YIB��8��� ?r����R�#zq��x�mįK��K];*�`(���Y��6Q���ZʢP�D�#�ln�L%I����(��c�}+H�X�'P��C�<H:��l&[�k�Y��5����ć�?��<����,�U��y�k*ȰHf�8�ӦM�xe#�gG<�@lD���y���Y���t������0!s"8���i��8�L�{�\ʗJvB����Nv�D<�v����B�n�hx�3�\���mu��&:p������1��&>R�G!�+"��1n&K�cy�&u�vL��
3-Ͷ���d^zh�`W�k��d~�hĻ��7oތo O�.�a���F/x� 4%o�L�RЍ���r��-[��G��a���lp�q�?D�F��+��U�{�1�	�e���EV�X��i��9&��;^qrõR�/֣i���wH���8lt)֚�z�&�����Z|i�
�CpD�/A}DТ�^��m�g��h����p�wtU�q@�)B�5�����;��hCW��ø*�X3��ӗ/_NMI�n��֖��Q�װy�/ș$;�c�Y" �g��K'�0tF2���>�x�}tD���u�VVA�ύ�" �(�$�!JV�g|���>�1k55$\SP��xӭ�qk�[�"U�<�z�B]S'^q�X]Dׄ�CC�.[v)����c���D ����XV=g( i>�T/8�d�(	��LxL�`.�M�`^=h�1l�~ȃvhҎ�@�ƛDHY�'�/e��%2�@/9Q�fZ�Ojd��˫f��IO���A�J%�����>	��
�����cd�J^[
�4��Gq���h��pdj̺>����|(�% ���6-�����K/������vD�u���Tܗ���W��@5FA�?Tc�HՑ�V�*7�!�7����GW����} �ӀQ��ߴ,qC��\ScX�p�j���`wjXoϴ)�]�V�9���W�X��k�y��'Ib|�����d����cAI�]��SO}��H�,����Z�
������� J7$���D�.�%�c<dA�bO1����r&3��U*�[[��~����r������$+�?����}�j\\W�'fC׍�b`�Qfb���$���F��cﵭ~S�Z:M��c��֭���AR�ƊSߛ�2d��T��J�����3����l�-���dpTJO��+H�̘�mB� ��@�!c�/4ʮ�D���5�g��$BV��Xă���:��8��eo�P(�O�l!�*�#	���"�bnxO@ژ`���",���k����cؑ�ŃB����ʒ%Kv���^��T2�4�W&�X�k9U�I��c��l�;C3�X��T��V��Zi;a��3�i��!${l���6j��Ν�ׯ_O�Ϩ�����i��9�]M�ճHv�A��I�Ɩv.x����,�4 
K����P)>��E��������L�hƴ��-[F�D�BnB�����aC�nИ���'皔bRM&�) $���5o��SN9��}X���/�K�q�� ��NK��w�LZ�������s�������z�[��ni?'�Z\!$]Y����`G��cE��#�n6X�7��_`4�eU�SS�Lڸq�n-��&��L��ڴDH��څ�u N
I=`?�*6���d��M�+p�	�*1o��fY�*�%�J��mDZ��Q-q�C�Uϛ$�)#B��\<�n5Z����g�,yOL�}i/�$5��>��1���_�==��w�P�+nm=��?*gNA*jq��%%[�L�[�����c��DCۆ"L�Z�Θ���G�z��O}�zYi�3nm#�дfP�+(9�#M)tЕ�{�y�LD���k�TiE�5!��Cu|��b<��&�#�����e�f�9�@7�P��<�-��P���3�;�G}�iR��W�F��O|6���sw�uq�zZr��x����jo�:���|�� $����<$ݘ͑�	m�&����)���s^�=L,1���4�L�_~����.�bJ����x�L��U�fn���q	��K�r�)Ď��
&3Ao@�	ᇠ��hĢ��	�&��'��r�<��DM�/�^ø�fy�u�p�������2�l�R9Ac�O����|&�� Lh�}�-ġ@q�x���塄^��*�k¬t̋AJ���8��w$��S��u,Nϱ �m�i�q�I3������p'�rт��rvB��E�f�OX+� �^i��;q�s@�4�	������'�#95����A|	}�6oޚ�T�:��X�hL]nz�w�T86.�a��@��k���@��8�DF��;���tX�7/@!p.G�	ۚ�Ύn��8���v,I1��p4gb��=x=8��A8�c�i��Շ�z�d$���nA碆��Q��$1�a���p�j�� �W\��<�����.�x#8T�u 3�IKF� �8�Z]\ZP$�4'�� I�v�Ҁ5�Bɽ��EА�xO�<�,wafe�mC��q�P[�7!%�M��-]�$;F����Ј;w��x(|����Λ3w��9z�*�>ٍ�s;�	�kT��o߮��a�E�`�d�l"W]Z���\%��r��J5�׃��tף���?�<Eͧ�z�;��N�Q+�-�K1��4x�+��ر[F'��^�AK�����(I�Azv�H9�$s��I��)n�L�\b����v�3l�4�g� � K�S�M�CW^��dIE��7|�;����?�-�oEϥq�Fz̍7SW��J�t�ȵ�4Q�2ś�Im����9M�u�;�sժUD۵Q?��h�4R<v)�x �c a_�z�w�e�{�l�;����Z]D�*�T�u����h�� h8t���1Ʌ��&�x�($sKO*q	)�/	�b��0L�2�AD�SSDd��6N1q(�d,	@A 6��%��)AЛz��������D�ұS�_p�g+t�c�1H%9OQ�ja?��Eq�Y*�!=��c�(�o��:�9i��$or;4�~*�#dcK9�G�.)M5s.[C�Zm ��_���8h���㘈�{n���U4���̕ѕ$�'��lp���C���� �7���[����''��LP|�5�jI2�(�قf�G��q~[-s�ZG�R?N� `9�r�q_F$�h�j��N�S�1P�O��db G�w��5�Ĭd<o*�q����
����BR0��եK�I��M5�
y��X'�\)��	E�f]7�������5XV��~�F�4s���'��0�`�X�ڲu�VM:N#��ؗ���9���t�52! Ɍ����K9�5]X�hWi���\ҽuq��H��>��XƴNj*�}�"U|E���/���g�[���y���5��u�Z��@�-^��1�@�ewu�u�Y:?�t�gd�`����Z^��;�,W@=�<#-�݆��6T::�Ǻ#{E�~ǎ�.�^Y�l��Hj[z��ź�;���(PY�-��?	��&#�L�I�E����v�6��~}&6��fo)#5�CLK������:� �����w�������pC��:����-2A�����ׯ]�6)���ȣ�@�VF^�����3�<Cl�
=��w��I�p�pJm�*ӟ��H_�������T��G#0t��g,��g%�hѢEH(A"D��5Z��ƣ���{��%�N�:�'y�����U�z���_��M7�t�]w��[�p�F��\|�ł�Zn-��7b�^�P�V��g?�߾6�dĵ������/�]�z����P���MP�}���e%�QXG�ŵ:IxK�W�uE0Q�<��s���=gΌW_�K��[��Nأ�z޶m�c�=��ɲ���>��x��SOI$;��}�=�	`2��u��i��gi@�A�}��?��w��]KX,�nJi�?�OPL"�`��!�K�ad��=���nD��H+�@�G���
*<g��_�:�q����초C#B�fK��C�TN��%~�{[�r���$[Y�V�x�HE�e�)M[%&y������зM��`�fzQQ�-�$������[�PR��[/��Ng'��}-!?�<�jM���+1�`���@ƯaL1Z�H�!���M'���j��	M��K&nf3�7J�[������ծ�?z���?4��}�,4�И����TH�s^Kn[K�sZXӈ�s���Rp����׿��j�Z�+gP+(!��O�L�+:8���Ÿ��{���H(�A��-�BL�JQ�,�!�}����x��11���,���B� �� ��\'�ɻa9�s��_�vH:(c�Z���Рy3�B�c��<@P�����1H�Ւ�	e���I�6�wA�8,���FGG,�8a<�c��FUb&zgr�ן"���al�ش�ү�ϙ��,�XM@��QД+�tG��!Ǿ���Tu�4��F��-�m#��������t�0T���z6jzu�ٳ��,πh||�0Y�f�J��,I���Y gp����Z�_|��_�Yk�-�W�, ���$	B^����Ǒ�V����首&�h��ǵ/�L���g�Y�f $^�*H ��z�w��������>262�a��o�,��$�B�r�1sD�-�{-��ul�k�������~K+�XȬg�A�LC&�M:|��K]V���h�9��mS�W����F���@j���r�Ei+HRs�H����I�a�����������Q���'������_���{�ճK9�޽[��mo{h��O�W��5\���Ӈ�'�,�9�v�!�믿^x��p�<؁�a��_�������ɟhQV�^]�
������9��eΟ��p�=�P��9�������?����e�]�9��c��ek��|q�����T�h�e�c��x�G+W��r%q�С�����M�:$���e��\3�4���<8��[�H9�r�Y����5(ܘkj1�3|�6�=)c$*��	���411���k5���W�6�i	��n�MR��_*���q��u�H��׾�R��6��m�s��O�S�3���G�w�L?���o��)С@D��-�ZÀ*ܩ����dX��n
��	:&�ʕ��	Y5�����Gƍ����EJ_߳�������_ዺ�E���w��w��Ӗ/_>p����)�F���}�P�5\����mj�JM�҅�dj�N�<�����0���d�Z���gR��[n�v7Y�lv�	خ��#G�J��1���e���H��F����W��7�2���a���@L�g*���L�FULl �H�zuj�V�7g��x_(?�̞Ml����p���3f�L�R�1��ksO�6�;�&&�Y�5ZQ{g���8�(����5.�ٳu��y�My�\4>{�Ҏ�۹�m}�bK��R����{�ҥ���{�G��Τ�U��_1�����گHvW�%�QD)g���@�TR��B����B�qU�~�q%A��J���%�3S�w`8�3�d�m�r5�ώG�'R����!�'�:p�T��e9�G.���^�$���s݆�ͭ��r���hS�@�TT,�&'�b<��srű�{/{����!���l.�t&_̧I�z#o��Lߴ�>>�Dxz�P���w���mECbo�o�3�ɦ�δ��&~��p����j������#��OȽ���GL��˨-��Ɔ@[�Xnmh��(X�c���"�R9�3/���l��]�h��[���|X�B��:ڻ�[����۶�8j�}"Ҭ���J�tuu�{�,�S����CC#mm�o�5uw�S6ci	�RU?L&����b�=���j������]�M�X.k��S�\:?:��D��!��B�(��l����9�X�,G��\�.9>3��iA"��Z�
��ٳ=0|�2�J%
ܤ(C*ͮ՞;�/�4kB .I7=$~o��V�m�_f ��A��׵����Hg�x�T��!�2A�����b����b�F;tx���2Pu�z"����|�3���J)�׆���/�N
��+�<묳d��ֈ3*dГ�mf�{V��p7e�IF�T�NJ��m��Ԓԕ�_�n������t��[I�'�mC�_�l�dh�+uĳ�4	�%���䐲2=�� �+)��SO�x����	\=�����:x���Hϫ��
���+�z+e�U4�Ծ���h�"����Ǵ�HJ��X��n�J���W��W���+VP�f��V�-�kX_
�ƿ�}�{�{�x꥾%���"y�tiL�G7��&�t��ҾP��qD$�d)�B���o��u#�N��я~T����zQ����$ J���L�8�?���zM�v�
��rt�ث��|饗p�Iz
k�W�ZE���w��@��q�J��
��á����=��#9������^�J	K�j'�]y�u�9�;��&đ'򳈸I��㨩�E)�B¢1��e<y�y� ̭��h2���ѱ�6��)�m�!�FF��K��p�ğ��m����I����YΜ9��*�pHe�U-;U��3p��A�v2����*VPሿ*^�-�2pZG�S�J�F�"����I���zNs
��I�Rb�]CFH
��%:�7u#�:ȇ��*3�ߗB���c�� y4�ZV6����� �t@3��jk��ظq��o��Ҳ�N��\7������o%?5 ��)������u`�Z��Z,��֚3投Z�*���0�c��S%�ҥ1����A]3:.��K�J�}�&-�|������w�d�p�K<'����R1�PG�֚3���pYa�<��W_��-�ݤ�XF�E	�ZZ�!!-2����W\�0>]�����S����IS�|�gN?�T���hc+li�*r�3Jd���D؊]gn�t�;�o1�iS��Җ��B�M����ˎ/L!�_H�:�K�cJ����jj�s�9����ev6���Xl�C��Ji�.�E�\1J����.�[�H_hb��۵>����\��1�.d�.:�����=%c��������1��i�.�Ց�J�a�T�:�CY��x�c!y3��m�T��4:�CY�0	�: }���8���\SkK;I�BPHT����ÂFì�s���O�<�%J��&eM�e�PL�|W� ��ո�	���tvv��%5P����x�|�I�G��31/��+hN}u�.}Q�O"������hln�<��Ȳ� ������fT[���A�<8��o۲e�޽z��[o���'
׼.B^�ɩN��rjwjJ����Þ�jM�W%)�4��_M#���B��L�w�4�wG�k�� ��F><1!�N�#i� }.Eҵ?�p�`B�
j�7�d;5:���r6+�x�����*B_g���u�������xwg�j_|q�s���7E#�c�1C���۹�k۲ҊʤCP3��\�4ҳ���
���6Yw�y����+V\v�e	}즄04!��}��T<g��%�Xׄ�6����V4PBދ�]h��#ʹ[�k׮ݴiY�Q�f�g��/��oF[ߡ_��;���������[�m�5�m>��s�N�&74�4[��L,m8�[��T�jz�����@�7�
��L��ȠhCS��7{POirtLfv�&�!�5�v�ls��+�;w�Z�tI[g��E��Ca�X������ז�g.\�ן��'-jj�����[�֭��MW���z͞=]R�=j�x�����	:99�g�=��ۃ_����B
?q1����dA�y<w��Y�59�A��Fx������^�W�GV9~�ޡ�r�{
i�6�87��
��OOL�����vt�5~���ÒB�ӧO%�Nt��w��/n�ӯa��|����R�&���^�l�Px�T*a*�J#��Z��s��H�j}(	�����j���0����*�#�[*x�)���"�/�T!���Wr�z�Y�M��j|W୴�&h�����^w�y祼����c�T� 0ECK^x�7�(�c�1����� � �SU�0�����=�yό�9뉒F��=�YG��HRL��mY�F��Q6:<"�w�o�]�F��C�tGɴ�|�+�&��MR��)�"�u�v����Ν;�c���P���:I�R�S����ho��K�W?-�C��A��g�J5�)j/$��~���{�����93=�=��I'JmMF�R"��N`q��+j�n�|���j9ah	ߓn��e�Ԏ.��mWW˩L�� �S�A��ݛC��nS�n������l��ɬ	�I���:��ӓ\HpbR��a�4OE���cz��8�"�_�&��y�8�P ��� =Dl��׹R:qSc�/^�5�������"�飏>*d�+æFړn7�$� Q,%H���cN�2Z��fbq��V�t+��@�.�dr�1.�࣊�z}F8C�&���8�[�K�PV�������wEȵ��3f@u!������$�Yz/�cH�2�5��{�M;r�pƏ
Y�0ؑ�R�f8� �Zb�^~���}�{/�[�u��q�t=�=��+�e��}S�4�ܾm�O~��]G�f�z��޲e�q48f�59�W3Ij�.�ݢ��I�����5�H9�Q�4�3�<�fY O�7��t�#�<"5��L�x%ql,[vk�� �N߅�B^�X�ݰa���%�\BG,zM��c��\��-� ��	�B��d��8�1���%��ȝ�P�h)�'�M�֯��{^{�[��]���b��FF&P$ n���2�����ɺ�fO���7l4:J�N�2a÷\�R-��
}�P�󂷚QA���׊g�� C	�&m(��(h$��:1�[w�2�!1���;���tɗ:���$x��ׯו�d�O���҃KR�	���� ��8r��Y������~c˱�ԓ�۶ms���M1�4/���O��Mi�F�_�OM��p�:h�O(���������ݧ1�Y�Fʾ�%�O��M��*I·�����9��ե�t�T-���ZO��&;��1��x;�ٳ�5��#�Z��o}�S��������� �#�Z��"�z2&If��e�b5͙�ܕ>���S#U�@f�)�"�H*��BD��vr@흰�A�G�#}pƔ�	�K�>Q���8�Np�U�F�$]�ח6n�T����d�QV�H����|��z2j���6X�|��ի-��[��#��u,!'����xT�?>�k����f��u�Y�SN��� mxƦXe�٢<��W󲛮���<��:F���n���H׹Ӧ���s�������ď��
<���#Q,��Y�#M����_x�_��z\ L�dO©��L-�����o�]��;w���}�l�0J8Z*f�)�&�I8�Xz���0�d�Tc
z�@䀒t�j�D���xs-��c��ױ��~q3�����*P08P�g�@�$��g�3酴��-���CG�JtҢQ*���f[FF�h{W3�∵�VQ+��E��\VNN���C�Y2�8s�iT��{�־��2�6My���t�UpZ�Y�gC��Y��۫/���<�L�x(�N��G�fc؅;�A`� �9�������#���w�����u����ҋK�,a�� ��)������/~��k�8C�r����w�.y"��ĳ�:]g,"z]�A���.��t���G��C�Z��р��tk� 0t4��V������ %MZ^:�����E��`�h�8�&�Pu���.�0H�QG(P��fY;s�Ў�{�"�O�d��Fq���W�Ǎ�ˤ8cx�	����� 4�Z2��j�^{m��q���.�TB�׈C��T�bc�EgIR�Izj��8��<m�B˭G�$T�������M;f���C�a&�p�PT�������/E������(E��Ԯ�W��7v�.[Z���`=� #�6	c\l�!V&�����Y�4�ʛ����Ե��"1�U�.7�f��r�J)uD��	%���h�V�⁡A��==tĚ�M��<��˗�Е��孙�!]�=pp_5*�����<����)S��[R�=��z{uL�ٳ�65	�Pʣ3���X�t��X��t͏N?kՄ�_|�E� a;�� m�s�?US�4K�4frY
�tS���)l��/8����îN�
<��3i��iӺ�{n��~���k�
�� ǮC�xM���.+�u�wj?���}�#��ޡ��Q�  5ȟ)uB�Z�b�[��KW]u��?��o��:���������?
y}^vi�&���t�aͤ���љ?�JBK�W��g�2�
{�j5�a\^Дm�2p��QL�dZ8HpTS_�e߇u�	PK^����ʁ�j�V�Z�䓗�u�YZw����T�m���}C0޲�w��|����a�$���J�����_#Q����f�8;w��w��'O�I��ȏ��r1osP�������Z���H�Z��R�>��_��۪#�C7w�<�h%��ZM ;�Y�2Z�j��_\;Ȣ�]0$/��(d3�ew�}�$�dтtqX��H`���>*qA����[n������ ��1l6sc��B��� �d6k͛� �:�V��k�j�7W���榜��T'��[��>K�
��f�'���2����@�^��%�#���
L��
4J�V��lP�%Y�q�Ke>y`�`~q6`0�Џ���#v'
��7�?)'FjH=;MZ������Ôyj�5��o�Y���`�o0\�h���>/�a}���<��C�,:E����>2	0x4�^�u��:�I���D���K4�ѨD�d��}�Q/�cl�LM^>I���y��IbJ\p���:�p�
"w�^/{/�$W�(��wMtX�r�W�����*���i+D�^F��=�`�w7l؀�!Rs��O�I#����q/�+:'w�u�Ԇ1�����a����=N$�248��#C�]�z�9X �x�0s�v^����M/����ѱ3&�+HkB�E������H�
�5:P#�G���%� ��YՄ �h��ah9N>�d)x�`�Ɗ+�/���^���ڵ�Իǽ�MN�$Ԟ��_e9��y�{dvOm�m�J⿡� 
���ɭ[�iT����z��G1 �_b�aj25�������PT>j���K�#o.�Lg�p�謹�����:pg'@HX�B�AD�� -�;Y �=���I+q8{U�=��Sͫ],n߾����2I��ti��)�:f���ۉ����/0����!��&����˖-�s���=N�u����y�t�M�6iH7n�zO[ˀ	Mr�)pl�Q8��S΂o��Ib4�A��&sצ��"_������g��ΰWd�d�������$��駧رc�����{�ǒ ��IsA)2t0.O�)�)�ַ��-*t�p�t�8��T;�¡>)	�A����u��K�X�"w?��h?��O1�p��F��Lj�/�~���;�5$=.х��e �.�x\��>9���jJP���P��L�0)�
'e�|����K&���_����ia�'Q��Yh�W�^-�x���FQ��eQ'|0��m|Q��j7�����Y�F3k�zϞ�m��&����&�o�:J�+!���l�D�Ri��,� �hGsS#;P�a�s��~)�z��+�z�'e5��q�8�a+�5>I}��m�R�;v�x�B~�$��%]�V�.Y�p��+��㎋.�H2�&�|���q�z��w�fc�7�ɬ"��et�DH�� 20��-n&B��u�i�:=�����3	��z�	�	'��UC6��D���HW҆��|}Lg@� .�$Fޥ�|2R�])���	r&n:'�7�u�}��{ ���r��믿�����L�0�>wn-8�/���o��+�q�`�m��
-��#H�̞9������@`g��)�7@�:.�nƏ/��/d"SJ�}4�	4I0�?��i~�\��.����w/���}�C�'�Lb4H�C�@P\�Cک��W]u��;cs)R��4��W�ҡՇ���H�;��ڒ�Ԣ��S�J�����Oy�'j@����E��y�C�SP�ꫯ惣�����N�8���|�"��O��cl�$���k�5�����fĻ�Sw��_ݢ'�cj�6l�|�5�o��g�}Vtr�!�]��	���|CcNJ�ŋ���ZTJu�ٲ��ϻw�:k��.x���@�P�����4��ISݺu��[q����&ׇ��$�n�:}���ٚ5k4�)���$5�N�C�X����s��9�EsSsk�1��m�5�GHQ"�z���>�=��ٳ{�iҮ�nj�/���]8E�h�=ny��s�Ӿ�R:�fɩb[;;���a����3g����|�	=�~���'���~�X,lݺ,H���3�:묩==�����R�:q��Ɯ��h5�/_��f��{��jl:�[��,�O6��B�p�ʳ�/^@K1m�C}$|!UFtJR�u�kx�F����~��{����V������Q��+�����;�!�֖.]���'鹉�_ EG�.U�`�ûA�r��"��K�=��]*��=Q�#k�BO-`d,6^�	q��w���-A�Zbr@l;?/\$�2^�Y��U�eAϏ}�c�����TkZ��p,�h��������0�f�G��G[K|饗�p��0���絈FR<>F��քt�z��ilnj�e9�YY����QLe~��X�38�d]�5
��X��j�r�P��;�^��%�+��_��k��/^�;ú.U>� 훤X����k�O{����T!�߶�}+���43�0 ��Tl�4�F���0�=�-�:�8pw�
�~���{N{Uv��$���x
& ����[۞B��g�����Cj�Ã�|I|�K,Dy
�qy�j�n��VAm��Bn���MIf�m:�K*N��x�	��$?�:����}įFFL(��I����iAK/٢Y�9s�ѣ������͑X�I�J.f��	GΫP���W��'KY�hrܲFG�՘�%����6��l��Da�X.b{���7@i�JL:�#�b�:���P �V���o�\���ioo�d�B�? nJq�;v	�Ǒ�1��"�i%�!����͕�{;I�oIZ��9�_��ڑ��o����0����+��ɾ��x�qu#�>��
��biO=M�D�ɕ�S��M����%ĕ���]_pGS�aX�/�$��~����G3n�����_����ַ�%9����:�S^��^z.�)������t���^7�t��8=�[?��a��1w��={8!b�ʡr3�x�1�:U�фK�L�:�#�][�/��/>���TH?-"J"Y/X�
'!k\ e�H���_����>��ө���h���?׺�S�����nݦ'���D�]:@+�u��o+վ߾^}5.�ZmKAF��۷�K9��#l��O:�O��>�T���nR��]v�T^���_ ��a�&!N�K_/9w������~����'?���zR�}]Z��"�����=㥸ے��a$Lf�7ig�@Խ�ϟ��z[�����!�5"h���-�IO}��4 �&��P�j&7mڴj�*M}}Ϟ�p��Ճ�ᡏ�_M�T���v!Q�,)aѭ�ܷ�r���c�?z`��v�n��vOS�=�x�)����8�~�Q=�[������4._n9d��y��׉V���|K�.S�KT���~�3]6����?��'~A��=�܃��K��2�P�(i'h	�c�y晍7j6тH��G��"P�B����o�i2��K�,�����M�V���CS�h<2^���ԛ(蜞��4]
."��4b4�"A��V�-��:Az������;w��9�7��y9�t�$`�%>0}kh+���s����1���-pѤ���$/�A��a�sk)g���>��Y�ΡU�W�A�����K7�f��X&I��3mZ�O�>6dQ�E�$t��JL��u|B�Ճ�(n'�������˿����������J溯]���y�zpV�����zW��ͱ5{�r%�.����>����M���8(�|~������=�1�|��L*�s���ӫw
q����@�`s"g,�j^����A�����/w���L�aR�£x.�S�	0�W�5�>� �?�#6��\u�&@!k�C�#�g� N�K{�GF���#��ΕW^�g�g���Y���{�կR����x�.ʮ��Ytˊ���8g�>�A]S)0.�]$h�R�jQ���\�6u���x��W�$K���c�4N�����V5���ٯAL���}�a��L뙾}�+�v�L�n��X��`��Φ���oGƁw�M��$��#\eRrΉo\8!i�P����ОC�Ԫ�I�Ʉ^Rt2�Z"��ի[�ڤ���� =��[ZZ_|q#��K��校r��o^��*K)�_�R=t��?)��rLgƒ�Y�~�~��~�=�&�u�F��=�.��`ܩ9:<�81�\�mT����� �*�w�w ��CW\qߥܕ��� �gR<��6�y�}� ���-ҿV���Bk���G��Ҡ�2�^x��GHW��FRH�F�t�pً�u��}�s��+��J|��'�(R��7]$p.Y���J�l�]��o]'�g�ncR����a�fM�D�.f����-E*�-a-�̴;�#��
26I��~��$��k��<��뮻v~s{^
�1ki��m�7m�dW�⻻�`Uhkkں��[o�����ք��t����믿^�����\ ����դQӚhk�k9��'D���,A+�IJ`�'!,��HTib�-��BG������ Z���&�����ص˗�ɳò+�j�ܓN9����g7���3Q���dKK��La}E��*�]N:i��e�c�����:ill"�X?��O�q([F��`��k����o{��U���66X�lהn���ζ��C���سo�O?%�;���w;M<u}z<#(&&��ڙ�������Y3�X�!Oj�����u���%ap��%=��Q��h�5���_���H���֖l:Ky���,�������ȑ����7]�w�`�I���i��)�]"��e.�K���d��!���Ս^}m7{��E��>i��-@��f-�,9e_5ze�˚��S�s���U�k�>�7�g���c���KN]B�q���4T�M��&��W���UW]%{[�cٲea��݂S:�����se	7j��� k֮�����,0�|@���y`��g��{���/�^x�e�_��m�o���1)�L����m���`q�)�Q�=G�m�htt2�?��?�����E�s�-�|�_��i�#S׀2^	ڋ�~�d& * ���[ś��X�.�F��"�FyBK+x��&�2��O����bTv�j%N�;{����@X��I�7�zL=Yw���E�����6���0r"�,wL!���:�H�o���ox��Z�_����5%�� &&j���{��W9�ĉ��<m7�c���i���?�I�>�Տ���/}I����k���G?��Ӯ.c�ӵ��7�������v������<�����ib��$�H��~��_'��\,�9{y{��E�Yx���g�%kI�PY}W/L�4f��L��f�,ٍ�1�mx,o�Xe�4�P�@n~PG[̦Ǔ���(�<�)�w4>��3�a2��Z�iX�4n�3��1Ia!t%}C#*"'�;a{{'�0�\�oB�i���B{�Yk�h&L�ԯ�����;==K��'��b�
�Ѡ�҇�LY�t)�2��>����ۗ6�5T]D_\�f�Ϳ������6��p�TJy4Jۢ�����p���L��{]sHƉ�e��{b-�A�3�-t�E�ؼ��7����5�3f�$�Tt��CB������q5i'��Q���_�@�z�L�ݶ��7��t���jtӯg�}v��t0$�5	-��#��-qӶ�z����X9�@�H��{����ǚ����N"����A@F�@�v�Tk�B�[,��i[��~;hI�|�g$�s������_��������ܜ������ޚ�����҃|�ӟ��.�!T�c��LZ(FY�`'�c�� �^�%���7����7}�!���h�'�b�M���7����lr&���h�.m�$t���\rI�!?�p�-A4M��F�T���p'����gj���gUV�ƭs��#$2�ٰU��4{�Y_��L�*6����FGF�X�����!�w��])6i�]+hh8p��	��8�]=����CgL�%���4�0�:��4?o�MlWWӐ���Z��\���=���������.�m��v�}��=�n��^^����P��)��y�J�h�Տ;y�Ԁ�(,�������3��|a��m�m�����YƧO�F�jժ�+W�����V	�Ԙ��(�Ƈy�����<{�݂!D��5����b�} ��Ձ˜��C�tz4J�u}�W�\����>�m�6���.�H�KӨQɺ��w������p$;Swסж�*h7��lh8|�)�D�����)��$�(�c� [��NU�Í�6���ɋ��R�.��x��][K�"O�w鮇 �8�c�α�G@��y�ڬ�����;�<���H;v����R���(�3UT��S=��ޯ���o�������F�K.ygO����5E��'M�gҴ���xS����E����R�*�$3_�N��ƿ�ۿ]{�˖����wz�da�R9f����L[�\��	�U�N��Zf�S�lr?7�e,����v"�ɑǂX�X	���5	i����x�CDE%�����*ƍ:�	�����mH�N��ʫT^�k_����UL�>��¦�r	=�qHy��$�D�R�+)pV�NM�S#�	��˒?gB���/܇�.Fo��#WKc����vx�����ւ�ǯi͛�$f��P�$���'�h,Ó��8 �r����������s{|B�)����Wɂ�w�D�Su���	�Ph���&��ב.{�@\�W��"Τ7����C>�m�|5譩I�~�e!x�!���t�_i#+�43thd8!D@�?�������m��Y��/*H�ݡ#*�v���!Q�t� ㌙G�cK1�i���y���=��駟�D�䕧Q����:�>����_��_Q���13}�~�3��w�+�uG1y`� ,�U�I*�Bi�F����t_�hSB!)7�t���4fo�3��b6�!=��ŋ5�����/Ξ=W�P�����嗷OL�54�0�C/����V{^ۭ�
�T��~���50�Vg�!Aŉ���5-�Yg�c0��5<)�3�8C�u�Y˥����3�$�(��;��H�kgΞ=CxEoj#��?��ƍ�e�̟?��^�a�2�a��V��?��?�J��^\R^(�%-]oR��ӛz ��;��y��'�؝;v��g��9~���BУ��,�&����� wma��R��g���Wr�Խ���8��l�Y�c�Ћl�n��G��΋��4���{t:��h�$?	絵v�ٴAW��������S{p����9x���)�� �ksk������hWw�ࠎ�ԩӄ���R	y�I]W1f�n}��ϻ�KwFǴ+z:3%Tz_W#�ѢEs��x����ۛJո!�K��hAK���⩧��5�D(��eO;m�6��ݾ�{;;:%�����.m'���ui��U�TQА
~#?t*�ԫ��kMֽu�V�}����{��mmn�C�$'����;Kv���=c=���V�L^��?�!~Ir|%��^�r',��g ^W8��5*����SB;T#��^9o�v�;��5F��������� �D$)��Ђh�m��]\��^�1�WBC����0c�wP=9{���9;I�g����L�l��Td�f�IS�UW]y�gj `w��{ߕw���_���Td�g���׃3�E�$�sI�3�;�PM�.���OKs�7h�_|�����TZ�ô� ��2<:a)?I,��'@�dT�|��l�9S���֭���V�	rIC\G�F+��,��N恤1��2uMB��pR�A��I��&t"Tގ)$��'q[������N��goi!��#���Q�����7��]V�MgdѢ���w�-["i��Ey�����L������Q��Mr��{�j�b���Z��|A����j�5ǣ�S���ᴩ���tH�ʦC��U,��Ӏ���2���Z{�L�m��6a5ÀJ��e�sZ��:����&!to�=�Z����8!y��p�"�2�2z�/8{�O#��[��>�%�9�#����F"CG�PR4fiߑ���Ik��/Z�7`�4���d�Y5��t)}�,l	5�I�K���VT�A�Z��������FG[�s�Z\@�$��)@_ݹ�W_�R}�C�P�N���J,�Z���Y�$%q�8gi�Kz��~��n߾��y}^P��g������<�M��k��{��v��#�ew�|;��o	�n^hHi�u�-�O&�i�|v�)��W��Y���/)�%3]H�;{��gM8U2�u�V�>�y𠑋���Ls��ч�%Rv��Yn��QrVš���n����J�������Mr$���2,��kO>a�O�O=z bXO�H&�$�:��5�{�z���7J�i�?���_x�;�V�cECZ,�y�ɋ�l��� i�1�z���(��u�.�q1J*i�iN4-�@�}������G>�-� ��;�t��^�	W�Ъ��l9��n�,p�-(6��ܢ1�id��l�5k��Fͬ��Q�6cKO;M�FNg��G���E�q^h]��
W]u��a`��o���ׯ_�)c�Z��>����NӉִ�]�Vs+�ь��T�j6����e�S�"ĩ��xe���,~ ��#Q����Z��xR˸�K|�ӟ֩�	�)	+�N*:�!Zh̓� �����/���������'���Jm{��o��C�C,D�e�lE!���8�瘷#r����98P#���H��Y�� �ѣ��2�<�*"��!C_�$c�ksb�Rf�0B��/}IӨ5ҌU��~֬�^z�O��������a�-~-�>iZ�*t��mH�j*��8�al�={hV�F@�Tq��zF1/\x2i@��ǽˬ���˗��mo.7�`����W���G�'� ]�0�DU��F���9�������٩���Z[�V�\��C�~�x%F~X��F4�W�A�,I�p��E*CGC���/�[���c	K�,� �d%�q���{���_+��A]�������g��0���	��T!֩d�;�(��# �@��|� 0�U�3�I*�.��Q�-�&�Tn��O�F�5S��nTp@w�Q�O�\�䐰"�j���O:i�ؘ���ѣ��ljζ����7�t�t�ҥK�'<[ȁ��	��ӛ֬�ּTI\��G�B��𬽣m��]��M
��=���V'h!�\3>儔����S��Pu��XG:Tk}U3I�$�)LQ�\3#���m`{y΍$`���dA%�`2����,xs'�L&a�f͋�����x��Z�m����|�P�O8�c9U9 	�?	<5;�b�d�����ب��."�':�W$�3d>�y�Y6�(F��-���Q�U�"c7�xG��\�������̚=��e�#!s�M�r�=y�����KH��]t�5��ҏ<��o�y?K�/��RW��
Q�ᡡV���EB���ѹ�����[6o�x0ڈ��N56/b�L�~��!}M�,�J6��r=��-[��G�R6+Q�5,���fɒ%���諭w�=�SZ�JK��K/��7����>[��_��ub:��	����o\<�ɦ���l<c�
W��I�������ǟܴiS�@w?z�H��w��]�w�����/�߷/׬�h��q�$���n]Y3����?����}��Ad'�i��p�W4�4
^�{�UK.���[�6�tuu��K�O�@�X(���}��g��F�qbU?Gi�
��%Db1͌V\�.64�RǪ��ӗd�ɺu���)30���7a����,4��󓧞*Y�T+葈���:��%�,f������w�H"�,&O?}���7_�JP����-E�� ��}{�
i~�x�md������M��|��;������,Є?���_��W�7�[[�T�u�����}:�{�������ro�
�&J��l����iE����R�ݳ������;v���F�	v=�A���$ �����U��� b��_����� �%�r�˿����A�iwv�: �! ӑ���>_+[��E����N��ڍ��D!���}���1ϒ$:�pJ�[~��ih�����[͉�g��S���d>ii~���4��+�7��Ʋ�wn��{���z�Sʙ�*A������vvf���FôS~1�o���Ã2zǧ����3�0:V���d%Z.8EsL
V�9Ҭv�$W%$��x�TC�h�+�ܜ�R@	��y���bA2L�9ς�W�zxvL�}�oŇ�J�y޳^<��Ks��3�'HV59�E]��§������Af���/����n�������)N��F�c��vƔ~�6�,K����c�����i�ޚ��_�~��Z�5�gLTk�i�x��I�+�4�LR���&��`	=ŷ���:�ӦI�g;;[��r6�#o�>Cو2%��{�5a��3����SB���*�#��l�64�k��,E!��/����#־��m�+/K�LƵw��a�9����/Y��xUj}-��5ɸ̸_�ZG~�ߞg��!#��H�r2�-�I�0&7�c���߀��u�����b�>�#uD<)��g$y�TP"e�����^#�r��N�("�L������G]N;Ul��.���	ie�Rb6����2�x?��O����|^�_���,�T��$�tS��yn�V&�s}R�VƫƠ�������{@�U_g����}F�
� �!�)�F��!`��l�Il���a9q�Vb�4/�8q	�qp�`lLM��*���)��o�~{?������Fs�=��e�g�gq�������d*���p�Al��U�`P^c�wۼyJ�U�1C}�W�z뭈�z{zf͞}�Uڢŋ�=�<�5�j�!(3:����	�|2N�QB�Z�� �]�a���� �6?)&^(�`q�ړO>�Dō>c�Ў <���*�a%+��T8[�~݃>��o~��ե��!�}�+_a�9rT1 dz}�
 Sq8k�; ���ꫮ�����k��������2�oOYe�_�Ĺz��/��=���WZx�O��O��w�ᬳ����¸g׹�_T�0r�[n����jiiCK��T�b27�A��r9笉�Ȯ�S�(&\q�m۶�w�}���i�'ϥ�`RKl��**�GU��h_iaժU�f�p��9ݽ�U�>,1�����tt6���m�]w����>t�(p���|����'�h��`%�q,2�P���!�}�}g�y��?~k��^��5�\�r�ַ����w��� 2'���O?-CEmÚ��M�e8�����x~����e���X;����0�j��t�R,�<z��͹k�.&*��Y�/|�Gagz�(�D�eS��T��y�-�y��s8"�+GF���Q�*U݀VՔ���(F#rV�S�(����	�I��/�����|�}��9Y��Ww��"�+d�
�1U>ǡV�������)p�J%Ie�X+'kG^T��4������n(Q�:�a��20�u�e~��eQ�;&<���ݝ�@�p�-X��<��,é�ӭ�4m![�����i￩��hLђP�J	F��mY:D�
�$5���	����kr�p2���'�LJ�W�_ֹ�w����e쟴��a��Ύ����5���>&D,UˆŤA��e�_�rA��E�?Qoۅ`D�|�� [lwd�2���Me��ʪh]5yl����а��M��AZ�X&qy�OĔt^�b�� ���R�~f8UTȿ��n�3I����	��Er�|��1�1�l��n���g477Ej����]����*�F~b;�Y��/@,��Y64�:��8��56f�B~w;�q���-��4�?P,��ƒ� �R7�l�h�I�ܯ� �'�X�&_n�!������$R�|����^� ���(�m��C���k(��I�jI%�#t�[�\Z4��m����_(3��a�Ks�sHμ��B	V���p�c(��f����т�[2Y�>���3�;���{6LB\M��{��A�rum��˫��
�Iz�Ϫ��) 泟���Sa������S�cC ��_ ��y�+6S�D���"����f����T%��G�[�#�Uf���f�J*�elH��y��ן�hB\�ȯn�d���%�hԉ�@d�3��	Sف�tX��۷+�x������B�EY<�� �:Fa0 ,h&o�"=��1�ˬ�3�ic"��c�RIS-Z�����G�OxH��I��; ��SM��0C>_[[��|ࢋֿ�������6l��w+�ܾI��.k�Q7��+����2�<Ň?�a�?�@��^z)3������}}�.;�U)�'RWl9*�0c�\�eE܀��G�v/w��L=�+���E��!yF���I���~V���Uٱ�93�[�F�'(��H3yr^���ۿ��#���QSS�\1:�����'�'�����ڵk%�<,^!"��:>��?��#�����R�b@�������[s���瞓+�ugV��o͓_�0>w�r"���g�P��+[6#����^k�.n
��H�{Z����
\(ѩ�+u��R1��������޻�mn�˺�}0�w�b�Ν��\A�dJ4a����UT��-җJ�b�2{�]��L��Ɋ���d��A�K4�"L8[Qi�|W)Y}��&&��H<Q��R�h7*YB)a;�{D@��O=��H�z�_=��/�����RJ�����Dżr���N����P˖ѱI��'�W̹����suffT#��`�U;u�B���j#��ܤ�b��7\�u
$�{ZO� j�r&�t�v�y��U�ԕ+��?�2����J��I��P��Ug�ő��ӳL������+R��f���x�&�Y���Q��X-{�[���ϭY�-�Yl��X����D���E�iLa X
E�&Yg̚�n�z\�r��H�v@�lS;X#�K�O�>@*bK{k2U"�߳7��ǐ��X��J%�a:�L2���cb^䫀�z������*A�ψP���w�����9��}�_���s��\wuu�י����?/�x�9�kF�1�Z��+�&��
=�*�INDs6��r6 �D�*&6�^�b^�hU��z{�Ms��x�`�����d["(WM�7���2����Z㼇�X_eʼa���X�)�BM���uL����0�7
����	w�f��(����3r!:��%������\�v1��2�z'�F��JͳmL���5z?/����O��2��诼��V�jU**�8���[ot��]y%֕X��{78$�z���?n�p�`<�����}򓟼��oa[�*�����o�Ɣs#}�dv!+�z�3�/B���.g<<�꧔���򗿔�V2M��PT<�i�B�XS#�%�/��i��O��O�eǮ]jY�V��p�ET=R\p��[>���m�֭�`��6�9}�kt���^���}�������)e\���]s����x��o˕o��m��cI5LrC���o۾��+�'%%5D��JI�6�ѯ��6�1H�Sɟ~�錖Y�pb���ޞ�)S���9p�ef����+���q2]?���e� S��j�������:a��׿�u����a 8m��s_���T�U����?8/���� <8�d�`DQèZ�k��'�N6?����:O�\�b�)�ͨCS��bX<��ш��d"�6,V�:gN����l۶��fe�!�p�fK��N���d�"\hc>re� İ�r���:%E|��B"���<���m��0{�	^#|D	V�CB=3�]=�JddۜӎGFuvv�\��I��^d��[v�����,�h`���C���>�'U)��$��͜5��º����Li�����Wn~p,+ư쌥bg��l�_���B$�(?>1����{���M�2�'��bjDs}A7K�rv)B��7�v�,���]:tL��t���{C�X5��gׅ~���A�u��-��cǎE�:���7X}C>�n2ϟ>��o ��;}�eb0�\���bB�.\�/���EKJӲ����uل܉;���Ξ%1b�%�}��M��G?��*������&�JjlR��X$��H}��"�I:��2��)��$ml<8�}��=�Ia�3��
��Qn�\:놥9w��3���fi�ʊ��E"<R��P���w5�7�^��A9X�ᣬ҄�ް�3�
����$fE[�K,s����I��?%u�
Z~���+l�,WX@?��e�Y��l>'��x�tW�B�rU��ТV�f�Wd�#����(�㻊`b�0c�|���ZA����^z�;�}�!�������i``xl,#�
����k�3���ԓa��`n�+�*pg,ɨJ5y^6�����
_���;�ٚ�%UU���x�Hj߁���B�"�R�Ӱ��RN�j�?��(�L�\,��nnmnkjh�þ���>mxT�fE�
[�T#F���
��㼩B����f��ږ���c�]�h��hD.�����r#>��N��ݘ��3��$�2����#�M�C�h����۷�9�ˀ����žJY�zwG���#��U�Ɍ�ꗿ�D�|$�Ѫ��?c�r>	8۲y+�@Mu��"���\{���xd˫�2�Y3fX��ҥ˗/�7,�Ƣ�%Fx��Б�ʊ���l߈�^��*��9��:����V61�R4n���a~����ҽ��^�;�3�n+�����>�nYv�\�ԅs��+B�
����v�
~G�)��ޤ�3���܈)���̘[n�E��4�C�M�$"qV�X�5Է
�q�����	����1��3��3<cf�N��U���k/o�2>�N&���l��N;Ȉ���mX�Ȳ�8�HU�z9���U�V�S����q�������ƑJ,���X���R}K�,�Ű:�H�����n�\.㟴Pr�LS�[��͛��s���������>��w�VP��7��q�	o�}�)����@�wn�Y���$̪�=e�#
��_��KҌ<1L��3�\�vm�{x=uR1/�ƴ�{�۷wo���h<q�9�b�d�`�4/��n���ڵk�j�GG�2���zc�Ovui�:ex�ro�����U���ʋ�HĢA4�Ύ����\�9-��b�XWG��]��P���H�q�l��E��;��X�3n���=w����Vkij����6e�)�k�jg͘����րΈ���:ڧ��f�',�9��:�b|���ꚮ��x,124�\�V5>:�J�S�����8�w�k;�ۻ;{<��j֌9g._���B�q����a</�
Օ�c�c�Hlxpx���m~$g��{sey67���Hzz{�8c����������ٴ�7d��]"_N%�y��|�
�6��hv�\�l* v�y�6��^&��>��o������萕J�T��J��8B@fh:��w�,tuwUUV!F$ߕͨ��\,:42��?�_20�c�8�v8{��d*>2j"�56>"w��~�N���T$*��Ne�⑸SR%���Q��N��L�V�x�������)SE�8�ū��i30���9��70<42g�ܮc]ȞH!(�-���S�F^�μ�!��'���ȻbPLy���U��*������1�s^ �����S�S��F�]w�q�h��HaN�Ԗ���i�5�ag����,�S�D<��:��!Ǔ���\]C��DV
>R��Nd#qˬ����x1��JŃ|���flx�7�����D_EY- ��B���
�]\���|4W�`X.`:�~a<� ��G�p����vM1���d<Ŷ	
l!�N�����j��1�yT.��gsپ��b,�)�Rɾ!�b�<�f?�01*�<�OD++�,R���8̞$��فHu��Tʘ�T�\]����}���˗=��3|E�k
�)�B�+\��nMـ�y5r��16'���c�ʡ�B[[�,^��r�h,�H������������E��X�h2:61j�����:�s�,�!�dy~c�ìco��d,��SI�?��N�r��!��h���?�{`���g�G�aD�(q��%CG{N]�&2Ea�
W�70Y�^��bq����5E-��e�������uu�?������]�v��a�f�/�����^�����TN�W3dE�l�%�'S���O�c,2,�qϵ����!�KJ�8Q�����W �m߾���[������q��-^j�4^]]û��`����=�\S���_B����یq�8�w�޳�:K�(���c~T�%�)��3l���7n���@,�1�VA���﹚(�3��]/��k��Fi�2ݘU�)���+
�W����>��<Ё���M�ȇ�:�t��z���<�裪�MO�.g:���I��P�!,fv��kP��o�[�:ի��n�EOO����Eu��ei��y��iӦW^y�x�v�әX���q�o�
q�y�U�-*�;�����b�Ͽ�Q�
�̤Ӫ�P~���^����-�)z����^��`7e!�������5bn�M�e�bT�/�nݪ�HLT;O�x@r�����'ꀕ��5�X(�&MSUQ�TѦ�V��Ɩ�6_���Vbbu�\�9�XU��d`�r9�'QU5b��^��l��Pq���k��_0��2Z~M��UW[�9�+-#
��Vd-�1,���b�+�1��2ٌJ���jD0Q^`.�klhT�2_iR*��~�����ŝm<"T���z��ҙ��y�ÜqP3rdEX�+Um\����-�j�-Z��Ъ����ƌJ�شr���Cb~��	g��B�	7�N.
U�+�ͫ"˝�	1��(}�����D���]���"r�U{��k�������S�z�.�..(�D>������dh81��|Q�#��򫔻̀�W��{j	��j��O����ZIlo����j�vT;˚�N���Y�T���H���=��b��C�F������&������oE�QdT���")�,(����ѓ��4$�g���	��0,��D:��22���$N��������"'���wrA�\ا�Zd��={�C��>SB��l���8��Ȗ�����Đ�����
�o��O�Cy��S�˃.��x��2������G�2[n �u~���/Y��o�@ge�ϟ?����﮺�*������v#ל9s&b����� �_~9�3�l*x@li�T��!��rab����
yȊ�n�Z2�ʮ���[`��*cg�Y���hTRAC���򪍌w\��bٝY�T��?@�����r��+�L�*;�-�D�{��&r`�3ZlQ��ciI.a���v�
E���b��cRY��`BḌ~���s�)h�@�d�EЛ��ʞI=�@%b��W	�t�Mmm�H���uy��u1gA�����p����G�玬9pp��e�30eR;��ʖ��i3@[uM%�� ��������V��9���?��Y�$���Ct,�Bv�����F�V��U;Q�esi��X��xu��V(%l+�����K/+�=B!�\�B�I���[�Ң���G�;5t��֓ʀy���k$�i�ߵ�^+b�ŋ#�^۲����{^&cL�qlB?��x��7Q��WUD�^a�5��G`[�K�T��u��ݠ�s��Ή@GNCjs�6b�@�"����Ԩ�ҡy��ZY�^��_�g��r/��]V�h[����2��^5���"������ã�!.�g��DHs(7�EĆQ-[��� �0N�}.[���k��O�� e�B}}\��v�L�6���2�ȩ���ɲc�.f��{bl��rr&��n&6��t�]���8���Wyv�Z��������С��|�;�.վ��8�_a����3Nl�ٮ�$�%C���_�����R�m��ڧ�306�5��S�N���~?O���K���N�r!��y�Z����̕���m޼��4�7�ݷ���UIa\|l|�k�:��IO��L9�(�,��U��p�I5�h��9B�D��Qoh�%g[��h�evj�Ţ��n��r
��/9�Npt�8|���Uµ�9�ɛ ��L�;�cN�:�
 �(H�=|��Ւ����sg��� y2�Cء$�{n]WW�{��M"3@��՛8��B�!-u"TVo!��1Y�P�cS��=08���)�U�u�#R��A5��"Z�0��MXJ�u�'&1_Oܕp.�P��S��b)g.��$'|��!�d�>���O�.���VpF!6m3ý��C=�z�j֗Q0�ʑr�Z��r)Ⱦ��5�o4.�,�XU!&�b�䨩	ԒS�Fo�����TQ�%�4�^�.�A��76��/]��o��o@`Hf��p�tS���P����_a�"Xn�������,*�>_Yy�GWO���[1�� |�H�(XՐ��
H�]6���T�H
K����j������8[(�2�6澠����dF�R*.����^��c�M�2R.���M�����O��
;"�i��[�2#��-�Ui[HX:44�3�	�Rb|�xU{5$�j��-�!�Z9N���s�Q��� .q�Zg�MbZw�~=�Ԣ���n߾}���C� ���S�cʮ��'�*?L���uL���9���^(��K����[EĪ�8c�F�ވW��\�Q�\( T�j�e%[�+����g�� �q�=c��V���y�V�\�#�Y��h����)�MM����@��%����hɀ`J�:r��Gn
��P�K���K�V�`��߿���r6��w��G����/�ؘ(��_��,�y��@L5�^v�e<;ۆ�iǁ�3�5�<����O3@ϩ��?p�r���$H�9���u�:;#�v����:�W�ٙ��3g͞=�'����J���� ��l0<�(���Yq[v-�"�������d=c���X#N����==L��eL��[<�r�O���y�Rէ[o:�~�:;�oc�ң�>jI��=���䭍7>��#*�0iu���D��<`�P,8'gR� *�H�f@KrL�%��?���d��W���G f�ٰZ�9x�$_��"ݭ��3�����_��A
%ӳ9k���Q��v�h{F�LM�::;�㎵k�r�8/�6��}E2����@�y�Ƿx@��+���%C�<"�Y�h!��/Z{b��+�,�#X�/^q1S�-	q�f$@Iv>0��*T��ΦUy 4�~'���I��(TD�v}���9O1Ε�;�FOSJ e�u{FU�b[U�R��rGN����*��tBl��68pD�YL�@sT��KC�6ށ�{E�!R���s��W��F���ȟ�JX,�`���I�y�t���[#*eA�3����ʑW��|o��X���P��x���m���&�tK���sapb�u;˺p�\.��֛�$�U����K.��{tt��|�k��?�*��r�%��H������[��n6�M�q�nT�|	�Lr�(�9؝�?3Y�!P��^U��#��<�r��+eu(ׂrY����7%�WW�6�ԱR`���k�(aW�ڡ�*-�R6+��1�%����	>�ћ���8Rj�b�K�8�	҉�:�뮻<�1P��<�ߒ3LO��"��X_�K`�Y���d��<11���(J�?�I�k���ٿ�m)|��8����-�����x��Q5GKf��U��'���e'R���	@	���~����櫲�:�9	و�d)U�A���jE91Q�ʣ��"QB�l�`�q�ZZ�=Nj1��wm��5��`h`����� k������СCL���֭[�10 ���v��Ȩ �P`��P �\�r�����UbVX,s�wʩ.��}g�\a�4��eۜ���ẽ(o,�O�"�d-��H(�h5z'x�5�E� ��L���%����.`��[��].ũk��&�Ȏ���*���A�
�@�|�ͫV�bJ��|�r��X8g����b�+�ظ���:W�YA��{lJ[;d�yJ�y�YR��Ч(�[��ڹs�<�|�1�L#O��@Ǻ����|ȸ�$�K|���U���-^�,n;UgK��%�IfLt*<]:�y���~�a���V22:b�g�y�駟>>1��>����Looo�ԑ��5�>c��g��e�F"��,��~c�7z<u���")�B��%O�y&�M$sEd�[�M	�RL��6�Wl㒘L\z�瞋Tڴi��Yw��G�
X�øG�o�αja���~ )[�����ũ^G�']Tqwl`FgP��_�Jr�j8H��DFĄȊ�ڙ��֭[���ӟ�Y[Ui�����/��qZ�/�((<x`ǎ�&~�	O��:��	��B�W�M�����y�Q�����&��f`]O�����9/�n9i�S�O�	0q���b~�L�+�ȮY��_�*5��g�s5*�q�׶����w�|�T�t��@��͛`�Bܐ�#����HqBU�'L�Ne�r�q5��"L���Ro9#/��>C����i���,,�C�zn�X����hd�Ϡ����}}C[���D�6\�r3�63$g�<�Ґ�t�z�3��R�E�\�_̡�+Io���L|Le���y�X�sv$���h���h`L�	���c��$�8�է�f�����^9{��9{���09l~6�����P�p�]��h����1ǒ��<��.���W�H���:'�Q��=��%����'�!>�<��Pi�3��@8 �"���Ғŋ��r9��a\VnN�����c��N����L�%��#x��w�ofL4P�FXL�
�>�\�����
��c�?�S��+�D�<��Yn�觎��NTK��K���F�Ϛ5��w�MǴ<M�`HҼx.���J����K�e6��
�sƍ��`����>�۔v�&��8'���9q&#�H1p�ʘ���]Ė+LZ����,2�.����X�%#'��5��aCZ���� [W��&�C"9.R11�+n�A�Z$���b�\�M�P�p�Z�8NFƴ����g[�Lj����Ȗ���B��l$�gN�����E�=�裿a����+J��zsS�p�������	o����K1�x�@=ϫ`"�HfD���'�SN9EM��]�y�%i����sι��eR����駟6rO���@=���i��dԂ����	䡺�hM�C�&S{1��������ꂊF��rȉ�c�_^]5��v�w�}7�����+�tø7T�~�J	�������0��b@�Tx�_<#�W��A��S T�Q���򗿼���V-1���<8;h�a1���?�m�k
��X��<�s����}��3r����8��͊]O	X��9�F�v��g�}�M7]u�U�c���u�9�Vy��g�ڵk3v�m����W��0-�e��O�(=��Q7�x���b@�� ��=`����h֟��Sd�*�3��b�C��8	S1F�I�x49_��3}$,.�aW�E�M��Xm��/������r-!��wqGV����%%m��nhl�gs�2�ġcW�-%��{&��ի�C������&hR�g�S6j�LZRY�L*���Cl~��S�w�)���
7e�8�\�i� �E����lH��d2�u�.Ϭ�F������"�=s�����B�+(��x����x^�
�9d���A!99�F�LV֦"PL�l6�B�]<�h��t}�ߋN�(,���%��`4O��3gLcx��j)�(PȞ��?@�4
}N�:E�5�Qu�:��S�*6y/��M��bI�B�!	p��r)9��Y����{���#��OB!���A����s�Swu�$J����Qu$cc�#�v��:K׽��!�����{�H��b������!8N��'P]x��~�o��1��Y
'�94�KQ��C]s�����=r�+:{�m�-'�j	��j!E�,�|��˜�,K)�Y��%���'�^,w�W�O���l��LS����N,���} Q������կ���b0�g&5T��x��>�0������c�CCi�L]Y�G6ee"�(5���	�|'��Jt�/��A����dLI��T�8r-���4���If"��3y��+x�L��v;���e� +�Ɍ�c�i7Hd�X��b}]c���^�ٔ�� �PP���)�\����e��O�*x�"�3fX3�SNY o����(��j�k�z��74<�tF�9�F�Z���#��f0(���c�o>��q)ĩ�I��Z�����$IA=���BU<����.eɘ��]��}m�0=��s[�l1R�tZ�3-��%KV�\)�_�Ss��11������I]6�j÷m�6�0*�����R�7oF��t���9��U++٦�6�)�/<-r�1�(-����ۿ�[�[���Η/_������	��3�g�;c{r�i���AH�>�ĉ']�b���rq�%���]��U%"�`��:묝;���1�3���Z�k����[o�� ����s�1K���{���g����[���G�*��&��hni<|��;v0 v�w)����1r&��9��P���޽��i����S���o���-Z�XyH`��zK>��������d�܅a?��C��	π�zꌜ.,�]�a�������d@H��`�F$��k&p��` 6{��揿�����)S�N&�`6zzѢ�[��E��ڸq���k��\sK=�����	'�`��ݿϸ ܷϰ��gϙ���������M]}]�lI����y
qG� ���[C�SO=u��cX��/<]��SOY��8 !�����JDJ*@v[%k�U4�9�ӭiUbǎ�\1≐T���v5�r�ٲe�/~��j�?c�0N���_��޵ܣT�B����O��LΙ�@F��T��,.{LB�0-Igv��D8�ґL��,g"=Q���������Z9�x��J�2�,�Pl�W��y2�
��;����W�>���X>��	�u�wȓ')�M�DEx�}c�nooWB�s�4���E�˥Ļ\.-䐢
�Y9'�B�Ə��*d�:*:����g��C���זmɵ�͛s�m���/"[�Ҋk7
���nV+N�!�P�Vm�P�bQi��3��S-������俄��\/�R�B~R�+ۤoM�w�R���k���?�� ��ܱ����W R�jEER,�*��wF9*��C@_GK��'e��s� ) �����d�؆�Fg1�u�`�Q�	��|�%�?zA�E6���.R����G�%Q�.YH0�6����߮Xq�{ڊ�z�H.Q��dLM)�S�� ��x�Ÿ��Y#�H�*FG���̡��(ƃ�D�<m��y�j.�N�m�F*Uq���&u��:Z�f��Щ�8�x��*�rN�@i�����Ņ��\���r��6s���x����l��A�#G�+X6*�T�B��rMѽ��U���
A�f��Ҧ~��lڴɅx�%�����z��KpGt	'�_@	�V�1d
���ۃ�B��u��R�Y���(���1qYt���_E��4��R޳E0���/��r.kf�$��k�tb�l��Np���-=�E��>��s�9�ଭ��p�d)k0^��gx@0��!���vv�kdx��YX�y�g�;O�!����ېi�20�,r?�����Y\�5���P��T[�a/��/��� A�nnh�9�J=�SD��g��VanjK̘9�k�jo��&bB�>h@9s��>cgD˕�o����P�A9e*�ӯ��*_��-[Ƃr�2kɘ��x���>����^ۘM��}���v���ҋ�� $9�w)K�+犼�--���WŌ�Բ�IVN8����U�u�3�|d�7l؀ b����e���Vd�n�!=a�n]9���
'e�sH��l���A�E+�@g3̘�-��%{J��������# ���}�~���>�1�?��O����*����+NG�𙶶��;_������Qg��as�&�{�;*{I�nSшi u��A*+����|���'7�H��4g_��}:bl�kS E�[����W�n�)�Kk>`mˏ�+����m6�2��=�����e�����/��/o��Ƣe+A�za57q#m��|�CV��[�5w������T|���V����"Oq�dN}� 7z��	}]ǜ�}�����r���������Y�:$C��إ�L�g͚��8v��#�p��xL�/O�HnyX��s�1� �Fg��>�� ���(�^��Aa�a*�]�n�D]���J9zU	����)��Tr�D]���e����������R�@']GL�k }~�m��͗]v�x�j�� ,����]�齼�to�
�j3C���&����]N�IΘ`���7�;�j2�u�ҙ���F��y/o��l��w�x+,���p�BQʅ~bi:vN�d�����7�FR,�O��#n��8��L��P��ҝ'�3g��<�;w����}��_��_s6�8� A�|[<|�x���O}�S�����/?}t4-�+��Tbl���B��Hĉ),�֒�*����X)����t�;Sb@d�sgZF��Ö\j�R*8(�������<���J��~�H���ќ[�}e�!�fӽ�^�Sojj�?�,�E��4
������A���w|����?opUm5�~�U��|U!_lx�L����>������Fn��mM�ZZ-�A_�\��,��#j_|ᅸW�O�����۷����mSzF�5�`8�
"D<�<i��@]�q�vo���Q��넎�6Ɏ4��n����m[~����+�T��fRR?;�2��5�
/�dHjL�5��B~�.+�lhl�@0@Ge�b�b�]!�����䨑�D� ��2ȋ�0���)�H܀"~����PYH��
��+��+��$���`�ƍ �㧷�+ �x�ȁ+���h��`�Y�wW�J>J�Ȳ3�+���+�R��ǁ,zn�v?׭[��Q�jɒż��5�V�K��I��������o����A�������P<����5Z�"�"�Y���Q�]��eb�%A����qY��u�]�*7�N�T��o�`�)��%_c��X�7W��������+YDT��O g��l��0�o���]t�y��u1�W]����ب8�Al����cfc(C����SO��}�#�����K/�Ē���J[p�C�UVTbN�z�\S�o����}2��r�.���z���G�/�W��K��L�x�R��kׂ�Yb���}{���0�����&9�3d�D���/�!n��n�����4��y��g���ouuu�LL*���Ш�,]v�%L��O>�zi���տ����v�V�b_�8?�я����I�K뫏�@ 2�x��1���Xp$���U��M�T��R(Oy�	u9�\�a�0��;Ԩ�?����Ո;fU�&�UM�* %��a�we��֒���20`e�|K�Hv���w�h����|�����e��t#��t�
k(����������lc�h��G���̬�T�)��+��sE������QԛYRH��c�(T�;�G�A��2���6(�2���!��F����mA��6kd%���̹qg'
E�c�(�'�3g֖-��r�!��JR�>8��*c��+2).�G�d�+vLO�n����I��_<�e�ٵ�y�����|.&N�c�c�m��cN{�rT�pf��/���dL�D>�
o'-�dr��dԽe6���$�b��X�C�MM 2�]��Q�^�,�^�H_�wv0f$�)�_�F�k%7r�AD844V[[�d�\�y�~����!NC� ѭ�Hᢹ>������^��}�~�U��r#��=!�[ݑL)a �߁�����U<4 jY&"�2o� fO$O��,i��T<1>2Z�l���s�UJ��|!�M��R>�ڏx��z)�8XX}�X��0����!��*��=M��,%��.����U�����c�P�Io;��J~��=�s�o�;�=�t$NuRx��T&���);��Uy�ou��pN��{G�Vo���5�\��sWP��)P~\�]����o��oų��̚5k��$8	�z�i=�>�,���O5�CE��:��� �$���(f��x������Z��^���aɡ�[���/���-��ݶG�ne��M�R�D6��pܲe[�z���Ʈޯ�hW�X�"ʚA9!j�FL5�l�����^L)��[�R2�cT����e�EP�M�~�	ܳ�mF����w����;Z쵢�y`H�>�([%�b��c
�#�:d(__�䔗_��V�h3�a��dL�^("�����{LN�0SX`���/Ph[^OK�vwzHm/��@�������ך�77s)n�_��C���#��~���޴iS�j J|1@��U��#���<��¢r<�2���֭[U�)�"?��/z���w�����������˗/7�d�Cg9�o����Po�frZ����DH���ﾰ�{���K��bC��TԲm�V�L�0���qV���G�R*w^�+��r����~��L�U�p��']��\-�D�r2�껢�~���lp��ח�K�p��Li�Af6dm�o��F^���˜b1��8K�9t*��/��&PΐxX�9��̳�
;�D�ʘ�N��e��A1Y�|�7��e���բd�x��eU'�z�K#H���-�r-Q�)�iկ��d?8��.v�#�/�G�;��������Z�
�D�L/�e�A����p09��f��f�e�I`~��*L2PA	u�R�(�x�al�$ʻ��������)�쾃qM����K&7��r[z\ep���\�(SJf	�ބ@��3����1S�S�@���)���S� ��yV���j��ޯݨ7-��)���C��
�y���^	�'�L�aAI,��|!������w)�[��)~�X��_+���\8A1/o�t���S�[|{A��;'�XWJmb���.�Ȃ��d�	VHT�S�ch�:�fF_��2l="�&���Wup[[K��5����@�Ϯ��|������?�y���hy�,����E8gA��U3B@>��o%��x,5�&,�ז�Lh*ԭ�iG6r#����Zi'�U&�{͔�W꼧�����'-�f�$��;�YtG�%���B`�-`�r�+�����e��I`,���R{r�[���,^Oo7���5+GA�ӧ�K(#(E�;s�t���e�򗶶ֺ�ڃTT�������Pq������0���,��>��/U�R��	��O�zΙ�@E����HAQ7
�bٟq��ii��c�X������c	��y��u��n����XǑ*�Ө����z�EqS��^��Ꭵu+;�U: Vؙ3gL�Ҧ�|[�s��bU.��������m({��O�~����^��˓O>������}w�駟��a�x�LOO	���5���F���B��;_WgG��?��s/�\x�ߵ�@���;vĽ_��[�D�W)^z饖�<s&�1���Ȁc���W\q��
ڋgd��q��"-�A6��ꪫ��JS_x��zc��Q�	۹�}ц����˥d�Wx�^��9q�-@�<#�m��5�w˖͠��ŉ!���ny��P�<�������x|܈6�]���HOd1W�F'B6>6*c`E� 
�p��-[&Ǹ�����d@������n�\�f��R0$.��2U���J9(jɔ���*��`U(�1����^�=��3J��>��>����v?��Ģ1�7c���,���Գ�Q���YP6�3�<�����R�I9'��'k����p��A��<C4)8������r2�K���)��-�vd�=̒�R	F�Pf>����/^Ƅ[#��6�o�1ϻk�.�}�{����٥l�k�h��Qe,1�w�y'�hﾷ���х���ij��S�W�����e�P/���.r~�F<~q�g-�/���j`><���v/�&�u�J8-I|ԺȀQ%�2[�XP�*R.@�:ƽ��R�&���q�o�`��<x4Y�R�D�@g��u��eq`���<��TJ_p/>�.CE�D�p)��~���3� ʱ|gtWhؕ��R��%b��D$��\�iٴ��QO!v�_|�?����}m*T��.3TMU�<����Kc��G��W(���*]���´���{�nL��b!�<=E4f�Gc�6�|�L]q?;A�ؑ@L���2�U�'��S�� ��'�@,���J�A���,��f�tTQa�r��,�a�\�����x"i�2f��C�S�"ܱ�w@&������(�x���|G}i噓�$?(�G�7�|���R�@J�2�k.W��7T�vr�Y�&���?E�VH��Qq&b6i�JO�m-V���V���"'p�;�pb�E
���^X+�*�D�2ȚW��[�ͻSф��ސ��C�2�*�vG9���[H\)�]����Ʌ|F\��Qe��d!��X�b��
N�2��y��:��rwW׏��-[����V���ޛ6mR�i�|�.�|]����t�e�7ʀ����F<8��K/�W������O�c�A���7l�����_qq�B�gI7�����p�`K�Py%;�[��l�eT)M�f�A���|�f��|�M�'26�0W�\�J�<�Rh�S����j�r1R��ypA��ї�,�&�Z�q���;w��ꦞ���y|N6�,�446"͙.η֯?w׮�A{<�z�kne�r����� -]y�̃��n�p�[��]�@����Ŭ�2!���ɑ�a4�5�\cAp�A�#A�0}}p��|�k�t�M�>��<��mlj��7���8+^]]�@۔):X�SͲ�'*,����͝7��{��%�VCd�v���+��Tr9��U��Rr$�ޚV/�Έ�D���[+W�d�S�Y0��G>��}�{��D�!~����/��d��ں���<Q�� ��h�������W�
J��?1a1#�Λ(��3r�L�}S=�i��:�
F{��ش���D�gKK��ݘ�~���V]���Bk��@�<�8�ޭ�����z�,]�t��u�l[�b�9��i� �|��Yw�O����:�I .���S��B�jj���m���)5 ��JF$�5�\������'_�^����o��1#�ho�ªmݺ�)3��d~��,�$���%����{�4v��*�r��$�M�b�ĉ%S��p��S������-�K��S��z�rX����;�RBŪfe��c�� �T�'�a9���z�W�W3x���@�������W'8TQ�������j6�#�Sӹ��*E���
�Ȩ�#{�����N�_|��O�cdR5�䙙�O���[��Z��Z�:��Ƶ���e|�$\�3pB:4~�,)R�r$��SuZ��T��ԫ�a��&�W*< ;!('�`Y]rɅ�O�|��VL��m�u*�a�S�)̊�2ެ��[\p����u�������Z�(e�a>20�Z�k_���y����ဪ������V�)��و�7n<��GP�r��X�r�syI?89�����S@�DyGi����i�+�D���Z  ��IDAT�b��aشz{�\���:�d�����Վ�,%�I5̂\Άj��l�ޕ�xhY�Z#�C5�u*��!���)O���L�d�:��l��F�V�={._?q��L1FuLq�P�FȞ����2e�Ux��Hg;��I�����ԃ�c(���le%��>�l�In*ysY�y��������\C�����;p�|��[o��Fv�ұU�U�xh�4k�v�ЌG�Ljsk� �a�FX�~=JB�f�O�W1��)������
�����5/FiԊŨPC��2m=A��������9B�����=oOoO̪��Ƣ���R��b&��W�������=\p�	o�e������K)/ �	�"_�̙�>�j J-G�+�c ��
yuv��yt�ĝ��	�M�^�<�-f͞m��UӰ���͘1I��}�ٷ�z�]w�6J�,ϸ�S	���͊}{q�Y�/|�W_�'��VJr�&u�6`��9��m�����Д�ro�4xҵb�����*!���YYk]8r͚5"<c���⋲�$fL�q�9�L�����<($�+��r��3��a��N�v�t���@����s+����'>�C���;l*�AW�;��[����])�{�[�ϲ2���u�#zL~HL�uC�E=Ę%��wѰ�N¥8��4��o�ӏ2����7���A�}���q�	l����>��z�p?�Fgcs �k$f]�8��G?������*�|����1g`Ro,1�[>��غ�4=m�To�a��zz-c�+3�'+�O`F�R[;�00�i�L�� n��@g�s)Q��m���CC����d��h��3W�
�y5^�d<2���49=���Uuu��eعC�
brx#�z,v&������n0j�,���d�:���D��X;;�is(v��Ⴎtr�&�iaK���8(�=�(�(��*sם�wɅ��l���IR.֪<m�kk������QQ���!�m�&Ƕ�=i<�-��*�����K�/��WYsG�[��BJ�ʣeN]����e�+"������\��JX�V9K���r*�➖@�^4�@�"�cE�O3iG�M��cu��xJpG �Iy�n��9kLA�)��T�;�?v}}��-�3�������\,N�v�k\9������� ǍvN"�R�4��Sa�@0�����{F=|g���d����� lޞ"SS7mڌ�ᑠ�/z
�t>����6�B.����ݘ'a��I8]v�y��=�1�D+#e
u�� ��nhl��y�#=&cE%�m�9ƹGhtd\e>�F���wi����b�ٱb�o���� J5��GD�u���n���w��RA���3�Q:=�S�r�R���j4ֆ�pj{�w܁��t�� �a_|�%ٸv.kJG��ܲ�|9�������>W(S�r��s�"Q��
�P����s��ݼy�O>)򽜃`FΣ�׏�}��D�O85�j����������8n٨�-=1��@����,Y�10�V�z��W�x �$��Z�Y�#��������_��tE�)�R�*R�s��R��+�1Ѷ���]tG@�|�-��GL[�y�n.�s�I9�E�����3G�gVP����"슴�F���>�K��Y��[�^~��I�vc{p�1�v�ڕ�dΤ��i�ڊ+�cO����g�rEe�x����.���7Y��U#�"j�)Cb$� G�ž�{Z[[�?�|4�k[��τ�]ؽL{���l_��z{��8Y0��L��\�ib��ml��7˖-s���2|gΜqRx.��/}	����|E
Yc�0�3��E`����s��r*k}��3�D2�b�TT�UM�r�ʧ�~�y��~����A>x�L#wg�����rr׮]˄sY��޳�Z�Õ��_(�108P�+��~��7|�O���V��ϝ7��j�wW�>��ǆ�j^x!���g?3�G�L/T�Jm���5��g�gX;O<�$8c��m���ã�4�6`A�=��[n��S2HNՔ�![4�씣%��P}��g��׻Qoi�ON���9TR�L�v2�]��3�)��b��"yX�zxd8�i[J����FMX��f�?�XqƎ��W�)p1��K�����z��c�����܊����Q9V�!+5a�<&���x~'�bT7�^, ����r+�v����L�S��u�1k�݇jEސFk$�SnE�W3trꩧrlYk�&�Wbl��O?ݻhؑ��H�����N�ʂ�k�1O����nW\x������:)�U4���R�h�yX������6�O�#r�RS�S޹�:-F�C�'"�&�a��J��'҆��9*eOz~���[�7U�\?�Qy����bUU2o����}jw����A�t>{ݺn�*�Y�h��ٳa���#�t�04)u�/��|q�¹<�W�i�Br�]��29H�%�Z�hPj�%�R��sø#��]��BIẔ��p��N�4œ�,�=^^�hh��]�y#�H���+�N�C��3���v�8㘌';3C��pjab
��xe� �Tں��J0���k%�ˑ�H��}���Ɂ�\��΢3"�ಳ���@�)�Y'_ �\_A̐�Ƞq�;�z�^%�O]}��w�y��W�R�w	���u��!�,����%|tt�Ed�/b���kAu����_gJ(������	�S5�C�
��0��(s�#*�ٜe�X�@�мPH7nd��\10	�==�D�V�ڬ-�+�����-�E@H�*�P)\%ec��^��d��_�����<�����e��80%Y��i������%��w�x�P�'>�I���Um��u������X��{����T���+P�<`_�u��!��|k�d�l��g�2 ���'����NVU�l��z�'@x��)`�����+3`��F��V����ʏ��,�+�l�ʊ���y�����ہ|�s���Ή��:��v���#G���V3�������o�}�� -t�(�w#��9�-���|����K.(��M�6+[�e��g?+b-�bӲL` ��K�G�����'���~�;�S>Լ�|h����O}�S�"����s�Y�,O��U�B�.\8�ӟ����˟y�m۶+��[�d1���'>��8/�O�.`8r5��ܖ�S�dp�"�����f�Z�{����M}VW����?���}�1�������r��>1�q�ͶaG���+/����������Y�������\�FGU�
��~�
��awN��{l���g�}6s�A���E�����%F���Ѐ�N��q��%3H[(4��6%�Tz{u����Sr �Vh1e����ڔ�*�]! �yk�0��Ju ,>?Y���Z��D)��"r�eMYg��FE�yRVA���nؓ��R1\�%�O*7ɔ)mǎuH�E����vԬ����A E���b�U� 2��l�zW?�VJZ���eGZ�C��,X���+��ʚ�p�MLel����.��ݤo���QH6Ap�b�4��/�~�G�C)�yNһz��&ǵN����8�p��_�hɭ�� �J,��q����R��ub4��3�U��8�����ЊrW�RwO+xe���;����u��-������F	[ʐ��rg$�Y�zh�޽�f�/ZHP
0�:����O�Ã��^xA���sE<yNYt2��|��b���+UT�S�J
һ�d����tZ���JrJm}a��,)����g ��d�jb����-m������;C�AP���*�bF��PGT#Xٷ������{�9��Q�k�
�&�Rr�+CS�R'AV�<r���Pi�	}綰�un��K/c�j����{�	!������R_����2L���V47ʀ𢡄p���g� ���3����X����䂈o�iy��"�<��Jn*��z4-�DƩ�}���E�8P�_qIun����_P���'W{����+����`&�o��";|�7���F�BT�|cq/?�[�>��SN	�e�5�h�.���6�\w���>�-�s�;��Q�S��X�ږ�\���[o�k����ߺ�O�m��u�]����]�CfT�l �`��:^~#^VM���߹/�JZ��@���>���9�|��2 ����3�\�b9:�Ø�Dc�9k:3�>��㹘����r��`���s��Z�[�����|���j�w��].���e�V�{GE^K�.+z�&����</��\\��d.UR�����ϻ
û̆��$Y�:e�����ׇhC�iT����Д���A���8���ZOL��^�0���E؟@m�����$iM�f |���RK����d��A�u�\�NyϞ=��u�h�C����=�]r��*����Rz���ʕ"�6p �c(����; ��9�o��y�����������eۈ����g��G�:5#�Cʯp�Z9�9VG�t��yS�ǀ���N���� u�Ó2 ��H���k��^���vw�2EIx�sU�� ��VV:��u����lB��H����Y��-M-��?"�cP�»�̊�N���^3�-�e��utu�㩧���W���`n��%�aG}�K_����@�]�Xe�H�pAv�����9*g�b��V+3.�{�2��������_�iK
�*u����+���$^Ӳ'�#hy��&v,@���؁EO�Ӎ�'������dqw0��%���T"'CR���TN�L��Y靓>yWQ���5���vŝ�"��~E���=�]�b�@���D�e����h<���x"���JMW�TC���U0�̂�8m��#�CV y��hS��
��S����i��Y��X�bEss��c�r��W�,
Q��2���^P9vkkS��G�����w�+�|������B{�]�ŨJ�1��9#uu5�M �=���E�\z�DR�?�M^�B����DX���<�\ĳ�N�1�C�A���i����h$e�A�X��&�1j����P"�də;����X�E�kh��%�JTV'��1��C��uy�K��V�zDO/]%�_S$� ����H�8:6��y�����׹<�JN�ș3g~}}ӎ;�˖�Y�M�G�G*S�hDy]`;dS��@�˿�[Ǒ#�mm��ӳ����嗊+�vA� ��ηW����{�54Y)�D&�֞���x��������.���~�׿�u�]���s�t:wD����}�ҥ��g���Tl��M����曹#2�ߑ�V�b�z/�l���#X���ESb)�5�_߃�A1-
��E�@�(��e��W��7��T��JAQ�^ٔ��B�[;��N%Bi)�6`n���(�X�e�>fbQ�� �}��3�#����"V�I8�Ә���\+��1��,Xȉ�Vno��e�kS���_ޅ^ę|�G�:��Qa�y�y�
�Xp����Wl� ���k֬�c�%�D��B�{��u��������E�i�y@���� Ѝ!��믿ލ����"���=�m
��̊��3f�J&+,8�	cL�гJXh��˥�3�*�$wa�N9u��'HmeeEg�1f<Q�6#ܡ��=�E-�����f�s�(���c�,s���vCV(.�)�)?4����;���<�f:�o_}cc"����	��Xg���x����1	�.^��O�*sK�O�����>��챶)�
)�7��a��=V���1}���X��c�c�V����=`B��x�K|���,��4������L�"����LU�V��A���f����cC=v�X++�����O ��.��MVT�N䌌E3�L>��47I*���:�M����&��YX�fe1���6+�����*���-�o	���A$�LU��M��=212jL��f�ic��
G��Hs���%�U�Jk}c~<�90(�z�������U���pl]����:��tnl���H���f���Vk�2l�Eb	��PM]Ue��>lnmD�"s �h;~�IiC+��jj��ǎ5�`i�s��qC%$�
c昋���i],���omn�'�J�hlhl|ĵ�x�X�tj�6���x}cC&���:�rϞ=�g��y���.U0�\���
��H1(!��XP􌗰�R�|�X4��G��t�[�[M���0��3u/Y�H�B��5��%b��G;Z[���4�c�8}��d�b�Yg��ÿz�(�GFgL���,���wN����rp���mK���
��'���(%�'��R�� t$�v^��>W o��(��<��	͘?��jV.�<�����'�V�1*��\+TTV�>��|��+ĚZ[l�������j��"�$x�d'jj����BVM'�=}ǧL�261�m��Te2��UT&Z�s�U�3s��LG��h��h�����ʸ����Mo��}�`Ҋ�wn$�^\ŶQ�9PF<�P]�{�ǧLm���O��u�	���uΌ�%��9����HMm���V&�L.�PBv�rd��7U*��"T������Lflt�PTVWW���Q,jRvb̄X*������|&�v�v,_�3{����2�l��Nd#�[;Q�
���)D��|A�B�p|r0;�{�P��]^Lȿ��-� rd���J%�9c.���� ���X��h�z|X� �[��<���/~Z�{؎�<4|�;�D1����N�>j��0�^s�A2��n�
No�>CK�?D�(ʖ�'�"�7l� �Q�Z��B�kyd�+�:�k��ץ�^j���z�%�p�t���nQ"�	�l�>���(s���1���ίh���l>Џ�+���+}�&.(Q���Y�l�I�aI�	HR�W���cZ�e�	��cJ�f��b���+����m�s��b�'�y�w�q"�%�P|�'�>Q�xt<x]5k�lm3e�/�G�/�첶�֝;wɐ��iAL|�Q���#K�t{���;��g�g�9�b���S�疯+�Z���B��EBa��]v5wy�ט�D�b��vhh�T�ӣ=��aA�\\>!�ǖ���Q'ٗCW���G�.�\�h��O���ʔ�$�:Mn��#9�YYF�CYew���ep{i��j^ek-��H=[B8[%�,(f�`+62q�Ok]��f?qܑ��<�����:�ʪu�s�����]���� ��
bd �I��v�x�u̘��j���Ϙ��'*���|Q=�xKse�-U���a��qU��TT�_��-L"eҺW����wʂ�|ݬ�rc�Cp��ya�R8BZ���qc����@0�S��L���JQ|�V�텓��zW�,��[wxD}�?��`x<W���I���f1���3ϰ�Ų����,�ŽH�ޞ��&��*?A�U�O<�1�&�*�V�>í	Ӹ��W�n��	ӫ�\�p��~S�V��0�P�&���ɤ���������I����9�,Ye;q�3�	g,�Y[[��o��A1n8�$�ųϝ3��۾m���g͜%�1�NvY�����
_����y�-R�D}�s)D�xѲ?&������D��	�Z�b�n�E�С����y�+�C�
�-(��KJ�*�`��c�ΝU^t/�>��gVvڴ�l�v��k:~����
tx(i���گ�>?o������XN,���Q�^S��de�<s�����(��)�[QE�θ�uJ��N:�
MP��X!$�]�-O��o��Go�JR�y�0���c�%�y��'���
qNv�'��/s�_�4u�eT!��Q��Av�g��{��խّe[�%ٲ,�C��rr�8�P8@�B�R�"E]r��ʹT(\@UB
BCH !��!�y�l˒-k��s��=�����Zn�p���{������;>vnjr�Z(`J�������.�������L�\D�	��Ս�U�5goo7V6�5���)X*�I�j#��p	�5#�M#,��V%ϙr��p�2�3WO�M6���Ba����X�(�����p��|hܧ�z���T��6<���	'�� ����At�M���@$�Yl.�wg@_��){���s)��'��07៨s�J"�-����H5�`]�b��#�y������0�G�Ԉ��Y[�쪉�����)/��&��C�OT���bM��f�4������\�9��i���p����qM���ڢ
����ru!J0��^3=m�9^jک�Yڦ��5�R^]�.�l�	D��E�̒���W�:�|�{�egl�u��)�Bl�F4��Xf�1��Ql1`Jwժ��?������E�u1j�#*֧�i�J4��w��������IħAB-/k��n|NK@��/�Kڋ�{r���7�l��"��m��`�%�jxX��\��w�IRn5�#kPu�SX;�������tf���·b���Ψ�.��rIh}
��XنA��!�ɋ��iN���>dN<�6�Hgv"�<K���
�|8n�R��� ;�(FM�ڡez���b��D�W������kn�햣GOJE�V��!�|�|J鷘u��V�nX/{�*Z^����TNS�eYB�Vh���
�ك�ù�bS%g���z��7��|~o�8kצ3>�rD_ڤ��*��e���+*F3�h̏mk��U����)f�%l`��MM,��i�I�e��(��:�-V�R�%u���:��u 蓅�u���8��Q1�5���lkP�e��}��{�G������O�Ln�%�_i�V��)OA��뢎T��'�k���R����r�R_j��7��rF���w2�,��K��Wl��;��cY�N��+xpD�{Njmǎ)��K!3(C��FqR±`Q�7RG� L���a��7�DE����G�	�en�W!HTd9�ev�����lK�P�+"4P��f0�%��S9��W߱��:B�r�c5��`%ǰG��|��b�K�Ŷ�+ŀ��/#�۱ϊ��S,��d�޺�:��W�:]��P�ÖXm8K�X�AP	����	�����RQ�PQ�J��I��J(�	V��'���6���Zq�I�i�tķ�4���tif��>��c�	��7��	�c	�A��裏bHq�)�BT��K[e��O�夎�
�y�ԩ�z�đ\)/Xۚy$��"�&��0�o��md�����6ɖ�c&*��m�f�6�uk�>��b��
S$4���5���,f���u�� ��fBM���qd6ONجO<���3���M���
9���̹a3�y���I�l܋�=��������jl����LlbϨ��/3��v�WrC� &����(�Q�6�a v_ �����DZ����^��X1�=휣�g�4W� s��ɍ��t��9�52������Ѵri�1�'�N;7(1�:�x���o�K˾�����^7
ŋ�j��l��rme�	�g"�a�'��Դ1B���$���~����.OsV��xy�h
�Q|�{[d1 ��t�B���Ī���(��i��K6��[����R�p�`x�adD�ʊ����,����Iέ|����P%�K��mDa[��LӪ�5�I����̒�+��'Y��ʏ���C'��W�x��ߍp8��k�%G�aW�:80hphtt�$]^���(��qR��[��i����Y������F�Cg�:=��B�3V�����!hav6ըb,�?�U��@<���o�^�:9p۽d��=�Ο�M��+��z��q4������\�t�&�V�s�'���c;Yĺ4��_:.԰o��}��{�q���Y��5&C�W	q�F�v���A�,�|sҖ<¥筵�
��l�?�ط�z+�
�+�Z���I�F�5`�wP�y��$�8p!4%�ZZ�V� �s~ m �y} 5�,�&���|۽�_K�<�l$�E������g��Y�/�,�;'��������
d�U��F���q��3�daa��]C���>�B��vJ���z�aͼeoHPҼ�a����TZ��'u�jG���Kl.�T.Zmtl}n��W_y�G�N�b��ơ�.�x�>�[���e��&5��:���5�XWOT>/&>D7[0�WP9�uI���nf7I��ٹ�T�]W-�v�\���V�ϔ�={h��XT�$�ZR��ӎL��%�	��/����<�q�RP�9f�����[忺����fο���y�j+.0
Ⱦ��l8�ySv�����oy�ma4�Q�mig9
J�Ҋ6���
�~����y��4�Ħ��ڽ{�ʆs�D�]a��
�>}�70����y>�Ԑ@nR0�r��#���"*�qC/�p̔�ዖpr���O��yd�J�d�3�<c�1se�
�@�3n��#b�@�&a��Ӊbj��T��ӉpZP�6�h'@�dq��ـ� ���xh��W��B�:*-=6��ɭ��$#Г�s�;3:�̘�p*r�ޘ��^#%Z ���9��O�Y1����=gJ�L�A�����0?�>v�����X��[.}��֮Y�h��ʒ�6�>ǦR�Xxh��k[i�[�� #@ZryE�dn5mS
~>��u�zj]��Tv�Z��(!n`�D2W���t_���+��ֺ���c0����r�>7����5V 23�h�F1���/:c�:\�ML����]���,�F#�fF�m�uj�I:�/4l�T��i/�ڎ��.m�(���YT�u�փZFggU���$�_��k���ѡW_}�_.�������{��U�vٞ+�h}�����o�Y�]��<�a���HL�:�D��ܴ�!�x�1yYyO���<OZ�i���&߮��drx�{���eDY����'��`�}�Җ),ش�jb~�+��r��?�K��YZgW\��#�U���LZ5�����(��w�hV�ʬ�J�̼LF'��F���(�T��1����r��=>i[�Z��=�5��j%B�Iq���n���b��~W1�mII
YV���Nc�
E�H6��M����7�y�u�=򘼚���]�N�����͆ƣ�ϩ�[Ѯ ��M566���}�=�:�̨���ٹđ�gϓlrO��S��iՄ��������W_}��� �)�r������Rxx͢z��/�:�~�9?���ek����(����ߞ1����%��
S��]hݿ�>�ָ�(����,~��e+��#������ĩ�����l�),���SVz'sF��Rj� S��1N.������N�'�ۭ�><j[�˵���L�@�N�@�6������#h)�K����m��_�e���oG�!3�"�L���k�I��fS;�55(cz,�e`<˱Y�aHL)ߒj�ք���G5�L̸ۡ��\�z��e%�KVԎyC���`��Uc��`���YZ#-��mٲE&a����O�����>OId�<��
�̃O@�D��ì�`�Z�U5���\�6Gq'�o�T��t��*.{��g%g��J>���U�h�m޼9����B����`*�-��G���l{��k��a`k�(�a9���Z�K�l+����.#鉆<Z?�Р#�6�*\� ?���, _�f�x�'��ȐL!�q��D���Q��=#���u�S��1����(D5e�X�4�f�+�,�क़ن��<����uht������Ӿ�툭�⭬����4�� �n�TIU�l�zə���3d=|&J��Yf�;c��;Y��e�?���?Ϝ�ݷ��{m.�l�[HS[31�D$/�3�n׮]<Ũ�ǜ;��M�������F�V�H�ZX�	�P�b�U/U�y+W�4f �G���b`}\9Z|*N����|ǎ����$����Ca���FCj*\������V�����FvYG�g8MS^�ǔ��PQ��-e��2�Y��իG����C;'䁱B��{K�i�=�Ը)e��=6����.\� ��3��~Ɩ t����<��ݬ���k����O�`���H���,���e�o���z��2{���-�i�z`�3��u����Սk��do�-��i��\��e<���������L������U_�\��VMb?�rV����z��%�����}�����w����Q*�p`j���|��f��X%]��L�;\��o?�qy�e\1p���W��:��������߿�[�r��8�>��W��U���Q7&�r73�r&tw�Y����&�-J5�ەц3���������$k�9I��c)F(#�Lg���/������g-KB�g��8k��!��Z��`tx���D7\_��+�+�7_z��ϟ�Tk�6��J�j	�n>fˌ�!���R}�F��3�,��_.�D�?�vV���®m	�~m���35|	i>��(�rOi�����e �Fs�6-���aZ�%ڔq����nE����ggٝ��[�ƄD�nY��HL
�Ca$+�t�:@�Y~P��v��	�)�-�6$PU�
Iֱ6�跢£��R\�3�d-6���i����v2�!�\�K]e<O���D��� Ԕھ,��^W+�䕑�)8�\k�=�~<$�yJwt��m5BY^�;��m�����;wCQ��/����y�~��T�Az9�h �'p��cE����X���/�QZ�"���¹�3�aFoc�����\�L2>pO$���#GNJ@�C�m�nc�Z�̱����i!O�YxӠ���G��K�Hr��r���=,�����N��A�k�qK��v0�psM�޾n.�X��L{	m���YTD*��U�(d]�t|��m�%��X1<:��S�2T�s^B{a�5���!��{�x�'%�����ޔI����JjAc�]e`��i�W�u���DG�Ju�w���1I����+��[ą�{�9�*�z�NN>gO�(i��ls��ŷ�z�-Rr�'�|���~�~�[n���~������;3o�����y��#G��i�:uB{�Q�=7�/�;��k�,ېے�>��46�)6�4�E�X�4fF���]\�/dt�߾{)�=���y��N���jk,òP7�&[E�z9�Υ�cѧv_��������\���*�R��^X���I�^�v;�-[!+z�]�2�+kX㛅f 4Ŵ�U��%=їLQ!�go�گCC+�`��T����}߭����U�e��:0��F����m���?%��'�!�[f�uO���c����׾���o�>.۶m3�Z�:ۥ���V�]������gϦ���o�Y&�-Aެ5ףC�����G?��h�c�|���B
�s*=/�(m�ti�4[�Hm������(-~��*I��
����	�1п��'UYI�[:Uwx��[��?NN�R� ��\o2�ڥ7�g.F�.���[��17[�l����{J黨�S����v�W.U�D�7��®;�U͋<����ޘkv ���q��g�B�@�1�lw���\���DB�a��qك�2/X��+�Ec�
,�Ou	�W���+|������&�����.��O\�V9c�Z����X�ۨ�4�:ɲDYڕG��M3I�dҖ߹��Y�����lc?�D)L���U��i� &LD���"UY�Uw�J��!�X���E,�3.�>K���L�7�LaqEM�0'@��8k�j^p�Dq�}�*�*n&�Q�b��V$�����+xx�F;��eӸgxqA���x�� Z�r��<b�gө_|1_ᘰ��Ce.���ѡ2U��"z���l�![3�L���bj5{��2� �`2ټlӭŞ�Mg��-d	n9�;���9a���~p.Mx#Fn�V�5��ػll-��Jk������j��`y�Ɛ R�&�!A8�T�[�V�����i�V$d��L!����?��OG���2#�l	]3 6EЗ����d!��;�f��}�޹�a�ː|�Z�D3%�6����h!����lv��;��<v���]�
O����^{CwH�.5S�PY8����T�|a��qOt�믿��O�u��g�&�m/�N�'M�ܬ�ZCCɬ��ވ��d���G�^���v��M����J��ף˭��7n\�o_��������\�?�(��3TPn������'�H�`;�Ϫs��8�"���<�0ߟ��᫮����AܫK.���}����wx��yde����HX{	R����R����N:�J�M1#��s��i".�twR��l�o�\��������?��w�4�h�kd �$�jO��JP���ׯ_{�\���n���g�
����2�}NUW�Ҷ�?WF� %�̓)�o||��T��`��q��d�aO�D6��F}������G�.�R�Hf�S��ۿ}�]w"�g�2��F!C�-5��wog4��N+Ȇ~�\�_%C9�@��%#��l�xa��&o�T������T����ޱ��5f?�j=�]�r��\l��z�gfO�8�u������sg��˴�ji��0�9l�5���sM]�D6�a�[��><�)��u�V7��T�/�P�����M?})W��j{�d8F�k28�����w��zc���U�֭�nиd��
�{2B���/2-��T�o�r��fWY�Lb�E�R�3����&�O��&����ym�b�t��x�T����eB���h�	�C��r��a�'Y)�
���MF���k=뚠'~��m̲}0��
e+B<�,.��75��8 ��v��C7�D�;8�b(ۍ��tsK!kX��R�m
��cMyA-NSi֥�'m�Wu��|�pr�b�H��{�oYgZ
�ks�
D+
�]�� ����(|�����k��;w�Yo�D�Q
xb%�e�[Y\��lG���Xl����6*��-3�����j;���rs��5�dv�j����*F"Q�2�nw�k�����+�7��|T�P�3�Q}�ӳ�-k4k;�c�ےI� ��ۖ��Q��蚡Q�chP�^J�^�Y���m611~��	��
Vqܖ}����4�}L��0Ӝ�w��ˍ�Dm�d�avJ%�]/�)�fma>u���I���,�aY�����xꩧ4�}L�V�0x���d۶m,=�c�������[䎿:���Ȣ{�GĈ�W�&O፶^��eݻw��Ȫg��1����Or_KQ��M�I[ (���qC���B��d��f�-��˧�OԻ�
Q�$޷�u��y��,.��j:U�zA]IOau5tƖVŊM,�6���f��!K��n�%�\£edo0>�[1��u��u9���D��4��̟={��ʴ��e�pu�g~�k,���"���C�ìȉc�y�����ɩɾ޾��I�2���u(U��i,�{�{n�9���a>JLN�؁�%*�ӧ�ٵ�_��>�O���ʫ
�b������G[�1Y�j�tv�0�/�/���}��ݻ���Q@����Ξd��4&� ���+ͻ��������:�+��L\k�֮]����E`ɧ�?e{#ՋQsj#2�,ޠ��]��T.�-���S?�SX2NWo���S��
}���#P����	���Zj��f�u�+���ι@�a�_�J��j ����n4��v
�a�"��1��)��I)��nM��c���4!iTD۰�jaRо�bڍf;"L��|~n�j��RWR핵v�3a!և��2cWY���f�=�7�4�#\��SN�<e�SF[�(ӂ�/D�]��&��Ĳ�tb��\����uY�W~L��� �<E��Yb�b���ʵv�]U�5R��
o�V���7���Ͳ�mn~�,�j̈��;��f���sϱ]��:�ҵcT�G�+���2�#U\���$BpK����E���<WA��qm%죏>j�}��!i3Aq0�(�ת��a$&�NGsR�lw��R֖Z�oͬ�F#H1�Y����N�7m)�S�,1<�~�+й�d�0�)`C3'#%Ѡ\�<pD�c�by4�d0�ܺZw� ,���Ohh�h�h2xKx�|��&W�8�e�GϮ�G4+* ��T�o��J����H��:����(e5J�Kp��\[md2��^z�&�9k��}˪a��p3�m�	� C0w��gV�9�Ə��7��ک<�u�Bt� M�Z��gF��3�V=��iˊ��B]��*
q�d�+.��T]_4�Vķ.lঌ�47�l���y)^���u6��BK�ǡa_Y�^�+)D�[���/���C_}ƚ���0��N������O~��'�|��Ĺ��N�6�h�X�Դ�h媲��[o��?�c�U�yU�Y��g���$S1F�]��&E(��Rs+S<on6/�A�9r�����a쎮Zu:j�Szwr������!+��u�ק���G*r2�^8���
�������@�f"���й�B6��RMQ���;��]�@}h(u����?���|�/��Nig(f�AC���4��s�S'O��T���+�$K2��L
�`��]�נ�%�^z��fl��5i�'n���	E]�B�>:���6m�Ї>�$���g�1�`$��Z�{>y��[�q�]w�[6m����1v���ėK���(u�O���'Đ�ݜK힖�7����טq~ �����Sm�k�]��Ҽ�g>����3�i-`ؔSX��}?�s?�����e���݁E4���M�� ���gΞ��_������ں�
���̚S5��<#��F�r:*P��PyU�b�`����K��a�h�����i�����&�������R��l�R�����ӗd�����,W�E��{|3����c�����i^\�<�g�k�?1lܠ��S	V����ˋ������#�n�$�²r(GZ�����n�cԋ!4�ttډx�;�l���ؐ���Tf)��ER�6\�z�����N�y�R���Hm#�,����N���*JyC����z����>��lB&�"�vC�M4��ɂ!e�Ӕ��^D�4L����0�e-��I��-)Q�*���7�^�OABW�UW)��'8fw��#A�E��#i���=���4�����&TS0��˶Z[��+%��)�+|�Mx���T�� n0�p���񏻢=@�����k1�$H�>޷/z��Ҿ ms��s�%��(�9 �r��g�Hj�e����K�=�kK��جֶ�Qma�/:=��2�1�5+��0��+�=�z�������d����
��B�#�?�ǀ�᫯������[�sN�ڵk"V�R`"ezã+d�2E�&�}<�	YH(g7�j4�"���ܘ��a͞�-�U+Awm}%��[͕�Қ�������t�fhq�nDVЛE�լ/^N��[���C��&�˶���w+x�G�d],�z�4;�l��@�%�*D��n����Y�볡�Y���?2˱�����\��1�ѩIϡ��M�I�'�#EA���o�~�m�}���3��;˳����֨���ICMKz������s��I7=�����~��$����G0�։�)�#N�L�w68�S>�ܹ�k�p��Ty���1y�x>��ؐ��h)��LMO�w�f�K�d�h�3�)���f�F�@�|���le��=�)��
�"�#y}�@������ӷo��u�gx�w��]���>�D1�uA�"9�.�������+��"�W�D��7F�?�j'=�D���ߺu�c�>��s!dV�!�:�<&S�qp�r��CY�LjN`��u���+R3E%��*���8Y�<���26v3��ǘ��y�k���U�A�v� �~w�<�T~f���)~�~�7~�7FF��k0�0��.��g��������_��_Y�0?JNS�ŌuEE,�*3����_�4�066.��V�74��ʺ�jؙ�̅@����n�Ms�8��KJ3q�U�	j2>1.�O:��f�]��..�<,K�r�$Ьy�1�y��g�D~��K��}�a�C#&c�w��؝�>Ӛ>rIV����݌:�2���ֶE�{4D{��ZMQH"{d�ք��E�YO*Z+q5[�d�9of��y\��g��s���E�V31~�x��?j���;�ˊ�kew�I�|�ܔS��y5��)-'�O��ģ�0U�I��C���t�&e.��	È��^S��`�I�/���y"O�ǌac�4sO�W ������FPr�o�����ы�b-$�w�}�Y9a�ģb�C����5a�V)6�3o,�d%Y���Fyb�D��2�?Ջ�
SC�@��r'�Cyee)�u�?�)X=:j\�W�
�G��V����d(�������GS�bFcB�xŨN�Y<䚡ķ��{�k�Ϊo����� 7T�r;}�� W~Κ�/o�0n>�
A-�r�מq3J[��B�Ⱥ� s>��0�ma�$8l�l-�n�Æ����s�
G=�X7�5�Y	��FD�Bf4rj�'U�.,���'*�ft�4g����%w>7�е���Y
`s'�J.���^���Z�	e�CR:+'-=��BӴz�{�I�+��Tut�����-r�V	|,PU��RT�a���wfR��|���|��_}�Gd��'0�,����G�5;����>w�7����<T��᱾QY��~�[�t����qM}����t�������gn��f-6$ ���8l��;wJ%��O~�={����������Ȋh��2�������G�FYh����æ�L7�ŊYd�4n�ˆ����

�K/���ݰa�;ν�~�+Gq�Đڶm[8<�� �8z�x�y�yA� �� �L6���k����G��s��o�N��S��e����_��8����p��mq���-�,_��^o2̫vleT���S_hX��"�hL#q�Y��Ī(��2�Ss �{LFGW��/�1�jMc�|4��M7���o~�K_�z��T�'bx:ۖ�7�����_��_��'.�璟i�&�n�#���$|خ[�\�/|��>��/��;GfL�;��|��D[!����62��������-����?������ a��XD�'�e������_��/�eȴ(Jx[-�'^`����Śaxi*b�2��ZWb�Z��.�����sӯ�������.��٫/��?�n�j͚ս�����Rj������uJ,5����DScA�.��?KE̬�HMUr�h��g�-��M�4��V�Q�*$��Ԛ����5.-�L���B�x(zi�TM��mbK�]xt1��:�$u��e��;�]?B�r�AZ�i
�c0�S����9c ��W��B�N��xb"7�������lݺu.�^A�h�UBk=�n\�9(QӠf��ݶ�(����w�^���-[��9qZ<D_oOc�5П���ބ�Z9<Z��$�R^���X��;�-EY���ņ��\c)��J<��SH�7B2ūjI[�b��p+f�M�$���3�FהR׼Ti�˥�K7П�������c������"_71���Y������٦�m�e��'j/Dw��gw�b��vڱ��T;� �P-K��ad��{�o��+�.�`�Q���ƙ`s]CtFR��ё����7c
��ɰ�؉��d�񦎓!�8P"F
��ھ};Ύ���X�-���L�5z;�<���4�+FF��'�'���xj.O ���q���~�C\�ү�GO^�Bl�a$�9;핅�b�c"�L7I�����:R?��$=׸tu<���!L�����f\|h
��/2�:H�L��c{�-onu�u�I	a��}�c���˿��o����	�65��r�y��J�� ��JuӦM������8�p�2�;��ys�	����,C0�)31�)�=�������s�Թ�1N��J��T����$�gƳaC"o;x���:�1fͶm[&&�?��3�v��u��ظ�T�ҷ�':_��'�䚦����s�nLN]x�6�Z��6�Z�y�����/���RI*��|�L^�Ž/��9��+�=�wǎm��O3� ,�s�j�`㥘��j���S��-[�Ѿϕy|���ҝH���P�r��Y3�˃FDX�a~�A�Q���}�𕫬]��ⴤ��x�̮�їS�*����/R%��]	�k�.�ucw�y�4.�~��1�ϟ�4$d�&,f�C�y�E�����g9�v����v�����k�g=���c�cm��آ�_�g�g���*^Q���۳���R�mݣv�-/H�B�@�`�H�Dkg|ua٧,��l=5�]>��k��gt~���x��F`���Δ�'�l%lIj���vO���$�O�9�AZ�4K��d�-���5P�#e��`0�fe����\��3��hA;��h���ݙ8��Y0�Ī̇62ʮX���i��k�)(��X�'b�B�/�(��Y��1i�ȚÈN=x�o����*�$��>+E}�%xuU�ըX���U��ٕM��-pcx�G�/�U8'��e�<1�&b�gS_�՝G�J;Y����k�c���3g�U�ؼ�%|���
q��PP�����=V��	q1�#�-��2�頤KU������X,�N��`K�T~����sbz���[��z���A_#�� ����<Z�Z����O�(~n����3B��s�ݼӏ/������Y��_�ؼ�1rc� nn-��z~��֚��L����R��2o�_��ȣ�³x�@�T��W�_k@�	�N�C%ޯ ̪]�Zʪ-�Y[�����be�X���� �2H`OX�v�*�evR��v�hS
���-y�l��jk����J�b@��d��s�=�fwa��v����T5��7�m��ķ�n�}�:�NZ�r'D����?�u�)!��{��I�`�$�H��U5�0�"�����gAQ�3M�,n6Rm�@��H'����
��V:�<�"�ܥ�[+YO&a1cy�2w�]�v�L�w]{����82�c�QC?�ʞ�n��wd6n��V�`����/����n{���n������jel���v���'�a>���L�'��x���ׯF�Y���nݚF#nH�8>g���ՠ[��\�*��X�D�z��p!�IE/��s2�(��K�KKo�y�ԩ���I&���l
����I����W�3�|W��r���U�?-<Q��TH�� ���'dm9�I�x��HՔص�)�T-W��� ��Y32__�w�\�f�m��b�c���<��(�m�US^��B���W5�^͚�-��mo���;��ĉ�����c�kG�A:,{�W̺RXIyñ���y��X��'�T�y�ęH����O���w��}��9e��3�2~1���h�OI+>3�4�{1���S�|^'�V̺��yL͒�]�f�5�z)q�е�ԕ3B������L	_�Pn���67b��f�1�T�@���k4��ӵ�ޡ#���.�>q�;Z:$����vF�=9
AR+k s�J��f
�a�&�H�B5�3�b�ŷ��6*&�5%7_�$��:9��b�C/V�Z�e��;c��Y|>r+�YdN��Q3�uz��Ub�e�PJZ����I����a�BC��y�� �[a�F�̆�OQ�XF� ��3Ԏ:v��N3/�y�f��,+E�����хV�J� ���8*i�|����D���|�ۚk�t�Hy[5���Q477Oʑ+#�y"�h�9M�7�o�a��Q���?���I2�(��k�*c`����q��a��(DO��z��,����i�//�[,�\ȳAD�/��D�+E��d�_0��]ѶA��9D�����������O�yOwQ��� q���}�!w`�,��+�'��1�Ӭ����@i�=FUYA+�5<�L�֭[׭]������
�|k�`\����hhU��m�`p5��=��0��r�2�v�W��-���bT���K��Yl�<�������:P#:R!3�h�Tx���iqc�f���܇�t0��yhr	S;�.us�v�dZ�` L�=Eyk��N���l[ɋ��B�&�ͺWi�<�����5�í�j��Z�m�6��;�0��ٮH?[��?��8?���6tH��g(��d��Txd�$�+WJ-iՋּ��5R[���*�_A�b�3~M�U�FT�z����/���f,���G��%��w|g~6o�t��qԂ��M¦�<4��]4`ւ�2���%]Eى��&�;q�ȕC���l�%�Ղ�� cad'�% JyXH	�T�ɲa��0�ј��Q��J
���k''g��;����LOLbJ�L�:Bn{�urff��[�j4vZ���1M�jWي������Z6��-Z��K����5�UU�6�k��H��G(0:q��!�1����Z�w�K<��7lXW�/����O����Vd�JT�8M�����B�0����~�5|��b�1�>�L��d�L��A)�����,h3����V��1��V������9��J1��ө<;3�n-
+ʓ$�J�mc~3ق�j�ͦ�G��TQ9ۥ�^���{i�`b���W�����b��_�^B2�ֺjŵ� �!�jll|�޽�F7Ō��8.�L�\��Q�K���':ǔ���)&�����dLO)kXԫ��Jś�B�͚��KB&Y'�+m�W^yE���O̜�2�Ԉ������0]s�5bM��7�)?�� k4˺��L���D11����B�$/D����8��v�9d�$b�r���}��[1g�� Q�F�RԤo,���r���Ж���O4s�|�I#v��w�9bZ}{e� cZ!�NXc���|U/gϞ=�d.���1Z���
\�SZ5�pbQ� "L�'>��'�3��-n'c�Ɠ��l�0�G1�RN�A�/K�0pe��P\�����i��gܰR���F9Cb��~EQ����|�?1MX���C�����y�v�r��,Vُ%N6,2䠎1i���������-b���R�	oڹs'�g�Bhf�R���k��T�y��p1���l�z��Ijz�%)��w�;������n2�̓8����X���cfͪ���ɨ�N��c���y�H;f�M=�xC��R�r��Է���N����K`��;���)�hv���0;-6�f��~��	��KJ&�N�P��n�9k8JB��e*7t�E�2?�tʲp)ʚr[����u�6�:�f,b��c�D���e��a`	��PN���p+I[��(�F1��Wf�d�S�!f�So�(]4����+�������[��5o����=�?=�f�x.�EёK.399/��*��x���V�)��Z�����+��v�0vA�b$�b3�(�`�j�f#yG�]ƷXĹzR�,�	���l7m�83�`m��<X|��C�T�d��!��$�g��;���~���<�tTe23��RT�ٳ�B��v�$�BJk�D$���P��e�V�S�pCq:��Sd��kι	M���-s�H2�bE�L�s��q���Ex�9j��n3E`t��v�Ŭ!�蔉����j'YU���$f��������l�lx��o��H�^�y��b�+߸��VQ�cAMLL7�[�(Qt���c�,�h�V#����VpD$���ՀS�7R9Q������X�o��o�g���6�(���������m��S���^\,���uo�xCϲ�s�ǆ�V���狓#�V=v��J�I&C��L���o��,�ș�yc`_S/�2u���4�R����@��z�tO�+�l6Z��N�c̢n޼� rcק��,}�hO�g��G]˷���w�3�^?�6���Ͷv�e��#)X2/�Ǫ@���������E3�W^y%��g���ӎ��=�ӎ��zhrj"�Hk5��Ņ�	jbr�;h���7�E���C\R1g9הeTf��m��;�0��>�����bT��n��b��޽[(��U�gT̆!-�Ĭ�k�����߰�z�g<Q��>��np9"�q��C	���U(�%�;c�V�6�]�@��6�Ih�i&Y˾�YA|6kG�m+hM�W��l;r�/Y�62�`�(��[�:EC=}�zV�=u�D:�݉��\8s:E�ϝ�М?�Z�F��1�P�)V�ϏO���#ǅ'A�4ԉW�� d$��͠rU�od�Tg�Y`�ڃ>��1Ag��f�����Z���c-69���|���V퉮)N_X�<��}`rf�9ׇ�9�8*k愅u�P�s��U���-�:2�L��z[�y��0�;�����������R.����l�����8u��Hϗ^�P��>����31��UI����ߓ�(_����n�O�3�:�B/��uk��VIx���ɕ+ml��(�{zz�Q�:6�'�ؤ@��6]��`>� @�hQ�3�x\�o`]�@^�{Z�jS���8�b��������C+6n�����Ddsn�>24�b`pf2��]+Ѯ���qBt����Ac�����P�.�
ыma�����t$�mX�n>|�C�~Օ��cG��q�Q|vڕ;���U�=�/I�/���du��lذ�رSb1�o�>�2!^M%��L2C{�Trr�F�-o�q������#:u6D�^���C�!*#ɥ_>���U�+�ks���]�izzF][H�~�!��r":C�z���".�s��.�\�2�����ĿGsNL%o}q��}���)>=ߊ>�e�T{���\���
G��Z)����q��9�ݵ����v�Q)���\<3~.�����)�VIA���Vm6SȪ�P��p~2q�!E�?�IE_�-9��֮=p�}�^����bgN�L���4��$+�������(��uU�Ų>�5��,�
k�F�}.��D�n6*xRy��ъg&�q�g
���Z��z!䱫B�a�����]_R���e��ٹi<)<䄡,��������ɚ��i���ϙ�E�'r�b���877/n��S�:z;u:��Q�=�ƚ�F��PK�5�S3�gΜ�.�ϭZ=:5>��&l,���j��l,��Ņ�-�[`�����s�+�#�a���rAF�RFc��J{I�
��6��{.ɻ.��F�%�*D���e)׎�nSل�Z�bX�o��3��QG���w9u��&���Y(��l+fy��\4	���	���r$�G���D����@�)j��T�Q�H����mSQ�#�-Af+ŀ�NB�
��-��q::;w�4�g�nb�\V,<B�Fb�#ar,��n��&�=���,��v�D�{0Ϧa��6��5ܰ+�軣�h?rޚq2�J42���܍�0f��;�&��ټ�P>�J�7Z"�h*8��/�5%��8E�$���^x�1�{ｶa�W*&��
�)
����b���!�����k��>�ʄ.90�̰��Ŋ�g�w����T���;���ʛ�LQ�u뢃G_�����MQy�R��=��Ԉ�R���YR[jDи�%rܜ_؊���#�\�=��g5�R�v䠱J�F�)��0�|��1�.�� "M��<yG�w�^-VЖ�uĐ��|�4��I�b�sݺ5���"�p�������4�� �]4�<;�}�{�g=�%|(ɧ�L�:at��_�<�rXl�0��4��vS/�8?뺹�΍��;e��� ���Z�vm��y�I�Wv	e�0>,��].�g̬�E[��p�=��hgm������-��n0��=�����cB��/^�tWL�v��ї�ϴ;#�,"3�a�B���QL�s��mq+�)��ĉ3f9���o�Q�,\��L �j�;��c�3���j�;�	�Lժ	e�W�F���|]���9���G;F��Rc�\��q-)�%qX�TkM��'\؄�Ӌaa�����TȄ�B�0��N�2��Ʊ����{�H�	����[��t�ik�eMC�X������-ց��7���S��	��rM�m��؄amtRi��<��=�E�F��O��_�=#�j"}�-�ef$�)�)52�c؅ \?~Ҥ�)B�Z����L��?-�� ie}Zߴ[r�&�� ���sܡ���l�Mw�WFۛ;�����9Mu:��7�#D{�U=0���-�W&����фxn-��,p���O%{մ�J���)��hu:�'��b�Y�����v�Z��9`l�~E�gDF)�.����z���+����ĥ����"�k]=�Ύ����ˋ������F|��_
�UjgN�[5�f���r �WW��I���@t�ig-5m��ʏ%o�!�c�IÏ~�����&�TN���Țv���]��ܟ�p�Gn&6�QVz#d�m!��!oX�'�|R=ǝ�Y�mۦY��ߩ������S�&�<'yV!L,����D��;(�����T9��;��N�f�/�cm��>�QS���PuN��\�U�`0��fc	~�a����=ǟ��x`nv�h?f��n0EkjC V#(��,Q�X���u�9cu�8>=+�f���L�j�wy���-a��w�����c��U����?}��׳.L��sf������i8�f��%6�䞬u�Zn���A�#�Y﮳�ո-��{�瘱��d^I�m���6��X�G�z?�u�'�d���?Z�s��M�V������K��29�^z�z���7��4:�Q�dM��s����!�s���B1�<jЪ#��-fu���;(�C�V�Z�['��/���EĒn��m[�r�P���h�ְ
�lC���dc�=��hHF�[�w��ȃ�ci���p�y�����6���$F�e�/�{9x:�+{H��s茞����/��H�GLs��$��]�,WҚPfلR9E���kDDƝ%��f0���>Kw�K}qo���*6�@�׹�V̚�1�>�]�.Kt3/?�zt45�
�/{�����>$z�ѷ̙��ݰ������k��W�ar���AU�֟��MЋ��}���*�fT�'_Z������Y��ķ��]��J�λ�"G�~on.O��8��v'�^5����a���I���,��b�m�{�yV2�\�T@<ˊ5�b<�c�������:Y����m�K|�1'0e��u\�&�hT�&m�އ3`�+��
(���C�1m�r�zOw����+.��2�%:�Ā�E��u>�2�NMM�����俫W]�v�X����M�)�T(4ގ0+.���-�b�rN?� ~�a��W�Ŭ���\����GA߲��N�:�_��̒�rj�)�)N\�"�9`+$��J��i���ot�s Q��a}�(4���dg���9r8-���z��-�I_	���ߎG���&�0P��_�ž%�T��b�𪫮�^�M4��E����U'��-�M����
�t�`OK8W�sÆr��1T`If�׾�����s�����ђ�w�����/%�e�(�RT�*I��(���3.�&�뮻�a_�җ��{�������|������p(�<>Ǜ_��Z���\�x��惒���b���|bS*7�kiq������{ｆ�������sQ��P''������xEV�]F���G�w�97� �����hSv��'�E�D�8?wf��w�}&+���bb.�F	�P'�`�%��l��B[�0�?�6��t��zg��</e9=��F� ����&+^m�ŗ��A�A�x����N,���R���u�h�D��b!����Çu����͉Ƴ�8N�8\`
'B>�P���j>�s�@i��_��W�c%+��b�a�:��SyG���2 c���}��9VF�Ф��V�57a�>P��I/@��b��TN�r	e8��de;�C�^��+��,��g��
��ί`F(-Q�؈���7���'Z�-�p+���n��-㌱	^�F��3fa��%����H��W�o�� %�GF�o�4�M���~b��Y�T#�Y9xva@"R����T5b���&#�W�9�{�-����^Ey"${"$�d��|]Q��	c�o9'B5���(T�f�jY�(ont�i�"�};����{r#G�ۣ�k��E��3gR�So7$�G3�[��g��	+�N�o����.����u�s�-\G�=�l�H�Z��Uz5�k�!V���4�GV�R�ș�%m%cr�$��\�[ZKb�"�Jv�T,�,G{�?�_Y�F�_Vg�z��܀�>3b�On���(e4"��ɩ���"K���E�nF[�a(~E�j����/�(�4�' ��G.��U�-���.4ז�a��ce+�b��Zɪk���v�ZH����wS3Q�j��kdۢ$�.�C�2ma�I�g�Z2�T�$����NR.d�ťb��!�4��W�R�u�:"5q��=U�jr(��h��ؙ��|�?��c�=6;;�⃕
6{ࢋR )�4�,E������w���+/3=��WC�K���26�|1�/y��[Yh���)�L�s+�MeF��똍����@صJ%�WZ`C�N�b%G ,������!�j��Q�퀽���x -_������;�.�
�u�d�J�1cu��֭[r�dL5rYvi��ڳc�L����l�X�T���cc+"���li�H�Z*����5��Ǘe9�g�Qv=�����(y{ݚS4_ǂg��"p���	y� m��k�.��w�eGF�x;��23;U(�&�v�X*���(����L�j<��f�v��)!S!(J@쭮�Y$)�L�3*{k�O1�`��k+�X��Wc�;3�Ѩ���=̋h���D���;��0�[�>���m�<����L�%�(�neb���J�#���a]_{XP��	Z�l�]��X?(M��!SBXZ�nN-����O�\�3и1|�6Z�Z�c� !�Ҭ����!�9�VLGQmq�k���~*�4�-)�27W?yy�n�����flc��I�c�YbW2L����
n�Jքۈ�gD܂��-g�5�$d�t�� ��D33�M�^T5Zͅ�b~��q7��CC�N�Q�3�?��O�y����<��ڼ����_�D|���,��ݴi����+�.�;<�7����M�LfY���oh���
v��$4�R�Q�:��n��h��Z�I�y�,�Gk=�p�h��`{p6�xs�����Ӛ��b��µ�I#�7�4�x�͔(�2�wQ;�=��x�`���OMT���o�d�f�A8���q�����*��L�ͅ@�i`y���*)}Wk��X`�Z̺}䞤g����+��� �Yo�B����-Y��G�Ӗ@���5|�"a����h��gYoϋ��-�Ψ��Pn呯$���������W�pD-֓��DO^yn���J�R��Cp����?TM~y�mV5*NQ�F��O�\�^.m�ZW�jtϳ�JŠ�IRF�@ }��QnV+�$g7K��s�!'�/Orgzڽ�\��l�5&���L�d�D=��O�F���_��ٳg���ئ��|���0�\e&Jl��H�O�_Fo�F�GQb,��4�ڻw��mˢT�ٻ��[炵U3���P\�2�pA�cjĥLNj�R�&�����/���k�/&�م@�c���n/���n���܍���5ev�`�/��"&/O߾};Oa�xM��n�=���	��L����H��n+���%PF�"Rk�o����E�����.oL�oڴ	����Nr�5hU0l�Ɣ�8��~�����Ъ~�Ůɬ��I�.֒Fz����Q!�Q����s��R��|R���x��Q1�<qǎ7nԉ��]p�KAd�i��鶎��@��G��@1:�	�"���ȨEU9���u�����/�[�0*⠽Y;5C�|��܊�d����h�H47C��f1��ka��e� �A�S��1�wL�0~��je�����al���M����piM��b??���\�������=�2�9\��b�#�8�<K��\�[�IѮj1O����#W0?����9b�+�� �o1���)z�� s��<���1�h��*�=��{F�Fb���n����b��Q�R*�z�*����l�
�C�nÆgϞ3�Y
!v�5������T3�:���\���|�I�p�Qe��j%s�L��<�6����?�bKmzᡊks�FSC*�m���k��,D! :��ľQ+=+��&c;�Ks�����ϧD��;#=�����b*���2�*N������Mr�C$�)i�Ce�0�5��"<k��rWc��\��|Ѡ�������ɬ���5���M�-
L�e+�0��rF��d"y�R7��.z�`u���e�R�i+)��]3To"U���X�'���.�Fsɻ]�:���RBv!����k���R�+Y�����Ԇ�d�Z;h����%�XMN�,2�V�?�i�ީ�Jyͺ�ã#��ύ���I�/�����p?e}"nԭ�ҙ���N��i�L?�d�ܘޘ�0�Rn,�.'�,���׭_c�pWF:5�)D�����.�~oo�ޕf
� p�'P087�8���l��?N {�+��}�'������s�taF��<���N�gUG�C�3u��ܴ�5��j���܇�͜�ڵ�W{衇�7�t�%�?y��8�\v�6j	�����5W^ye_��㗔/C��J�|�;�h�Gd8ӈfJ[�Hx����p��G���*���~�i��ܿ�P�b��K!y䑙Ⱦ�yIp�fsU�;D�#���}��<�R�=f�R��t���8j,�cޜ�`&���@�칟�������v��`xΧ|Q]��n
Ҫ���#-�MD� ,��-VUID7��\�$G��7W"��g�cnQ��i~0%������.��)^���Hś�]�Y��L"�A�vW��)�@sP��Me��chd�ΌY+Յ�a�a��d�؍s�`�XA�jI^^{�VF��_n 0w��t��y_;Bn�r�	kU_�<b$��V�kJ�,G��Ɋl_č*^�NAA.��f�eM@18�X&)��i���/xx�yS�/g$�p���C^�\��w���@�P�&���a0�G1��Hj���V6j�o��s�'M��(��$_�h���a��:Q	 +�7!.����/.L��LLM� �4L*I�ar3�S�;�L�}�8=5u����P�	by�Ԙ����	����TJi���<:��AJc{�"cZ[	Ph��~ː��WKj{�è��'���h�,�)yv"�7�H�`ع���c�wQ>�8��G�5�=�5���k��vW0w��<�`5O��*4L����B����k�\�o���S�(�Df��(�J~���ZBQ�r_��P�:���$.���y-Tݤ<M��h`=��@���gg�M;�y�F���F��_��gs$��f�S�Ռ�N�<��]��jHd~CM@�����b��.���·�5�b<���Qp�R��N��B��oEr2�?�)���Y�-����5�an��b�-��������C�+/B;&lYW5I�F3O0h�КYhFA�|4O�_�N#iw����2�����m"O�D*�S�`�f039x�sѯ�K�Y&��R �ި�n�݌�ܜэ����24%Z)�!ô{�.��Rޑb%��`̀�x��Ӌ�������z���K^z�%S�Q��c����I��_|�E}e��RUdg� ��j1�ȸ��&Q�7��5����GdQ�{��	c��P3�1)���ꪫ�ڶm�����=���b�:��-f�T\�1���s�������F6���>ƺ3����9�.�xgf6]rɧ>�)|�_�m1�XA�cv]LO4��L�Һc}K�o��v˺*.�����?����+��b}#�\�N5~̃��R+��<��S.(��	�n�yD:�k����j֞h�h�cc�ﶎ�Ew��u3lܸQ� 	+�����	�~��x/SQy}'�,�P��qM�0�~�~��h���H�A��5�c�ypp�|K,����@��J��v[�dvl'��U1���E{����+�"�CT���Ί`-�f���+ _�HkINc�^�_
�]H t�j���|��k�%4z�2#QKD�ƾ���
@ ����u9䏰����p��$��OI��p'�Z���&���w�Oq��C��R�[C�)A͠4�?K���cL����RV����y��$�2��O��}��WJev�����`����A8L��E4�X��I�I6>��}6�����ѺWc����y����	����4��	�V(���9q�[C}B���+*y��a���9��(�k�d��F�
�4�f�F�M��;������f���`�y�auU�	D]_�ψ@1#��J��)E���T���Z�Mx�w.���U3� �+�"f��o�0���bĭ��%�gY��u�\wե��fv!6�))�a^݇}���4��V"����+-lWY��[��J��ܱ*��Z��tO�5R��BV�Y���y��,�����i\s�����
�Powm�޽ӓrp�C�׋\kv���-�8��"�Yi��T(���B��2	5(�*�L����&�6��C`�<�s����]+�Pg�>�$�kx�
�X&X��G�%+�|2Ţ�#���7�ԛ6
�]!��wVZ���Ic9"0��{}aa���ޚ�:�k�\)������Wl��WN�<��O��=�=);�j7�o�8�h�B�-��b06uv�� �OT��hyL�)�&�5��@��n��Ŧ��;３�1-�&X�b��p9������;���'���l��ke�o�m���W_]���Ea�f�Z������'!�n���g�y�h׼�]�BĄ0®ML��p�������c��}�{yq%�����v��~��R6%rȡ!�̢sc��}��gfJ�-0�;vps�Y�3�Fᯨ"����8�O>�$�yb�j�,�e�������J~a�T�,���
��4&���^��`e�fX��}�����������0Ɯ�??�6k�	�^�����������YM�$pϻ�m��	g��]�sϞg��^^�T�p��?�������]`V�b����~��v�Nݍ"�;4�½g�sߍ��[�&�TK�+�9P(ˁhnX!h4TؙlI����!e�,a	�ƥ��r+�Klr%�����y+$y��&MS�qD��ڵ�켻�	����� ��D�f.��5�+�qJ]��3��,���;D��ֿ�
g���`���r��A�:�z�2&�m�,4b�7bK��3,"3K����rPH*9���m
^q��f�x�s�R���g�͑#op����>n�����nUO6��7���L����[��FdϜ�J��+���OK��-mi6�?�����u6�L����'O��@ǆ�hQ�T��L�ϴ�X`� �C�utlLz����hf��A���2!<��J�3�l��^*&a "4�Δ�h����r���u�b}���lϝ�7;�T��+����Tv���6�Ǡ���V���&0�_�
{M�qv$$jE�VN�G
��˰��9G��0�B�����k	��f6^�,lO�;G�J�v�uu��Ϛ<���r���ҢN�.!���床�w6��R}������H���Q�Z4��r����3�8U��zCH��YW����BVmZ�
\sP҅����j���������S�t��������O!�8�Q�P(5c�g���j֎cf\�taO�����sМ�aUQn�Z��牬��;���z?��ZJv}w�W�Z�%к F&��Ĕ�<�US)k`��M�I�2�]�3���_~a$p����d'[J�Q�f�&I--��n�JHd��&Q:����퀤\w�u>��n��ƀ�����[ P�#/�G�_y����3�A_n��l�����/����`��h�����+�G��xZ�K_�_���*?�z۶m������>��o��3�ӎ�zLR��9�������W���XZ|�e��9�x�_��ך�V��������SOqFk�V��w���c;r�X\���eb����i�<γ���P����2u:�|���2�g�|���~4~���U��ZWl�~����Ͼ��B���W��U,<��~�ӟ��͔��?��?��Ev�����}N�"�����}�'�F�Dlf�BW��O��O����Ȋ��篦>�3��[��.BBד_F�c��?��C��W~�Wn��ݏ<����ݻ�o��oy䑤JK�������}���sW���7fwaX�/oY4ʒݮ�$[�B�3�q\�f�=ISl�V	���ib�>�(�r����l��9�����?��X�1�-�ɋ��/[Hۘn��M.��n���9w,��d��ڲ�Z3K]bF��h_ǉ��C
Jh���I��G4�eC������������3����p*�Ҽ��8����eYcx�$!�)�J5�*G��g]��l�rc&����/"I<f��P1��D�qO|��u��8o�R
0<��c��֞8�׿�)5t��?j]
�r4^���Ĕ�����O��J3t�~�,}��mW�??i|%p�C��Ǌ{Ö��8{v̽�!"��x��f�+����%�5���>��f�"�hS)�:T�Ё������b]���,լ��=J-���_�K`�3&㉁Um �3��L=k�-f\I����_��0�ٴ�0g9�����3�'RM�}���aJ�h(�\G�9Qb��Q�:T���=�����h��9:rO��xYB����F��[{-k:�� �ρ�Y��)W��1`V��me��<f��x��VF����$���SJ���!.~���F����;�"U���`�k^-[Z4pA��o-�r�PL���hR�����<���#�p87n�8H/����(�f�0%j�Z�]��S�M��G�6�ԩ§X���#۷_��Ea��#"}��:�U>55�X���F���=��)-F-w��^�#�Cwa�dtN<`y(�2O�R���/~�?�я4���O��P9]~��[�bq5OG��,�{AZՏ�ѕD˾��̆�Y1�rE�Z�Ԏz7���?��/3��d�=f Y��p��w����6��t����h���1�^�ۿ��{��������5M��?���_��g�
�#�3/�S���2�Mx)�T��Fd�����6߯{��Z� _�}�e��j��BK����l���2��P؅�2a�lݺ��_��?��?a��
�h��",fD��w�k~�S�b>y#L�2�����=,M�v�I��lY��*�eb�Y �%m�={��~��y��&e&a�����_4���b�����x�<���ME���y�:t����o~��c�v*1V]�6ݿ��͛y�g�{ZKт y�z{�5S�t��9.�Ї>��|AU��2CC+"�R3�fx��h���g��s���� �Nj��>�Eκ$�D�#���5�=,�-Ǵ��Cfó�]����LhhD�=NZZ��CV��C׵H�Ξ�x3����	v��ղ�$6�0�ad�+#�1na��8��WI���N���6's�d�E1�R������Hp�nŌ�U��4��P�g^$6CX��ɽ�@����h�{�|�� �o{ ����LZ��@��4�2��]F7=�DW�X�gl���Z��'Rb���gY������G9��q�;xvjj����8�b}A�����:�Q_Bh��jP�Z����%�	��R�Jpio5��RE�O�;-{�&|U
�)�5��ImB /�5k��&X�Ywm繪U.Y�!6@�X`'\���Q"`r�u)kО�V+�X��v�F��\�����eBS��U6��Θ�4\��9�
 �yt������~ѿ�E��zο�CK�\%*��+.G�t�Eط.��.y�˽&w�rܽ�� ��U�7�o�z� 0]�]�f�Dv �v͚DM�j,"�,jq�!ծB>]�����d���^~�AV|[�g^P��j� �2��aktk^X�#������`sQ�MO$އ�4&эvཎ�� 	�����I�]e��pԿ�1�q�o00�	���r$1*azfR� M{I���ùkG�2�2�9��s.l���LS�lT��J���ca�$�9}�(��W\aAeށ�#����z� ���������w�av�UHB�"�Ȯ�$�Q��Dv�/d�*ɋ���q������]kG[dBX ľ� @0h�����}�}����|�9j)風����;��y���}��/��_���,Z<u�d%���ʣ<��$���w�3���~�;���H66����rc��ὸ��y�������/2�����s���A�?��ϙ�3�<3�
--eC<�
�Ȇ7��r<��3�|��Wg�S��L�X0�	w�1���n��F��aH` w�վH�o��	�;W*�
@��'���������k_C�0C��$m3���7l�^g����{������l3�A�Ǐsv�b��7�����K���$�z4�`T �W����w��<���f�i.����]3���γv�z��WY�[o��G��ꫳf���%���^����քf�b�Q�"K�x�|1+87��x�nE�b��K��Xk�{�Wjo�M�98�/���to�P~�M�|��Ω0(�íc5o����'.>z��՗:�Ե��#��ΰ�B@vu��a�q��@�����r�����pv��KF�@*�k��N>��i�)b�XT��C}�r�k�9��"�05���5Ə*ģ��=nN�o2��L���|0+r`�=�G�-��ff�=by��X
^��9S�H����.�EW� ׆u��R�`���i��	�X�ʻsrk����+�CF^=��5� Y�c_�4W2�i�T�Uj\�����f�L��}�v��~#�w�)�v�}����k%�0���ų֠�j��ø���Zc�i�z`�jP���Y�Ӥ�f�h��z�,}���B2ď��F��v�G�V3��RVg]�B^6&�]��\�3�@�ߌ��լe��F��im���dN~����q��ȯVK~&yōP�ԅ\��\�L-c_���'��A� b k-sp�!��@�f�$�����Y%��8���9"���Z5�j_���ȗ�ޑx�SIr����<�ש�.e�_�[�Е8�R����b��2��=��K�(�l7;���[�;�B��Z�6�����y�H�d���OJX6'�47�t�)>(&{���r뙑v2(��w٠�$,{|���E-�u�u(V'���M��]X�ro�h��r7�.��K.a�୧�~�^�IT�bad|�}m�!���7��������s��Dս�u�E%�"�;>��Sȸ뮻./������,�Y1�
s����1ʵ�|����f��t��Q�<̎D�q���c�P3��J��D� ���'�D��0��s���r����fA6)�.�v��[�΀-)�"ns_z�u��^P��|�\t�Ew�,%�@'��|B"K�����a�Y/�����9��E8�^�13 }Q��eB����2X�hN��<�����
")�voz�Wp󫮺ʜ3@��ۆ���/RL�Z��Q�������g��ֱg�}���q����	��Y&xtt�_��7�����Zq|���ոf��w�)0�����?���@c�o�]M����U�$��6��^����_���.Ql�dk!h�����,�S���T-F�8;%j̥z�n��ONc�]���GףT\b�����,%� �`�#K�6^�Z,����>�gM�e�i�UúQ5���������}l~�����Wr�\��k���"� }$�,�@ɏ4%B�<q������+�4�$K]����`��qg��u^׽�[ے��R�넅fs��/�%c�}AgmpG�^|�Ҹ�4�V4W�����% !�+U5��dmQ=X����D����Rr�e-85�g|"�-������ɡ������dd<u[߲e�����gY;���OF��Ť�S��|'���	��1�K���h��	�3@��V��4��*��,���QBgleU��(���	-�����S|}�Νi��V
�����h�d5��HY�c���%h��;#k�z��"q8��B���6��)C��J<�c=�K<�akP�z#2��o �D����Y3����{񴐁95O!�;3B2�=(�k
��sV���y4�Y;�
a�v�MW���x���#�S�X\������{C@��f��s�&�Jyi�.$��O��S�������`��:������\9s�9����v~��d=�Yb��⛽?�WJnA7����]�6�Rl��Nj�R��z=�n�����r#q��%���i��g�19�,P2[�]�������Dd��	XN�����q�h��pA�4K��B%j�;a�*Ԍ>�0z8|�p"\�c�P�RS���/}�8�a�dN`R'SS��sb�q��-���?��,�����g�~zUt(Bܼ�ꫬ�i��r�C=�ܙ��>���\c%�g?��#o��*��4 v�qX����-蓅Ĺڽ{�\����t[:Y��CZ������-�"('5B��(����u���8�O�,��M&��������d�^�j)G#	��°5�4d/��R��00���t?�>ク���?�`o��V��r�����\+�#�7��U;p��S���.(�ggfxT��Z�NțdX��+�@ٌ׹^_�Q7�����rF��Ia��V�Q���,����.c����k�d7�g�~r����z���J h�.��a������_���W��� 跿�-c
��|)7yѸBO��� 
]i;�pg���FSN�����d�E�-�_�g%o�Л��A~siH�6ϖo+r�L��M����������E\ ��X�m,�������$þzWj�����Ed0�gS4ӎ
 �i^6h�� ���Q���t�[a�y�M r>�Y/ �I]��wMd��]?ŬF��uhU�<ݦ��^b�{��4^GBT�eU��H��.�.<w�N��]4f�Ҫm]����E7������i�w��u�9��q��H��V�N�]��ٰa�%�z��Č�R��f~9�[L�a���g
c^}�Uܟ�gގ;�Z�G��L���P�m�-����ie�36`)Df�eW�G'��jE�1�Ky�H��\9ڮ��N��!d�yk`[�҉�L�	��/���u�螰�U�X��u��,F�z�P��3�RM�\nRz(�T�Ř㭺�Kۅ��0��Oy�ږ-�&&&������V$j,g?����{^g����.d����d*X�b(�,v�au�<\yTsE{�BF �j���PL��� b��/��zU"��_�ǽ����h��^aELs��~�,���?�-����7#���"LI)$�bƸ�G��%k�'�~�F��$G1
�%\�n�5��b"� �f2�� ��B�4Iq=��:)S�[ы��/?22��2Y!�,�?t��r8�]K^B75Wr+�5���>��3ϸ?,��g �wdf(:-̾���Sa������̭>������A��&����ђ詧�bZ����}�9W_}�UW]�r>��`{��6;��/�5נ�xz=kq�+�ݻ����@!=��F�ب�ti�$�Ɍv5P�-r�ӟ�t;�����Lr�	 E�Dci��6l��я~�����w�{�w�E����VQM��X�L�|O>RG�����Ō��??�
��R�15_��x�=܇���?���/���$>ɾ�Ǐ��Z�gn%)z�q�E���& �L���<����,$��t��Ѓ�`�Y�^�b�O�.i��������G������������׾��o�[���>����v��t�GIWQ���ڷ��[�	�����{
��'�b������������]7n`'�wߏ���=�����+�:"�B
	oׯ_ǡ�>���F|���mE6UC#A�Ldt�$s��6X5���|�MV9�S�������G7�Uf�ё�\i.�qVJ��+[(��,��-f�F�����z֍͈�G[^K:4���������<�)hA���?ZH9?**u�%~<�ͩH��l�����z�,��G���ϲM�/u�K���&#�R�u�~��uO�9O���&�V��^��9�=9�Y���j~�m[y�WC	<;=g��DC338��X)�&8_LՈK�Pfp�F�Mx�9�l@>�9a�'�a���N�͛a�&�Ŝ,1�I�>?��O7
��T�̾hUbf�h�' �c�l@MI4wS��pjrR���a�Ϥ�k��<��@�j)��mݝ��� *�>��"s���M��2DZx!��<�����T�~rǧk��]����q�G�b�5#�f'��,g��ݬ@'c�/d� rO��'-96�j�����8'FH����΃�Pԕ����_G��D��8:-�zM�Ǥ�em:B��+�cK+Z��\�N�{$¦��F��k8{|�z=��Ѵ��vȹ��K�Uϕ�,+1s�E����"~+���Y��z�-MI3yI�	JY�y/�Y�2�� �Dm߰>����Te�|edMJ���H���<фc�*	�5S^X>D+XQr�-ݤ=����F�h�ʘ���/����PbkS��u�N�"�Y3�vu	����i6ǂ!Lg>ݿ?5�:��������[o��c�7y��e�LVK���J���a����˼�Pd2q��6����;���sa� q����h�+���|�;���'�x�g?���?�ys��Q;������CV�o��f}�A
��sX�8����|R�lS�!v|S
���TC�i�5�F.ɂH(Iɰa����n��&so ��{8�
��!Y����6�i���X=���x���;)�o$H�ϼ	j �ǎ���c2��}�{� �Ȫ�=9��/h-|:�!��J��`�r֭/� ��/�Ø��n��[n��{@*�x�Ii��n=v2���g?����^]�(6D�]w�%�����믿�^��4����}���~����Nx��P��
-<Q��P���R�6�/�/��b��Ϳ{�n��&�k�3�fet���+����G0$!x=Z:��ƛ��$��,�#�l5���Q��1ɕ���y_���~_�pyS�t(y��yeF�*X=�g4��`Wt�£����S�x�ID�[�޷x('���5�s�x^�Ʊ�y�I-h�!��#x({&5����(�R�2�EG�(��2+hű�/���b&�	1V V����3#SF<����@��k�m�^jKCjA��Y�)�x�"`n������w�����R��|`�2���R��X�GfCٷEE�)��������u�B�B���6m\XH֦��&/�\�퇾(�(�D=����/���=��綒�\[V�T�t��QRiJ��bzz�Wz�db+��Y������酝�������;���N��²V+�f]�f�r�)��/ş�Jѱ���ì5x��tPo��c$��*Ҿ��|-�V��*�w3�/���P�/j�C�B^E�&1V�x~�液^,bpJ`d�,�$�3"�"	$�׳�Q����3�̶gZ��VV���a�'Kcrd��Gܢ�զ�\�S�Xx
M�omݴ�_�~RcP��ʎ��@�83���۩��lW1�t�=�=V������S�\0�Z薒���-{A�����Rc�<a씴8~��ޯ�ӘH�˳s�O,����:�/�m��'W�2��Qm���@�C�����k�C)w��")�):+��)+NM���՚e�����Bq$u��ئ���*�?��ĉ�O;�l��wk�"L�����@�ƍ*��3�<�^\LnN������z�Q*s��;vl���wܖ�����@%�	��55N�-���qa7����?:��0-�+�Y'�Ĝ43�[����)�94��>=�q��5�SNn�S�?p����Pi(30P�PN���Ul26=���yyA!�OG:�v�7���+c�������.����%�f:�
j���oG(;�Hdva1��e A���cUDj�i�(F�Իՠ3@I��7DZ�'�d�nDI#�~q��IF��8u��A�|��X�R߾팭[��+���]�7mŦg�8?��{ο`�W�
Ldtgr~DL���"W_}5~��_O2.|ݝ�1�x/.�2KPY�rx�F׹���E�]��P?y���y����n�����SX��e�#@�m:��}���{/T��Wo���+H��'���C��|�Xb]�N��(O@��<����jr�5O=���G߮�p����1:��]a��_{�u6�ڵ�8��3�i�FFFLI�*'akB���U�S���`-)8�H@70uhh���;~<q�u�.@'� ���[NcqG�w��X1���������Nn!)��<�Gv���6��8�T����s-(�PU��+�.�Cmd~���4��<��s�4D�,�r�x;m-.���]t����!&��������Mv{d�nD���r�r���OaElڴ���B;�R�����G��`���,�c����v�`څz��F���N��Z������a�:����|�P?uBØ��x�o���U)�x2�֏%���_:cǶk��� 9Ag�؁3�!�qG�[�n��y��'ƇV� 2��IUe�陙���%�<;[�֥"Zϣ��a��e� �s�R��z@4�	Z-.=���t%b?tv�t�Ν�3)e�њ�]��o޸%��N'_�%���Ncq���l�蹨UiʦH1q
�.�h`�lݺ�T*��-�J�L�e�җ��O�k��rӄ���1(�h���"����E���L�@�Eӑ�' y���ˀ�"��� Z�fʊ�:ږݬ�e7*�t������Q�j�r3�aU_D؊��CƋt4�jy0�ƙ���~L(7����ȋ�~�uþ�k�x�hf9��2Uq)�7�,e��F+QTg���<��+��-�Q&��i���OOM�x�k3��_h�ׯ^s����bilx�p�����sSi�U�`�r�S,�X��qq���W��3�eȭn��i䟕*���¿�UJV�6�����Z����r�?�q�)۬�Xv�t�FqVAf�\���*�f�9����-������Kr���J�ܠ�D��b$rq�z�j���0���Z�` �]$J=�����ˁv���͋�|�лѨ!{�W�����5%0E�r�Gy4�J05�uβ��S�.Iy�:-��Y�V�|Ş�>[Z�I�'CE�;Q��)gMv�?Z9o������;�/��"����ypG���}��Gm-�A�+�|�����K�)2��X�{Ϟ}�C��m��|.c�Łd����w�,r�9�x��BFe��?��3Ev��L3����� �zh��Ko�����S�3�n�R�G�7N�\-=�Џ~�#A0��}�=w1	~R�ʹsR�^x�e�=������L�n`S�b�U^����H���Ck!b�Ũ��R6�V�Õ<�C��F��LOM�+���|Q0жg���w��~4M)*^���2b�4d�e<��<��3��!���+��b)�Ε&:-�A����Ǐ� �`&�&�r�ِg�S#�^x�����+2,�Ծ���r��z�4��憺�Q�,�P��b�𾼚޻r�K
c$W��vח`�-~���oķ6gM�dֈk�t)�3��H1>b
 ��'��5��I�tK|:��,u������K��?�R��m�X˚�"f�y~g��0�cn��<5�|Z�%Kf�w\�_ݲnB+�{���b$�ML�ׇahI��h��3�T�)U1��Q�$щ��K� �ҏ����T޺c�i
�<��/�,SJ�-����f(4���-I�`2T�����`6�-��ɞ=�NLL�(E�,EQ@P�>XJ��'����ƍk[Ye�Yk���k׎��-8x�Ϣ���Y�~�PZ_�_��7t۶M���7/D�f�&f͚!}`!K7��W�(Wl�s��4�_%2���54}�D�٬It��(�t�h`kTص"�WP������� �&ob�C��#,��5��1p,JU@���<��엩h6oh���G����H˨n1K����t�9wH-����Z
�,z�^��*�T����{*"��K0�ÃC��|�k����O!K�_B�{���l�?�+=�q*z����B����\7(�X�K.��5>���u�F�l����Sm�@]�G�K� j������mAn9��4B����2CΤo�o��-���}@��x{׮]7�tq|�D���@��f"��_�B ?���OOL�F�i�r�ͷ �m(
�_���Ͽ�(p[���;N�OD��*��d-d
�v�Q�
1���#��rc'}���b��NO��?]|��L5�Y�RR�����;5�8J@$�{'�Ӷӧ-A��f�$�?��sY�&�n`�|8��PD"��q�^~��8�Gz��&�G��i��" Z�x��J^�	g)cgYL�4��%�-d��c��~r2�Z�f�i�E�5{�����R>�r���}��Z�_b��a8L��Ba!2Wl����]�.���BJ`tV1*�%ݱ����_��Wl�v�:�#���uZ�W�gSg
�:�;�`�y�'M%��{����.ޒu���b	�&����̷t2=��'���Ă�TǏ6+[����F:܁���3�}ؐ��)%�#Jf;�!��G,G+U���RJ jX���6,e��l+�h�����<����Eg9�5�t�����6pO��cX�jb1��BU�6UT1g�R	��bW1�����YY}�&n2<Ee�����P^��v�f��7s	��V��,ם��L]��9�A}W�Ơ@È�%��Y�/"���TSj3��I��5#Ʉ�j�RP�q�ӧ'�l����l��_:¼���j�TrE�Z�[�bkc����ss�;��~J�-'A����a-p�@��A	C�ִ*���O-(����y0Ws��q��H�)����E΅��B���|y^��R��ibVA�|]cruTJ��=m�S��ܜl��(��/�/Q�lݚ|o���o�38�eÆU,A�l��A��˅ӧg���b�G�H�K�H�_���XH��}���1o�ao�Je]֐��uTu*%�\Z,��%j̆�s�� ��z�����E�h��S8�C-�1�N�"�w�lf�Y�F6Ϙ���X@��S�{�f�2��V��T*��]���~.�Dw�7�{�Z�7�?c���/g�r�j"��;d0�,ZRs�QK�<�:Êy��oFE��@�V'�������X����x;ٟ�N7i�k=����W/�����f�V�TV��u-D-��kg/�vUl��ѫ�C�2�VN0�d���R���g��D�����E�ZƖX�@�;'���+�Lar�n�N0�k��I�㮽��믿�SA���}��u���Q��`��驩5k��r�H��x���O�t��+�T.�֑7߬T�j��۵+Er#nB���?��Qp4�3	P��&}��Ց�O�����F=����2�%c�Qr����ɲ���%�m �9�_x�Z��5��,78�U5��m�ڵ�\\.���h��;����1�͈�0z��������{�2���JX$!ܷ]��޸��?o����g>���/j�Z�V�Z�����./�]=5�O9~�&!�	���1(��uy[�����������Ͼ��KM��[
3	�c�$�5J��/��P.������{�l�9�@��/�9 �IN
���o�Q�,���"���/��L�6ױ�hl����6}o J���ǬaF�e�_�v[A�aE���b���cdDk��/d�8���Ѳ�#ұƈK&3�XA�dq���Ya�.�y�@�y�,&�tr�=c���k҄���&[��z���g<��(Ǆ�o��aF��hd��c���;��]:wm[��X�r^G�o15�'��&:�����U��3Z��ΰm�Kz�b��,l6�護~�zҮ��ª��f:Fȵ+G�l8��Il�C��h�򸄰�S�R,����"+�ue���F,�f'Zkȧe�T����_�̛f4�m5�AӐ��,(�_��)LR8�G��C)��n����#�f���:�S�\��%'N$ǘ���c^��i�x��R{>��c����z���,��{/�.�ɭe�l/n�����ŶY�+�}F4�� ������q��{�Q͊�S���=z�^�"�U�����8�%O���T]ѓ����z1�)�XaaaI��-��o��BFÄ�l����8Op�Ls��s�m\�uS�Η+8�e�/J�S˄wc�s�ƛ��Z�D~!]sE��A'�����k�[z��k�^���ף��n3��FKТ�V'_Rr���:|t��V��_��
��͟���^̨8�	o�&H]ƣD�T,W���j_��N��p@�����K)j�n}^���RU�_��ɘ��p�ts _
��9׺��S��60�����un)�)���@y�5Lʁ>���|s~Aqr3 �d������ѬKT5`�C!�?`8�y�;�����/���v֚i�3
�1V�W��9��@g�����<t���x�M7����c�#�g=���,���RVC��|�{ߓ�G4#lٺ5h�{?z���� `"�M�uy��ә6�: Pr&n�m�ż�������'��v���
��}Cեf0�V�0o�&Fb�`2��x@�p׮O<�!�����k�ߺe{H���?�����T�7=3��������T\�O� �\u�U<Ŗ�����hҏ>'c�n	)yM�e�n� ��-�B��ˁ/��t��
\`oK*���U�����Ƒ10��#�3��x�t�m��P^�s��<�Q��zd� �_�:�N�!j���᱔L��k_������^�kl���FWX�������~0XS�3�Q�Bݾ}�hdʤ��^��ojL(����ڰ���ێ$?�|��LA��.���c��+��,�ܻ�B��D#�0�8Q|�ʘ{��=��lz��ѭ� 4��?���*�(g�������(u�謳vNMM#7<���X����˴�Uje?�mK;��bC�L0/G<Ѡ���I�B)�RG�k1׊�Q�(��ʾ�m`@��r�1խF��g�Əl,���#�i&������2թəS�Y��,{�]<�Ѻ[���'̞		����^�v�)�*fIZ��%���W>[�x���<��!2�ڈ�V��ʤ�dy~gMU�"�"�]=u�4F���C�"�	L�H���J���`LС s�	L���nؔ:n۶���ٳ�<�򘀭#��<�U��n0k誨Vzd����^�R�0�>l0e�^9�Ry�L���u��t[�"n��25�ؾ�O�<��?�����J��j�+8V阺���>Uk���ǽ��:��&6�����REWkΨ��j<�3n<�T?�=^�|�9�s��O���S'��o����Q	a���n	2׉S	��^ub||)<�֭O��ͥ���evX�
���b��A��ʊQ���"������<���v�x���c1t-�v�+v5��v�� P�F?�v+�7����΋�zښf��FC��7�A�UX������\k{��c�G:�e��%��/��ycy��~�|�;�����GE��6� ��|����}�}�3��e׮_�О�ZNi�TE���+<�$�u`��.C5J�8����ZԥTBݚ��2���.i��d���W\qEt��[��Ν� �w7�x#��n��3'�B�\PB $k��3��5��$Ug5��I^���Je�ؘ�Yi��C��b�%�5��� �K��z��p���v��HXE(.��e0ڭ�G�С���eʀ	~)�V1�9b��M��9�����e��d|DŕW��_�ej�L`�?��?$U:3S�RN 2SZ ���|��|Ν/��¹�}�:sJ+DdE��q�̰�$��t�0�jD�r�/"�;w���O��O��������$�l|�?�"��w��iy۾}���%�Ț��s�C��l�]E�9aL�͈�:$���(���5�9�nd`�Y�.�и6A�L��Qw��k1���U�Z�"���ם��t>4ō��u�����@.�7W^v�^��	+��~�wY�f]�Ε�H'W�����Y�.p���E���H`�};�?I7$�k2�M���"ɽ�_,e$j_�X�Vp+(*e���Fߏ�����B���4(ʒ��%�B����˼�����HQ;㌭G��0�"@�uǣ���`�Pѭ�<+I���J��b��g�ԟ����}y��b i%�s�˽Jy=�լ�)/���Hf9�%ʷן�|�?y\1@��D@y��a�J'���)N��U֜M�<?����z�����S"�EE�^Ù�C�/#�T|=\,������+���FVg���f:��W^y� ���. �i?��?��QS?��[NA���hRdY�m�P7�3�Պ��d)#Q+d�(OON�}SM��1�hξ���#�e�����\���[ {s��EL�P�%B�(���U�l�N�mL��	m���Z�NF�[̨b�!�FgR�^!�٠N)f%y���Ӥ� Yذ�W����t&�T~+nR�dԵ ^�y٥HuC��r%��z�L�V��tb�a��S�WXl����SԁY��7�ijP,Uʦ���%�賤�$�6k�
۾����=��3�RRÝvafzNP,�f�p� h�R�A�"J�ڠ�Vk�J1q�ഺ���fH<����*R���M�T`
����ln'����ꫯf��������N꟠���$n@�}���C�z--�Z��]�z��7�<K���'���/Dcqt�;�<�l;p�:ʺw���ؤ�3���<����@�V1/��8BW��}�k_-F1H4���y��_~Yd���i���ˢ�_{�5�k�Aa�F���������i#�.1���'���Ԙȍ����4��6�
}���3�p]؛H�$��c�S�	�͈��N�/��b;\�ȏR��A�kS�.��<|���Fy�Ŋ����y�M�V��<9΢OL�z��tV��͕T�^r�%(�9��Ln�{�n�g~���o��eغ/c�6o���/퉼N��U+jY�tm�²�t�M�����M�t�,�?�A���ӣ���dD� ���	c��#����}}�!\�25�5~=(�������3Ϭ�}�T�y?�i� ��u��b�zׄ3���ӇNb�s�8 ���>���hx'JI�3Ԑ��6gf��;�!�!0Eȥǂ��T���H��
��B����m �˕�Ul�\�Hͨ�?wcs���d<��A�<��u��C�a�����U�9�J���>�_^��uګ����<��1-&S[&������tc��"�Y�=�"B�}{xx�?z�T!��)�ʅΫ�ҡX^޸aC9�:��֬]_����N��[�˕�,��bV���V�E�-�g���!o�61ĩ.�{����̱K�l��o9BH������*�T����Mǈ9�J��+���.L:�䥎r��ɾ�ǡ'4y��fU�ӳ3�Bwi�����!1�D����r@��w���ե�^z�9�.��-�ʡ��X��Ҁ�HE?��]9Fi�V���[4���*D���mh6t��Tnck���b����jT����8�E�*f��&��G�6�OK�	��u?[��h�Y�
��j��X���`YU�[�:"i�&bz��Yg��B��jAX�����0U���UyV�U�}\e�����)��K�Z_�N�1Eϋ�c���a�뚗�@�i8��B>�Ni�r�R��J�ޯ�{9,?�w����'��Z;?��z���ż�d����E�h�'�'�嚶b�$��A�ؚ5�>N/�[�t7	��[�~O~��;��p��˧�l������zȽ��dx�P�V�c�<��#ɽ�y����D�l:t(R_�)�y��;���n�q/����04Sl+�e�w��-��P#��q%OF���ȆV
Z�Qx�g�}�d��r�~��\`������]���n�Q��s�">`��~������gD	s���Ky��������v�޽��{��G���
��C��T?��={��ZVb$D6�G�"b6O�+*>�G�-�KQ�X��b������>��H�}��1�/}�K?��L&����o>��?��\�?��?��ĩS��2�۶oO�^�Ϗ��)M�^{-6.��@�ĴhNQ�Z֍��������}	Ű�u��A���	���{�pvf��%����喛_y��O}�S?�p7D�'%1|6�O��Qf���:7�������BF�㔿<h0R�+㴡0�����k��&�Ac�w�[t�{'վ��OP"��|�5>~�asN%k5;DS^|iR���8��s�p$�D��4�a�z��Ye���
{�bw�T|1�n%���� �Zj���

�Ќ�c�:��|(Wc��}�jU���Q^[�b�Z�UPh�3�AsX��U��eL�jG�8/�,)��ZQ�0�zF#^�� ���r�L���s��B��&��7-���)���0����*ظy�i�G��V4�-s�-V5%���Ƒs��tj�~��``͚,R�#��L�$��_s���K�i`��`l<Ww�����0�HьIY��Ʈ�3}���O:�X�'~@��\���
�4h�[�hK���k٩A�Ub�h�єh�~�x�)<�3b��põ�A��Ԯ��Չ%���a��y���āI2��R�:Te��|}�w�c�c����\n�#��䅢�(ɔJCǞ�Gϑdj^Po%k���x����C����Sڪ������`�[��՛:]�Eg��rt&�Ci#l��;��v���<�@wO^�4
�t�+�������Ӓ�����Ĺ8�"��GR����۲�"!ۻ-g��ݎ��^G��o�
�jDЙ@\��N4h]QZ-RGUH�`CbQ-,�u���٩��>WB8����bVo�pATlYvB�{J���ƒ�VE���gs�Q��a��auE�;�HB��p���F��{�-� �O~�_|�^�.m�!h"��u����3�Y��}�Q�ҭ<�2p[s=�殻����"�)����楄�����ͨI�����h��������?-GЧ�,<bϞݫV�6�@�Cocb�������b3��o~󩧞2�	5���'nn��D�J^z�g���@3���d׮]�8�����,5�l6��ދ/��G>b/#Ќ=��g{dd6䯇���2-�Vƀ_
�B<7d�PN�ƃ(�$$���aJj_���u��\�$���Y� �=�����a��zMS	,�������/�մ���o�ѧ�d���R��YcN�Ʉ�+N�L $tۅ^�h�����ʾ�/�## ��.~�{����8�$�ijI4���v���W���|grrjdt���|��ds����g��5�'c�.����j40�EVk$W'��h�w�[��e� ��yÜ�u3�MOaeEr��G�����YW">a���lN�-�o&�*K�v���k��N�q���2*͐���>:n10���&�H<Ѵ}a�q�<�|�u��]Y�+� �� ��+����8��2���E[\3,V6�-�f�x(�1Τ%����s�M׾�f��c��g��H?�Q� �[�/2�r�J��/%�o۾eh8uGT��܍R�uX�	�..5˭���c���+�ؾ��!�`b�q��ؚ`jHu137�uƘ����k���#34:��
a�D,S(S��1�o��M^�]g&��nc�`vN�On�h�0�K�h����ߟ{� "Q��o�S��p����C%��׷o?#I�#o--4�9g'�adx��ت����3�y��G9_���[n&#P�m�Y�s�+Y� ��T�TN���
蓰|��f;�Z�oq� ����1\V����O�ie����'���(� ~1m���[����-MNM��\055m���3A�h&��_*�à��D�z�����tp^���d>E��	1�3���Y7
��	if��V��6��HK��\(乏:z!kՕ�|�������Y������2d5�r���VU�D�CH�3�>2�;�	8kR=��S��܌qu;k9���>7���h5���9ɰ�2fn�U��:���-��!K�鯧���z'�r�g^.��zF�,���m�k��	w� ŋ�X ��	Z�-������^���[g̞��8E�27ZI��"a7�
5�Q.�E6y�����'g��q3z^�p�����xU��e�f�x�����k���Sݾ�y @���oH��{�^t�ElV#��((��c���t�
6?��Do��'��3����?����Ө������
��4�㞈4�Ӧ�0������~�N�#����;����t;�M��q��������֭���/��棋���ҁ�����y.#Ԭ�-�p�!�6����'�7��?yܗ���?��?aB�g�ыQ��+�|����#��e�]�e� �(�O��$0�I���%��)\�i%p+��/y6h%k�1$vC�#F�0O�[̛^}�뷾���{l9:��Q�����W�2kU�O>�:�]Ǽ#�m���h�ͬ2c�/2���q�UA��1�/��Ծ����K�u6\w�u;w���TU�9+\�5p�����< 'Y�V=�l�ܖ(wՔ�����5�ѐ�� r!�_z����Ɋ���2c���^z���l�T��b�eL��IO)+#�Rv/e�E4�7� �`�ZVv��jbђ,	
#*f�p�X��I0�mۦ��4k7�O��ϝa-u=��'c�Əw歃��:�M��D:�&���o���u�Q�#5'�-ܟ�%�8��s��e�T����re˱��K,�az�	��T�r���Ӵq&���&}!��\�1h=�k���$EK�<C��DL>	���'�F4����S���Jn�b�l��˺s��#�:�?YA&������}�/�f�5ڝ��(fƔVn����c�\+7�,��S˻�$�0؍Rȋ!k�	0�+���e���R&
��Z06�~gf�H�}�n�8{衇�����O?�t+�`$j��͜�0ӊh]���}I�%�K�.g<��M+ze�-�^�z�ECB2��E�`=�v�m�v�����*���c�H1#
�<��3�Оy��t2^.�%ԡ:&�Y�$c��Q�R�cU���W.�&z�ft�.�Nh�úр+�/y���H��uk1*[�F�L[��a�<��tg#�H#��樆bBt�b�^k�82�4�5Y�{��ͺ<���z���(
�z���A*���:!��,@4�ݨs�T�%WT�7z�2��n�ܼ�,�Y��_�������qS�Z�0�072:,�66���H��nz��pmJű��9�w5�R��銯������X1$�u<|Ko��������,��g��̦.ɇ��6ndx� �1�5�4����K9�R)��������������Z���(���bF"|�s�{衇:�sD��V{9oc+FD	��F��K���'5ўz晇z���^C<T#�*�m��s+܍cȩ�~�3�+1���YF�_���"��B�X����p��J�̺�;c��ؤD��_�����_�����B2j6!���/������O`S�E�A���ژ1�.G�'dP���Zo�;3i���\���ꪫ�"����-�QX��|�099��3O?�������}�Q���RrP��P����c��n�J���f��=vN�P֥�w��]�}�{����V���$�q�%����̾�Z2���˨{H�(H(�_z���9��d���OO�Z����[A�ROA�pWO�:uվ}w�q����V��b��J@K �P�n� J���=faKU 5�~J����j!��87�B��ද@���Ex|��/L�n��ž����Ե��F�7009��U�R�ż�ڛ�4���"�1t�Z�/ف9���,d��)ΐ�4��&c+���S��`cH,��}�6a�zB�����}���^��X;k�,˗)��v��+<���l����I\�(Oy�����;vlCwLM���K�
',V�d�zJ��T������?\NM�����9���������'���ҋ�"D�R�@J�_��
R���y�֭���k�6o��*����L��#���k��I��/�K�.�9F�0�!���66����I2�䅁���ۆ�І�?��eL*�t1���k��ݻ�6��� ,��7��%�)KY��v�|�^�O�T�-@�RG�PF���C�vT0�RZQ�
�X�U�?,V�ĉt`7oN�i/�|���Լ����{���-�ǐX��	�;d0(dD\n��Q�����RV)&6�S�f"�kӐ\k�5��9��d>Y'+���yzC/����D�〧U,ؗ5W��g��u�ȸ��g�ɓ��Y�	���'���9wZ��6�&�"N/K����F�=%e�F�g�8�>�Y��+�V�-6�
�bTt���\�n˪���v��J$&fs���3�ڱ�3ME�SY��NV��~	���11�G���~���g�^-��L��@�_�H�S��كL�咽to�l���XJ<�����˒e���&&�SȒ�8)���k���#��wg'���B��3>�A�HI���r��HC"����77i��~��k�7�y�뮻�P��R�m��rL�)X|XK�_=��ɱ����_�B[!�8���ƅ#іS�,lZ^Jy~�%�`̦͛�;
8������SO�	��L&���H��w޿���z�޽�Lw�������b[˸|�?ʃ�V�����ÿ�;��~-D�'�(dݸ'��<	.,tr�F�!�K.�d8���e�yN��sKxt_kxy��%��L�xz�g䂠�1WE=A�@Laʁ����jcI_L��ճA�i#ǂ��
	pƊ�|���J���k0��;�x�;���/Z��a��_@����~����}�O*#�͔Ge���XVa�ǡ5+��n������w����/z0��%<cΓo0, g�C}�7F�-�/�ſ����K/u�+��>���]C9�H5��`���̘Ҵjt�Xs�!m5jY�o��J�*x74<m����X�˄3Âf{�",%O7���yk%�*F���誙�j�&�|���lf�g�΂��#�mX_a�_^W�^�,T:��L�+F�+=�L��?�0�ndX���":l��b>��l�<H�[Ș��Ça����щU�FË��3a8q��'QT�xV�Z��뒣��GbΉ�������sjfZ����tJ�����ΛY��E�/�(@���z:���U3�wKSY��˄���E�,�,��ܵfTL`����L5��ZQ��O^�BYFC�ط��-0t��o�׭]��Mҵ��4��j�����ܷ2�}�L)�l�]�YP�qY�6͠[7��t�ء�x�Ȇ=��?��O�{�����뮻�>Ԛ2	��L�,��x��K������9��Lд�-�Vc*i�=^�S/�L��BC�򝩽0��HWi���y)g���>�d١e�����_^������	�u�sqƝ���0݌�WǕq0��Fҳ�</I1�?<�#zT�YMl�!��2�r�v��:��
P�R��L�7v�b)�4K)�땒}�����1:�}�-�3�Y��?�B^���`��F,�f��%w�!��S�(o��a�괻c��ԣ{�ĩ��d���U_Ze������CnL���/&;�ONO�����Ds�L�51o�¥|1r�����@4�W���f$*�G:�<}!o�q$�P9Z=��TZ=�=�쳖ڤ������:�V�T2*�ǐ���� ��
�ᑑz-��W��F|]���ꪫ��P��@ޅ�Ic�v^Dig�!z!�Q*�b�x�W.=E��LC��s�D��� X�oXy�Os�q�5�\~��	d�O,�/���f���|�`�Z-�GR��Ɩ�[���2W��+�L�<q�8xb������R����A+�9�'��Ka�\|��g�y&���� ׂEЌ�Vl�UQ������)��+���;�.DI�-CBnQ�#�/�-�����G.�9�}k�0�7�x��O����/|��_�j+�0��|�7]w��:��ݿs��?��^_��S�{)k�t�g�}��>���~����i�F�<>�����W���k��ƍ���	��ۄ���o���#���?�#�������|�������g�����/~��|�͌Y�O)h\�d?���Y���f��a�M��!�������f��!Wdn��4ݠ�r76�-�Ⱦ�l0��+��R��QK݊f����s�90��ѣoGc�aCu1*�ܷzG�����~9H�+A'QX��"׃/��A������S�G#W��Y�'w�����B&0��Y���X���*����eY��
>Ӱ�F�E�+4��W���3�1gH^c�lw����h�tz(M��?q7�W554��f��j/�/�x�}���N�595�nl��N�Q�,,e@J�4Ur:���u�	�S�P`�j���{sb՝}���u ������~�A�'&NF*f������W;t�ƹs��
�d5w���������ƅu�ە�k8��h�mR]
����:�Ǌ��xn5�bS{C�Rbu���>��Z��n���UZ/x�#�\P��;u��M*u#qN��\έ����r<��>�я��{�ɓ,0���O!��sj�@�s��*������8��7`�S�H�'E�K��nU0w�/^�~�!��<��N$��Z7?�A6Y�~P!i�D��A8�p[�2�h^��Q~V�UH"+&<��NƢb(�Z:��)a��yΒ�,�/G�Ŧ��W:�z�g!��R͜z-���d;5yz��#qei>E 8��N�[��nT2��V�95cL����$���^�P��t�3��J��C%h*mdQ�V���:t��єϴ&�PŨ��p� فKN���YN���9���[_ɝ�4D��i �n٦�q��XTN�%<����t晝踇����5�iM�<�i�w��]�@��\H	�4a^0�+��������C#~���b���K�R�%����,��Gy��ɓ�����Z��ס������]Я��w�Y���\�q�L�׾��!L��A�a��f �=�]r��O;,^�q��>�?B-[ܼik���2�4�jw�9�g�g�^z)�-W��[��ñ�0�>� c��n�Ys�w�o�gT(��|�#�4)q�9��4��Yp��4	�\�&������O~�\oW%s�����M���Q^��G�2�[n�妛ޅ��$�Gp�?��?Drt��o��if��/�pr��é;��?�q^��`u�|]�T�C��ß������%�ٔ^��u_qg�+��1~>g28��F����xV��'�`� -#��bt�z�,����n5膅��w���ζd���xAN��iDq�v�M7�/y/3{�O�Z�b�Z
%��?�H�c�N�O�<�"���@��B*��t�58���"kķd˳˙�\�T��:��[ʺ$�����o ��t���1zݔ�a
��5�ӋOؐ�k�;��lyķ��rn�4z��V�?�?�e�����-+Z����e46����'��(�F�E��� ��n4�F�.dc����5/�����.�S&�ܴ�dfU�`þ���b�6�]�'�A{�������������䯼/�\:�<�7ysgSY�� ��x%��m�u�r�Ey��}�/�|X83`�S}*~�r���	�iD#pN+o�c�6+����^zɔD�����ko�?��m^7&�/��	F����Bu�R��Ղ:�*��Q�4[��4Vͦ�f�g���!��v��=�f�(��\��o}�?��#b?L��S������y=�f����_Uvjn+���VW��:5Er��sg	�Ǽ����� -�*4���)7�aY4�L���R�<�MK�}�j3���`a��v�ݥ:#[Ո ȋ�e����@`l:� �ET
1��D`�H�~��׋��0�]��P@&���Gߞ���/��JO���RF�,�U�ƄL���cz&E�&��f8*Z+��+f+q����-���5�ƥb!�B�Ϋ>,���]2J�
�.������L0��F��*���F��t�0��� N"b.�T 칅�%�"�Y���5�R�(�ٻ(�w�qǇ?�a$u�q7�d�-�kl5Jt����֢�픂���'>!�X�n��"�?٬�T4����I���5B�ɬD��e\~ٕ��g�?�8ԃ�UmKf���S"�y�)\��=���r�Qj�z_ʁ�'�1���6����C���}���������av6U���}hh=�v<�������+��Y�a�Sz�E�.�|��0$<KM�� �^w�u�w�M��R�.3S�� $�!rJ��|��k���I���m���3�H��H�uA:s���S)�\nUO���� ��.��<sԒOq|��)��o��(G#��{I5�I�}�ٍ7	ل#�ɳ+�&�GsE��0��&p�jLx�t���I��)^�u��#G�2������f�y0���Xb��egð�27�+�3p�9精L�SO=�,��"�x
+k��WX
�h֗Ox�ߎ;�s�I��3{�X�6jb����sz��Ō�C��]X��`3]�״��B����)��;�V�G�V�ِ��͜D{q���3;�3�1w�����F�,]�Ta�K#�[D=i�yǦJS8�Px��?�~Y�b����匆����{��k��\�x�p5c[�?��ͬ%���>����6�'�X�f+��*j�z�H4)�֓�2��&�E9��\�{rf��W���-�h�*u;�R���/Ҍ���4Gd6U	��f2�\�.�O���۷�FfMXĪے����1�~�8׳jH9Ύ���~�S���}?�e������zG$w0;���0M)�[�1P�Z1����NU5���I	ݦ��5[)A�T�����p��5kxw7�7W�jZX�b��c�z�c�h����糘e�;�ڨ`������.�q$
���F&���J�,�w�E���}g#��Uz����pP�������cB!"ѥI�ScP��1���|}]�q$����	S�}Tn ς��(��qС������kF�5�_߸ag���z^ N�F�@�&��U��A��"�%�`�X�]���Ҁ�%�z9�}}�B�T)7�Rbn���63�͐r="�RVj��&�Y��뮠9P����=�Y�������,ȧo����"ȕ<:�dd#X��|n��/V�X�C�ߑ�V��<~<��0�M�th,�Z�U��YӴ��Q��o�#�~2+) ����)�%��\�Τ�޽�����V�m�;MD���?/�%JN���-d�ƭYkE'�=���'?��]�zͥ�^���fm�2HD����1�!��<x�F�˱`Dc�?�я���[ˑP��3��W�����:4�$��G�V�m��[?��O�����?��?U�c7?��Ur[�gq��uc�T��u0T鬘����{�~���)5tD39ͨv���e�]&��.+���3'�t`�YbC�֞m�裏1ԭ�"rbT�MbH\Dfǃ�$+��泛���ȵ�֋K�V�jjG�tw����8���kOw��4��ݘ��t�y��}��܄�1Q���Pr��.�T�N�u
���Hxglǎ�O>���I�D��Xw^_D����b��ɇ�b#�%1&WٟѬ�l���ZRcp@xӮ�sƷPrڗ�~4��O�T)�uI_|��Y�l�r�X���Z��Z�u�RMe���s2�b�+��7�f�ё7�)2��d���䋚��T�;���E�3�הdֈOpssCe�0��Yd9m���$�=r%�=u+�+������'��*��ǜ	���a�_}�UNw���B�����q��Ԡ������[q<�|g����c��U�)ݓ&���y��e�\1�R��B+P�,�j5υ��&q�.s�os��8�?qB�+��a���ڿq˦�(���3i(��V�H��"k	;S�=�'rll�IQ)�ѲCL��֑0���Z�c۲��<����eڷ�J��6�m�e&�����_��7>��O�u�]���<&�̚j�y���P���JF:*���c�����:�#�Jx.
��A�dJQ�r%���������r�3�228�'���g:��O|����01�UQ	+)c��~aD��ڤǼO=jRs��fX�rĨ�R�~�t �_����,�^y�h��5��,ma瘇��:8�jS~dX�֭�M�u"+W�?�X'K
����LW�T/C��qҋ�'�+w������dF��Rz�+�~破j${��W����z�x�5��<h��8l�Lw
	Ȯ[c���_V��$O�Tʧ�TK�4'�!�Q%��$����+�����v��;���=�o�����#���f�k���|"�o-��*�������mL�zӍ�V�Gwp��qR�W��f��L�H�dfz�^ްa2�x�Ћ��i����%OŒ��iMM�~�د.�~;��s�BЇ�r�j©V��P�qp�ٹi.@+��IX�=!ÖV�Rjc0�����7nrw�81><<���`j<:��K/�}��C��������z)T��(HD�W��X�*��Ϫ�L|鳈i����26���7�<r���5�]*����D��D��*�'�h�w�y�����F�TX`��*Bn� [�iI<�oZ�zZ�f���DH�����zC[�Ȍ�ְ�5�Iv<��hU�zFKAʅ�`$y;��r\+j�tj.��H)t�
�g�}N����F���3>�qG��T�ҵ��}�^�Hz�A��Uc�S���7�j�L;�����OJ��ȷ��
[i����`���y.��%�o�<y*,�ʩ��{�F��������sȩ6��Ӈ�=0zWP�dnA��IZ�%LQ����Խ�P�b1y� �j�����X,%]r�%�`��!�����V��};"ͨ~��D�#�&k'��F#e|���g&�������r����4!�k��������o9�V�H7�ƪ:�jhdd���7oIA���ݻ�r��
Mf��x���'�U��������fTck�V�}⛩#G0g����-,5��&�k.��#"˛6mV�Œ�y֙gف����6;��%�����T�3�^|��)�����a�>rt��M,a߾�#oI����d	yZ,//-;z�wl�X�Z_�qC�Zi���&O����b;m�d"�8�@m��_�{�pb�X�nL ���6O��l�[�8yz.:R[@:?�09��R5F+���}�V��~�:>|����b�Az��U����곁vضm�U���ի�R��gL�N���5�������)��b�:V�Ԧ&g��}"m������[Fg�K3���V�s$�6�Ńr�]sR�mRp��	���X6������f�f_<p������s)�fxtv:�b��0�׺��q�h&�d͚���_0#>ɖv�h �~f���-2��Vy�<:��`�K�YX)����W�:�i^��z���ؠ%�Z��bO�...�o1v�3|��z���/|�g������
�Ua7���S�M�h�?��?k�"���e#ؖ�uѶ��<�m�q�g$1�ݷ&i��Z@�͜���VtmWBV���ۊJ��٥qq��]=��ڬLf.U��9*k�`��k0�)/��6;�bE�c��.(zY��SȪ>}��A��n\^n�"eP��^�kT;?9������V]��j��X��.�*,�<���K/�G�z�j?��a�V/�+�s�iu�R�T���n�=`f��$�)���tK=���y�Z1�o��%�V��2����Gյ�Ԍ�s/t���`�^�F�k�Mi�	;W?��J߸G�o�z�:�#i���}݉\\���Yrb�[�W�����������A#�I,��m�Jٍ+�$�w�F��g݌R��"aUT�#���$ o����?��7�x#�y��[w��~"g�/bO�*@K�-[%
�-�_)&��}�WX�oDC�`k�=�:���
M���J'��Hb����6�9�,V�y����*n��~-��#ѝڠ��
|(�v�����~S�s�C��I/�E���D�� `W;0s�rc���ML������4���=_z�%�،�a��n��yNT3x��+�׬�c6�����h\��ŒUӉL��|L�T�����v�h��+'��;�w݁�sӯD�ѕ�*s�q֍�,�Ҝk�����~�ܝ��r��TB��ؽ��05�
3T�-q�ȪQ��&gfɓO>	�gn�#������J�<ٟ�����{&r���#vTX��6��۶%��s��߹s'6LJ���5Řw�e������Q�\1�Ο ��b$�igilObH�"��>������{�&γWU*�z�e��ä"���ᑔh`)~tT$?k1a}�p�g��+[�b9�>iݔ]��Lj�)''��1��ba�݇�H�1M;T��1S��s�n�@:�jLlg60����q�����Л�
#���#�$�ھ}�O%��g�鵽o��LTZ8�4��Ɔ�����g�0{&&op
lc�5眳k����o��o1Z$� Rk��<��Q���6MQ�G� ��>���EC��T��y:�*�,6���̺U[V[s�ꮝi�Q7+-fTj�U�1��?�����O|��+����r�T 2;g��YIU�91���s08��Q�*5BI�5�����F[Lc�l��U[�EB�?.��?s��jC���+��N@[D�W��{V�+3�@14�̈ u�����42(�O�s��̀M/v)Bmg�a����JA��g�FJ�̍T��C���<P���ϴ{�FP�
Q�a3S�z��Y�P����]�V�2����L�����s��by£��rV�[MP��ܰ*>���rC�?��e�PXmb��Ά��(UJ�����D>vhַ�a�I��ɦֺ�2gf�������Y��j�M��1ʰRC�������� eK�
�d��={�؅ڪ�]kĦ� i�����J&Q�E�̤�V�����xe�u¢C�ig��슣�4d��rtsʍ3j�8k�}i�O��u+��{����:��;�<q/�s}/�X5��y#�&s�Ŭsª��ROŏ#a�|�>��u����W�R�7��S����f;f�S��<�j�Δ�rpst�y�!<W�	�>`��֛�հ����Cy�����m	���`�:�qǩ����Ia9\n)ta���ϋ�`���\f��\t2�0�fD��b�^�l,�&��Z{o��d��3���6�	d*��ı��F�*H	�@�F��s�Y�iak�mx}6�](�Xp����$`o��5��,@�4O5,܏4���(˯��,�b�Z5�#� ԃ+1I�S����k1��c�LҾYGѹ�Lod�{NONik�B_E*��V�BC�^3�2.U��Z�a�X�h��M�qaҴ�y��P`qn~.�9�����ʕv�is��<;1�B���(Հ�ҒQ��iO-c@\��O��'��t�Z�*W��Myww��G���6E]�bM�}'��b.ؽ{w*c?qB�f\#�hg��]�L���k�Ω�d�S�.5nk�>��t/�_���x�D[��N�e1\P)�8�s�θQ�ƾ��ts�[��kul�!��R��ۮ�*¯J��l-��D����v���ޭ�u�,F�<�ʧ�ӎ�hy8ձ�BE�r�=���_��_]~��X@���Q��V��Naj�.�[����v��T)�e�1n��@�	R��l�����W����àn�4�Уmo�8F��V�tQ�:W�6mP$ژ��5�W�E FƜ+� �¬�Z֣I�"��{����Lw�3���"�šHQ"�Y�$��u�ٶ%���i$0�8���	�h����� �#�h۲a;v$GV�زeM�D��8�"E�"Y,���L{���s��%;��@�N����a�wM�0��,�%�!���^�<��hY�J�I��TC�<п�S�'�1k�Y�A�6	��ܹ�?LZ!�\��#�,����� ��ܣ��7��t���]��j�~,T_�
IK.3t�~ׁ����N,�����t�3(���6��R�>��5
^�N�,����s�Ա�� �p�'R���Dc������ȝ�K�|/���n���1~�i$���̧崖�0�&��lqB~�Eѻ�HKDb-2 �x�7H;�N!��;�V���� ��ّ#G$"ɉ)��i���0��C�h݄�S��^��>���� S?6bB�%�	O5yfd�@A���t���b�4a��7����$GG��9!��lw���$~{��z"=�5�;�Cs�rrj�JP��]�s^��	XϜ��tW3�5<�w�O�M�6�]	m:���H���U��>}����e��ڐ@(x`C�Q�Έɮ12�+����tsj��Pg��v�xO��ɯ'��m��P_�S�x�X�K0�.�R>B�p=B+x�M7�۷O�A�S��Ux��  ��IDAT��kz)m ���#��&���߶m�4� ����K�3���˙�-O��95�0�jV���i+.�h���)-%{�:Ԥ@��w��0���;�=���j$�.h���@#�ygG��B�ǉd;����� �v�?Qf�1o�Q���n'�V#�@� %1� a��)M��D^(A+�%FK!��W�6�t���h�ML95����}���Pl$�k�d?/]�DGL�k֚v��k�s��X���\&�=�DGSl�z�[�%�촑K����H.�۫�W�:u�����&Y��~/�:c"��:C���y�= !<a qv8�.�j-q\�NP� �--`��!�huJJ�����TVji~�h��?�� Z��/R� <�p.P�"m�����a8tQ��M:6vZ�C���1�	�_�9e�LLLF��b��;���,��^KpP�FKZ�-�re��$j`PEjs�!����S�j� ��0���Ln�@-�C/�XR �m�򳙷���y��]�������j��5w�b8i�"L��,���hy|;FlH6�2$J֫�Sk����Щ�D��N:��6��acF;*��hi*��CЇ�5�tJ�ꍹ%���#/^��� ġxALD|��	q��$b]㼃�X!$A�V���� �<*`�����)����%�dR`���/���0�&�T-`%2�>qLF^rZ|N#��_�Pi:���azk�aa�֡���7�L�v]�v�Z��.�_�	A�Y����2v��M>��*�0�ٯy7���f�%�,s�I���V����9--�𪐹B@��� �+\P�q�B5���*f=��=�5{{W;��^Y���/8����+zGW�.���hJ�N�C��[�'��o9�9���JS������6 M�ǡ�֕J�5�T!mI�b�֜ƝN���Dh0h�s���2K͍~�֔7�J�ۯ)ںuk����HN�Օf r2���������p�]w�>�W<7	%֊�>��c���L�K����d�ʠK���o���^S���[o�ݻ���o��k{��,Nd�@��t�P���㡨
ˇ��2'�v뭷ZQ���C=$��t�3�d,]�~�:X�"	�m�����������7�??
e��,m��׃`��F���{���ؕJ�
�}`GT5���f�ҥ.��=�^����TH�i�������	:�>���Tӻr�L8�k���	N
1A0%N5b�1�==3C�$Jo������E*��u͊K+��+�M�5� ��հ<�JMf�i��iN��YS3�\b��c��:s�!5�d�h�����|�'�x�W^�9�����p!�#m��^3�Q�wWͨ�Mg�g�4bY�����4C�m9>`�C�I�a�۲��
W}$�t����J��3�<������������O�,^�h��m34��|OO^vl���2W��'Lw�;-���r��kz��;�b�A��#��ȣk
��0ږ�_,jz�o���r\6�oب~�N߭HMBSGY�����1�rQ��vDc�!� p�Ļ��T�k1B�xZ#�p�^C�K���h�'��Tj�jG��wK;4$p�YgӦ�_�{v;{���\[Jp��L���f;�ۉ�ip5�j�S�һ�d����f���F"�Ǵ�����g�$�|����0�0�4��&�Ѻ ���w8�p-`��%��Ǉ'���Za��g"S�X �%	�K�$($N��N�-�jz)%�W�ДW���z) ��  �yZ�丆Be�w��H��Ǐ�������x&��cs���V��(���K�^4�ut����Wko�nt�����8��%��`@�n�p�-�.l8]8u$ mٲE3���%�ʄ��?�M7��O��n9}�
40��g�k����EW�l]�����E�4�5�3Ē�_'��O�����6V���L�̢U
t�4�0J_�{�9�k
�'�W�8q�� �IbNYiS*=1�)������{��!fX#߰a�t�i[�<M8�pM:�|7ܰT�{�!f�`�ƍk/^�"���
��;x'����n����#_�8��\�f���43 �C_�M(���c;��@�vŊ��=���g�I}�񁍍�9���e�����{V�4�={n����wY������b��U?�_��m��o߾k��N{�s�b�L�L����J�&zHL�{��jM��4�)D�p��P�Ϩc�E�5�aT ��:��?�L�V�B�Q�&�Ƅ��hd:�[��P=v��]�h	��!�oQ��%3�jY`�֫'8J1uP1�DF�.#��[�y���ָcw�ܩ���׿���pp�,��bN�V���F�T\��˓X��E���E���1GM]2�� 5  �[}���/⺘hMr���h�j@���y饗��կ>��cw�u�6d�\��U
�b��
6*u��mFFFq �
��c�8�rg�B�d^'������=\�c���pF��a���(d�v�VD�6�ƾ��xt�K�F�K1 D��ː���u6yr� �D!�90�Ñ�
�*\eů��c{�X!�_,�?�`��Bz��e������5��1�0ɤ���I�v�'�����㖈��$�7�.�-qp�{�c|ll��s$�u��<����ݽ~ LO�{��eˬ��ڵ��O�6��"�b�-&՚Qx����O�;�����qz!�4�-*���Š �Ϙ'�,(�Tt����uF�C�K���@X34���L�{�I�a?g��("}�6B��
�B�1L�̀'�����w�>)�$o*��}���0zj�o����b��H,b����-�L�Z��dn�B+C��v�^�
�Ǐ�� Z��J��$�9gp�?��ӇZh���EިQO�&[f�Yo�HD[�"r;�.#�CY.�����:��G�9��H��w͒�������[>��/~�#�r�\�8_1Ԩ�g��7�?�l��`��"�����g^4NÙ�����)�˴�h\B���G:	�����.�%$�a3衠mR�u��#G�N�=��=���##c��4���7�Ϻ�ahhɡCGI��0�����رC��O~��t��wk#i���Ҕ`��IzkM8��h�#�ځ��>�R��Y�z�o�A��nױT/�!��:������BCm����SJ/���0rQ�ɼ�	�V%3:z���iO�'�'���u�
pj{g�)4��ud^��[����_�^�}��~�ӟ�5E6��#��✴B�8����N�<�b�J=B7$�����#�Y;�M�՝�43z.��ZwU�-�i����Y;�P+�?i��P�.p�ogfg'��N�9cY�i��y�����@�����\��R�Cd/f�V�l�����ׯ��FV|��3p���.d��:D(���}��e��f��p����鏞zJG�,�q�x�8/�$�I�.���D3
E!�no�:G�������q�<ӿ�$���G����P�f��CHm����-]��g�	th!��LB���Ǝ��s!��j�<��s|r��uu�a{&JhA��i��#�.Ͱ������]r�>��D�V Do�����;���SEl��%���XZv�ȋ��;�x�%��X!���	�vh�m+��a���П�ϼ�%b�Hl�"���,��h�n�������uc��ӑdm<���;�I��|�9����˰�,�� ��@I@g��_ �rr��9?�8Ibc[6����q;���uuu�<z���Ic>����Vjd=�o��N� l�a���Y�В��Ld�Q�1�->�X�<��x8p�A�pFYv0��GZH�9��җ^zy�)"���W*P�6�lْ�I���<j���GKl���^��3���քu8`z��c�%}J'� �B3%)91��?��I��¾Ͻ�t^Bs�OL.z�j�����x�3��Q�4�����!EB_X�������<�ķ���-���� �IM��O��)�Z�=�8,�/�0��S���L|/:^L�9�L���]�v-���	֝��_�Z��u�M#���=8p�@���w	|P�A�u�/����cI��+�P ��Z���w�޽Dle����ʤO}���6�w�O�e���6(��hR���O�Z��wT4\�t�=�g)�'a��$�1I);U��[�{�?����kؔk����i�uJ&Up�,�p����qVjUR�0!H����c�qo�H��\.����%�'�Y	E��=
E=W�R�*���s�nq�~'ŠZ����/�0������ْUo�B��΋VǬOl�h~�X;w�$y���糟���ݻ��jT(6�i�P��:tH��h�w���ǜ\C�>*��S�'�.`�>Pw a�$*��4 q�$�]��R^#������~;"t��%̩�=ݍ�0@�V����A�
���O���O?_��g������gr���
e��P�I(&	و��k��]v��,���@̔�,�v��hi�vĻ��p!��Uk�Byc�H�:ܰ�4������7�^�}ݚkU�7��b�9�.�oM��~D����SK�SO��:�:pGK����"�ꎖ�<��h�%<����]#� ,����gY1���L�umo�mY�����;�"[���A���>f�H..��`}J���а+*\\H�+F)�z�̹Ї�[Du��R!�!Ӣ�}������mZ�u��Mr������E�ڞ�a�P� ���Ծ:c���?���#k�A�����r�D$Q;MF��"�l��t���<���+��(?�8b�l\aM0\�ٚ�J�4_�%�I;��B�|��׻I
p�a��S��xA1��E�E^�\���q�x�D8��S ��^'�5�n��Y��Lװ�y�$���J
���G2]�C��.A�>���~��"([*2�c��?�M��,m�MjZ+���ˣc��U���Ș�%3T[*��&}7nğ�G� (ѻ�PZ�mip��H-�������{�16(?F����H"�&��5Z�S�Ni�	#Ƹs��quH4q}JL�N"9��iх#��]��)yAu��l�t����Y�p�Ӯ]����;�Z֪�m��hP�ٚ=T-�Mp��B��ai'^��i�a��O&%�Ç��Qc�jQ@9�~���٬�3Вx��i0m��g���ܹc��k8�}M3�{l������%R1�G�%� ��T#1J��	*W���a(]}׈{z(\�����P^�*��좍 �������������*��*�\"ZG�
,�b�W톲.>r�H,:6�f����#�<�;�n�뭷R�Jy��M��v4�^�h�-Ȣ�?~��ظ%5v���|�hAd�M�Tj��Ń�R.��j7�-�r��B�xi�n�U����n�X�:�(���D�'OL���kB*�>��?�i�A��q� �t*o��f��x�V�X~��q뺶a�L�Vfp�jL�4�|��J�mh�\����g�n��hv��}�~��j?��q=
��vVv~��k�1��Z�U�G/  I�Q�Kە��5HmX_��|�Z�ַ����~���Ǯ\I��^36�w�����Y|v�FniMV�i��T(�Y^-W�$Ga��'-��H�ze@��́cRT�7�i���<������Q�~�N#�,T��bQH��E}.����PV�~�h�J ���D�q�T �%1T��yA��Y�t���[�LLP%���t�I�0��֖��1]�O��X��zҡP|�<W,�F��$�g�(q�T�]m�@�?�4�MD�F��
{bb��  �<�2y�
��4b
8 m��ϭ����5����R����Hy�!7�2e��r("���~��۶��艴��b��n�G�%���u2B�Kھ魾v^��_�9�+(£�b���' !���~��ƍ��I�K�P�^q��4�YH�ywN�}8��	�ف�=ƧIw@�"D����180P���Q `vN��N�v��Կ۷o�+��q����6͜���8?��)"�	�Cĥ��v#��υrx-�6�w� v��R$hL%���@�.@l��sU�{o.D(� L�KGM�c����"X=@ 3���'��J��9�[�}O���^�BY�KI�)��˾��@���[��J��N4*M ��'�=���@�[���_���@�{��VXp1��k�BJ���Y��^�4��j���S���\I�3�O�t��W�Q����G����K��� L�n	��D���Q~ȫh��!G���i�Jm&��{��U�\����"m�n/�#���$� ӧ2�9�&&*�U�O��h�\O�l@���Z�`S� к��>^i,�Zd%���^��^�Ի�X*A��AK�ujb;��Η�%:hG�O�O_���ib[3+���}���gM�ZA�¶o��r���Q�|�ن�`��E��#��Ӫ[w�D"�2e�#�F:���"={�8b����駟~�ᇿ��/.Z�{�%���5��ක���V�HK8&��n�{�<�$�Odak�R�̹�5 Z�+�q]6J<���[��7����>�n����3��^�%|\�F�D�i'Z��_:Ŀ�<g�fu���y�T�i���k�ؓ���E1��Y.�r}\R.s�d;����V5�O�G�R�����B��CfW���f!�=⏘(q��@��¦+��x��GΝ;O��C
)� �G����7�I�c1,!L�t�k��a~�C�r�	|O�P�ɴs`Al`J�X�V�OL� ��6��ڍRM\Y���3=��CwT�
a�E��\2�Xz��� ���� �3�=Y��HsB�0��ى^�՛�x")k����%���&�=��� i��+~>����8}�\-.��?K��;#�[���t��m�W������5�wa���˗]�`y�K�Ѿ��ݲh�#t�`��R���&k��|�D�q�¡���F�K+�tŵwD�	��@��h�9�`����}�����®M=���$I����c�1y� ���3"��?E"�>�>�/��B�O�^ƅF��
��G�Jr�[���N���d��"A'���.��v3y�'N�����S\5�6"F��Չ����4B�ZN]Z��b��$p����/!�i$8L������~�
�t�o�O��8�xr�g���������͛7󾄶o��)o���2N�Я[�i��t�z�ot����P;%��+X�c"�F����N�
�ɞ��Z_�F��x�o3�: ��8<t��M�4�}����W_}�{���+��ĀZ^���4�:�yP������K�+�c�3��6?'�aT�sK�R�R�> ��4KI�?|�P�)X��`��k��[&�H�s)�mzj��ꪻ���k�TN���Z\~x.7��%��|x�C}}�*󘒒�*�^�N�.�`���I��(�N�E(j5Ե׭���zcɀ9oV�����Q=ˢ�Vpy���,�vf�������+�Wz��J*��`Ǡ��a�K5���M��j�*�uk�ႂ�Cg!��{����׬"�A�I�!mݺ��{����ם>�^� �a�T�τqR�Z�	,�N�{��r�*�ǆ���'Y%5ޢi��@�q�0J�e�$������t�ʘ>�֮;v져��)��y�[���&@�c̒W4��p�g�D�����I!���`P��r��h��=��C󁁴[�7���Nū)D�����j�5s
��ԃ:4��0C-�*L��lA�v�R��f,�[��n�t��t�0d8���~�B��'���O�ٳ�\9m�����A@�D�� 
d��#��K��p�s�@�y�o�z��'DH�C$�֍�v�	�ޘ���΄Ġ>�Dq�~���Q�@@th�l#ρT�<��j�@޶[�$� Xd�`�BU9�8�h�c�?��[�f� ��6�-ͺ����	fK�
Z-�W;M;RBU�.ˍ���4jb�f�G�6J��BC� �|h<�/-մ*d,�!,(ix�Ҩ�Оy�g�>G�+�䍟�Zb9����H�;����F=w�y*:_��f{��5���N�b���q��8T�,�b��
�A"6���)��^J��٧���۶mc�ǌ7���A,�$p��A��
Ls��}�Ӈ@�F�E���ps�ă�1��`�R��8�G54�-z-'^4\>T>�qiB9o|]������'��4Z�b�<#C�He����&�㶄�"uLs�5%��5E'b��y� U���HN��=� E�ue�D��8��/�}E�=���RԜ������R� (�������֭c/�µD�%|�FQq��v���X�m	ᜧ$S��5p�ל�K���s������>�)b՗�cK��=�ޛ{�0��E�y�OM�����]�ۧ�������o߾]�~��7�^�����v�:}�4�'O���5�4i����
7n,:+/I�^h�]���6:rI�t��tѠo��;w��J�kz֚��{ｚ@@c#Օ�ޭ�9��^���U;x�&��>8��ܹSH=��Hw��9n�S���1N��SO=���{|�A�#�﬐5šf*�JB{ȷ���[�ӽ��H� ,qL4T�:Y��޽[�0��%������윛�=p��n��w���W��w�ޯ|�+g������� ������ĩ��a��o�����Xt�W8nI�cc�Ŋ �o^�f����a!�BTu�-�Rd�B�"��mp�k~4'�l�{��r�n��8uٷ���'�|ROA�J��,f����zz��Q߀ �b +���G�D�h#1��Z	�f�ZВ����?�w30B? ��'�h% �܀M�Za��gHH0c�9�/��w�w_���|y
)�����5�W֮��� ��J�L���-�	���A(,hv1G$B���1�]��ʍF�gp�G	G ��wV뎇[���ܧHYL�9��1�I��U4My2ŉk<Ʀ��F蟸:��X�%g S� �(�;-����<$���2 ��(ԢoU�0&�[�d9��:�zu���w?]����~�2K6�?�_�?֋h�3 �6?;716�k��ӆz~�4o�{��++ӎ-t@�풛7�|�z��f*f`���z�Ouf�~�G\��%�C�zOL�>��Y)�Q�N������	�;�B]�*��{�{�Rj]�E�]���{4$-{�mD 6��eN�׊ZB��D��_�EM�p`��7"���i(�DN��C
@k�x�o J�7�5(s�W�[�%\��q�!�'^k:i�5��iT&IQ�1�����s�`��ȝ�\�#Y�{���42�p�"
U����͑����	�>xO�I7�/h��Po�3��en	��Y�
�i��j�s�r�U��&t֔�jz�h$>i��'��hW��^�fY����RP�S����M4��{�+�@���ÇK��8q��]DKu�}�Q��h�qH����,=��=�]��<�X;E�c������?���S��K��o��F���x��,�w׺G�Y��{�0�ڵkt�_|�C�&1��O~g�@�����?��ϣ���p�^_pM��������w�u���ea;����g�J�����n r�橉���W�;�رc˖��3Ma&�wa��K�<��'>�;���;h�'F.]�l��ɉ1���[�fu���w���4�\ʋゲbؓǁ��N@��M��U� !T�������������W^yEcC���[���o�Ʈ];N�:�(�:	�o�y-.˴��&'FǮ�ݰi#R{��w;�w�_�.B�z�����ͼx�<'�6������u<�J 1Tr^��D��Y Q�D����S�`�P/U,$���G��;ߑ�Ш8Ps�����	�޹R�ԘZig%��%L6�2#�B/��eʮ���<����BG������a8��Ħ5�(�F�V*Ʈ��5=:(����;fL���}o=�쳏=��6ޥK�Kn��d7��ā?HK fE��'��g�>h�5��]���|��OҴ-/�tL��s�V+�a�R���=}��[��E��T�S�P�UI\n��X�;�00 ��	��.I�$?
���k(h%�?f�4B�1��EC��\�Io�Y��l��K�7̶���<�|UK-���%SL=�^1$���㝨q;p��~�V#8�⛡9F��I\���� qt�I���[�X��u׭M=�� {2��b~�lG��A�K/�@A�0���Ze�Аd=L�D͉�^P���B��O$t=5�9���
��CG��p�r�}���¹b��qa`�;|�'"�4��]��zC�SHXF�B%��6�ɠ��L�+N'02�PB�����g�	�>|�D4��DzB��Y�~�%������8ƤVׯ_��I]�+�s��AQ� ZP��L&�TX!n�t�*�L�1��+��W
�~��E~�XO %DZG�M��o��ƖƉ�_�|�[h��D�W {�k3I����/�b[��.۳g�Iz*zx�Ʀ�':�d���n�w��>�E�������BŻ���ܹ5O��t��������ϥk	`��4������?�c]L�a�������7��p�y�n��c��t�w���?�}(�3b���
ĴB�&�m6��<vHm�JK�kg�S�[�d�{�g�F'�$B���S��hr$7�)r=B7�ZvӦM|p�~:zi��_X�Ko����Ű�i�^���o����'ɫ��*P�1S2��h̸mƧf=}$�E��]�����F_��T��t��/y�I�E��$/hyY-�>ь��}S3S�Ԥ&Q�i�0������(�N��?���{���?���ݷo��Ptڑ'�x�c6��[ix�v*{\��b!�d�g�������>ť��d��K��0$��Qg���C{M�V�^L�vT�rZ�����֜а��ӔX0�b>���?��n�T�!��Do�O��&�Ҷ�*����2]��	uE�<i���y��1�K���
>�-mR�
�B��:���B�@�vJp쒤*�ᎎ�u�C�%*o�F��GM���?��c������/p��-M�5�O��V���;�r�������!�lM�:zp�/����
,��h)%��
z��}��n������2�z#�AKOxL��>T]V��$!Nŕd�3�O����	�.c`6�[�Y3Pt�z>F�VM��$�SELb��Ԉ:�&�>�V�R�QwZ������fnh����6VZ����)�3Yth�:,YM T7xb0wfB=�IKU(&�Ъ0A:3��L�4f�cIn��s9R$q��$�d�IRDJ/�:��/�=ɚ��>��q a��	}Ĉ�ia(p��KlSDs����>@�L�vH���C���$|����N/�bFw��>1>���7�t���z��Ђ�:��_r���Z�-	�'��#�<t��U/��Ci�FNI�j*Ȃ"|�#��@�r2�N�A� ���+�tyo%�;�RT��[�Д�3�
<�{&m��:�	5-19�)
�Y��dǏ��w��#qdƗR�<诐�a �wZB��v�E�g�O���I#�5���p;��kя ����+�:tH;6/}D�l�����+ž��̀F��co�8q�_���2���=_����?��O��@gDdtw߆/��|W�_D	,*;�������w�Hz�!aA!��D�5Y�����r�$|o$x	����ҳ�ޭ�8���c��¨L,-��3���[�}�v�$�����9 ��#Gt���:8��/���;n۶M�;�ٺu�%�;/?�ӆ����ճf��+c����V�7���s�j՞���F���.��Œ�cR9��i|���<}�]�˙��}׶Vn����'�olO��U���hr8P��s���Z�M�7<���ż��\��������/}�K�\�J�tƛ�x۟��`����Xۀ��dS�;o�&P�Cޭ��t�7o޼j�Jm-!!j�3�������ї�:K���ա�X���H +�Rp?���U�%f�ծӫ=��ST�Z�bn�Z���Σ2I�4ON>�L�rV,!"�V��<p�Zl�=�-
eG&I9�i�v+		�4�n�|�ll��VG�fy���į�0�V���P��,���ِ�����{ɥO�����(Eo��3>8�xt�
�$�!�Lќ,�� �^=�hX���$L�NB{7���f;[Л�8	��Rԍ�C���m�\ww��Q �d�K�qAR�{�p�L8�H��=󄑀�j�Y �^.̏F�0t�x��Di�ma�<�h�Ӭx7��� ���O�X�W3;[%��Y\�|a�@�"�"�Rs��=�ut�t�M�?��Gr���P�#�!yW)��!%�Iw�馛L8�Y޷TD�8��애(�5RZ<�!�n�T�}W�f�"8z#�_�9*�A�e�Kq�i`��8�X��La��'��h���L�v�o�e�SOs�>����� v��)0�t-�x.uO���+��lʾ�|$��H�!�����=�
�|�Uoo�t^.�UCռ!;pa�ޏE�O24�\~�q@J�J^�J�^��?=H(�����F�{ڿ����}�/��2{�B�0Jr!�,��w�;�k�.���=jNm�UH�'"C'��.����P���?�I�ߵL�y����Y`\�\�����z���]u�VB��ӂ�1$DwT"�19��u��Rv=��J:h#�@��'O<�ė����2F���o��o
��W_}UO�#��n7m���o�R��
l�#O;���o�������#r�]w��<��.d]������ug���.�@B����jH�{��}�l%�������ީ8Pu������s�i�n��VR`Z�kO�)���{z{8��]�"Z�Z���Y�R��N�-�܂^�=q��?�{>��n��{饗�lشa�ꚡe�^Mb�Wӳ4���ps�m��'��]�t�2Օtҏ���4�~��g��C�:���Ҿb�:Τ�*gH1-h!���F���������ꯤ��X��������?���w����9V�06�e�@�v�����Q���}�	��I�5ֽ�<P��TU��6:���s��F��{�8�e@4�@j		J��I�+9Ȃ�ZV<(Z�HG�n��`;8�QO�@(m�z�c>S}��*�*S�r�C-�YX��u��� �����{1
H������A�J��q����4�,0y���$[�A_i��ں:�՚��}�{��s�Y��U�^�uR;�L`�[ YI�q�a�B�ߑ��+X��Т�Aϸ0�9�!���|�J�8	jK�^�|����k�����X�7<8�A�
�#8�O����wz�qⰕ@Pj�nK��'D�@r�6�2��zh��}�)U	�^Z�F��O<�EdB�] /炦��ܫy��ظ{����g�G��G�\h?_���NR̓0�]�>a���X���_���b�XZ9�����P.,4f�,�)���뮕�:��9���}����T}b�JÑ�ƥ95;s��q���H���I�|��Z�i��/��/>w�0��~�a��;Z��H���M�'��O뿱+�Z����|S���Y��R���4�f{��l�թ������~[��Ń���l�S'O���r�*���D�[����7��/�|��Ĵ��w��/o���\`u��E<I���L�Y�HKBVsE�: H~Q��cs�3z��,����HdS�Q5��O��N�Ug�"�	F�ك����Çy4�To����(+Ʀ6m�Dy�Jh�����EK��j0��i�'��钪誙�p~Go=���b�/mt5��褵���Y2u.�P�.2r��Y��v+�Vzjծ����Y�K����?o��������ɿ��l����u�V��q'���֜P�#�J^XD�V�k��&�;.}�xA
f%�hT tB^ 6jݑ��i¥�PS:V�c#�%�='3Fgd���S��^j���ڮf`LY�R���4��q�xd�����zJ�������ҥ���g���P�%��C�d�ze����!����'R�R���[A�h5w޸K#�4�~���;��^�X,��W��a�[h��kԳ4!���1&X 8�Y�<՘�.z.u?�) ���hVu�Ν7#a|rb��MG���H��fxbf����2���z�����Bҳ�p�ȨQi�i�{�}�1s�p?�`}M��m޺�仧Ȥ{�z9�ڭG,0�N�ށ����������$����w�u�j�z����+Ѭ�b�]���隕k.|���/��f�&��]�ҙӧ�u=Z/�M┰��|ChD�L���55�[���T�z�w�5��}����Z��i#��H$���o������7�q��׬��\��[�7�練g��B��=}�3/�0��]���ܹ�pT��u׮�T�v���Eֻ�l������%cD�G� ����l��{j�mټ����q�.3L	��I�$�
n¬�c�-������U+����0y�hѩ�'=<:t���_���E=�If�˼qI��@+�D��"�*���Y��y�⧭�`n�b�!�a���l�y�\̥�҂v���5�
�Bښ�/������K�Z�iܷ�Ĭݒ�k���M���c�庩s�
Ϙ"O��.���J�8K�@��K������n@�X�Z7�̈́���Q�����+/�Wʝ�wPK�I�iZ5Rx��|�
�4!�a�$����M��(��eH���\)k�3�1����Q<�YӒ��D6�fbrα�?�W<i�#��& �v��H]'�k#�OZG�%�\+���6-4�".���B۠L̿�ۊ_@ƞ5b%2� q2b��� .����ImL�3[�g3&��n/�pm�Qo���{�Jlt����!Iے�݅j+봗�=�Q;4K핳�Cw�â���P�γ���_��8�?�n��V�	o�N�.\�wj��Δ��J�' �,�,-�fB�#�gU;����L,Sjb�tR�%@�$w(�&I���`lS���Rh�M|�TډGdjޑI/e�ee#��T/����S�ͮ%��I�$�W�7���$pɵ$��4���hU0��{ ��N!�zZ�`�X�+B_uÆ����0�"�$UyA]�/J�OLL���˺ط�R%l,H���^M2Ŀ8!�b�hY�T�����o5���C�.����7{�O"��|�D��4?"1�z�A%҇@9�F�+p��#	�b��i�i����8m<Lj�,����4 }�@�#Yb0�0��RpR j{��ɠʡ�@�w�,��Lo}��)�{J'��4� X�k݂}�M5�|�dM��U�45N�˴`(
�����-^�d�ҥ?#�G�{��{zeh�
r�qM�妗"ɏ���б &<�3�e5N�ٳ�u[݄���6����Z�FH��@�����1ݜ8M5��6�7/ �խ ��tT_V���=9̢��3Z�iQZ#�0nWj8�|�@�ú|�O�w���I/����i�y
�n�Z,ȱ���$*�&BZ�j}��ԼzBc�'{���5��|�m����%���w���7�W��BˡiԻksꯂ��^M�	��\��[k�a��_��z���˿�T�q���⋏=��Yz��(B�wh�t7=K��@*�]�\��������AJ���P�z)z�]\D=��1L&�|B�S�h�jΟ����GZ�;�����ѣ����.zJ�����f���i�R�9�����̮&��*�l�L5�m��UFBQ�t�$�\����3)��x���)�������Վ�i��SE��4D!QXOp��t�7�.X�C��4(��o��ڍ�%}����a%l3TK�w*��x ;�Rk�0Ն��:�����
����^����r�ew�K�=\խ�����qj�S/B$� 0(z-<l"F�3�zd��k�B�v�k�g��NSRn"?T���p�)�S��~��V��"�I��������[^݌���5҄0f��b4r�9�]�c؃n{��\� y1_���~��!���g����Ie��u����81�B4k׭��\*��0bz%wZ;F� k[�Ф��%�]�ٴ��Z/\�/�a;ꜛ;�+p�&iI�M���6�]fs�/�:� �������Px\�=����c�"�iS#Q��&A��H`�5�@�{O91�����3b^T_U�jù�x(Y�ģ�a2n��q�-&C)NMZ���K��d��H�gCd��'|y��څP[���u�HR�&t	!&�%�Y�X���_59��8$x��%�T���~&<�,����*p��]��G�� �Z�4L{���G�@�JOCB�ӣ��)� �~�}��U����(0ܶm�Z�غu+��d�:`����'&�P&�N������C$�q=���;����,6�%���-�W�2�3C7��#�"���~w��R��7n�t���Q>�v�H�}ts�Y�xNN�ޔ���0��G!z,磊�>1W��i`A����=��������[J4�Zz�w���>��a����"�Q�����7%��,c��L���s�:a5Lm��t�6-7([A-a�B�#<A`+0Jh���Z�/i#<�jE��m�9���,^l�v3/�B�	�..ۢ���Zq(�cV29�P�����]H�GUh�(���ri}���o�ܨ�̓��Ӑ��[��[�����?������+���7x�����!�D�A��s�\����E�%i��]P���4z����WAJ�T�j��	���ArƩ2���!�S����:�#X��8l�[ZvN�m�����韞|�G2/Iu%�5*K�W{s"��L[Y�X��j���p�!�ߩ�����Դg�Ùѹ_�w.[�2�~���E���f|By>~�4eD���ke�w�j�t�ԩ!uj,Y\��S�V��<��SO=���_P�Di��v�6?���3����ܐqA�����ǝ,ɮ*���u��fnm+Zd�\*�{{Z�V4S�n��h5��]��o�@��Y�/��G\Ũ�W��M`i��{�BLz)މ�9���-����B�90�=�8��,0��!霬D��P �A~1���(�-�<JX_���N<�1�޹���/Ű(̥W+�C;
��c�&����0�G���?�f;Ny����u�]��:�z����1�Z��@x��_�h�w�x%F��݋����X��:�o��y�j���-;���� �,��u��~���<��5���u5��k�I����Q�竔�ĕ1��[��˓�4S��S�T�J��&�KF� �0-0���tsIõk�j'IW�b�Zh�)�$�����|2U����i��GHȲ��AN?E}���J�U�p�s�$0ᨣ4o>t�`����XJ��^��ľoq�Y�g<+�}��{�!����Q{t#i@���Cw֕Rd0���B�9A�ƨ�`~�8$$�q��+T��7m�䦡�h5<a��;w�b��@H��ش�z �+ޣZ���zЫ��JQ:�n���)�	˴ם��5H��9�e�h�q�6����i��9rk��к���b-�'��}u�E6�FUN_���җ�$�;�6����趺 �
���T۷o�>��曁2(�O�:%�裏�˅/�Ϥ�)�t�����
hHz}][ZS�|��4�]�vi*tm6/�Ç�U���L_��:�J3O����ȌUt�;\���Ww��q0�Z;=����8���y�h�;G�������6�xJ|魅 �S�̅��k��x���%,�)���j��"BJԝ_�.�߱	sk�l�x����S��R9�����
��E�ա��Ju�&Mc��G��*V��c�����
����g?��'?i!�qk�aTҋ/�H�\�W�C6gɹcp�aGQ��ׇB��3z1oƀN7!4�P�PgCW��S(�ɭ�4�~0W�s
�T'�!@ P��i��%D��!�E�B�X�L1��)`i~�=9�2�9�[X}Q�eN�����t�T����,�,��4IBl$GM@��U�_����y� |���%K�I\LNv-�a����46����ѣ����o<�����t9 ��r�+K'\��	�ᩢ&��Qk�
�y�Ӝ/Ќy��gT�Í��<��1o��rd5�F ��+�(S��aM��%-^��k���+��*�/N���=���� �+��-��Nd恏I�.��[��$�#��m47s�s�)�G �L��Fa�-�W�JY����|]݇����/�E���'�Ԙk�m7��!���G,��|����J�כJ��]��x�����,���СCZ&-4 C�nR]L�0qτ�o��N.i��++���lz�V%�(;^���p��^QH�78`-��lk8��t�.X�GDu���!,]�j@F֏D�|(v�v��_�����x��
�s|�tB��3-Q�j浮�2VPB�D���;�jz���+�l-�#b�
A�#��J�s'��(���!5��uL�#h�l�R& ��q�fH7tO8Nqe�$S0��KE0W�ի��U��Sj�H����CIˡ;�ٳ��;k�`@�P�
�XZo*X�]DPթW? U�m !=�M����N�8ǯ�x;M��v�E��u�{M�yz�i��T�I�!C��cW̑I�H�(�{���]���ߎ���j�?��{=5x�sM��x ��k|�A�5� �vg�P�K���{&�������tX�������׺����������ׯ�V_Ԅhr��dO
"h�tC}~�M7�O����{i$�;w�����b��n�~i$zY-+z���w-��/����뮻t�i���jtD��Z5�G����)���tOI$�g�"��)_���+�v��JS��dM
{9�d�i���+zcM�B���]��ַ����O�����Ci0$Ժ�BH�Шt+��)k @�,����e�Ii��->�/~���o�v���5׬ɽ=�������(��!5�(?,�p������[�7Պ�M�x�4��ͪ�=2�Zl��_[�nշ�'�P�_sBNz��um0������ �$ه2��uqo@d
E;���I�R�Ͽ&���r�"��SYiE����sWCf� Z�@��,lc�ж+lu�6>]�j6���<bxLٽ1_
C['.�jv{�C pA�9�)6�2}�Ѯ��ͤ��!�=TUb9��F
%[L���o,<��؂(Itf�#�I(�R�~L����Y��;Uy��B�,4�����PF>�y�K���L���F�؝�%� t>T��-#���$��B���Sx��{�S�FMu��eP�O��;o^���<��"����Id�8r�w�՟tz]Z>O�<�C&I3���G�BYn桅�/�_�l*�7p)'s�hW�B}�3��3{�sttbuD7m�ҡV��k�d���
Ǿ�~�"��2�6��.�ۯ��Mz���t�9��-�	/��619���*���T���F	.	�PHHd`�F��2�Y��
��*'6�R0�!)y1#�
7g1�e�.@`-'�"�*���<��D�0fvF�y�5T\ҙJsE��D�8�+�J6��N�/$�P��6b�Mĺ���,��ȈN�ho�a��(q���3JAZF
��l]J'%�.F��Nw[)��'g�X0�f�DiH�P�T��i�l�8uz906���DP�˚jH�W��5	ǵ[������u[iM��`��$�!�I�q�(�g�"[V'E�b�>��	�!��I�u��ZΣ���`XeN�Vp�������?_1Y/_�����@[N�����$o��VtT$^��O��9�91,���������ɟ���t�5װ����.�h�Ȁ�6^�~�f��r�+G� 2\nP�j���B§�=
�"2��N�Μ-�r?���B�,E��.���޽[�R@[0�Ԋ���`+Ͱ6����nFkrh8A�3��?e��y��(ш�lZ���8�*x�U��d���	C?��c�S�˗-�n�'w�q�'>�	<a���N�Ն!�/2��"!����*j�a �}�?);մ�w�}���K�KE뒎蠛��B�~�mۖ��'��zD�D1�-L!o�xFi�;:@M�@G»#��{���E*�u%�"Z/P,ʕ�(�@�9�`�B�ֽ/;]+�r���:P�o�o�3CY�W���R�jA~�9�� �Rq��>��N4���ǟ�ہ{"tV�>K����� ����I�AR�� �\\��l�a�iA,��g?������h�Ӎ���r���Z����ܺK��XK�U;P���� ��9O�$8�T�H���>;G �'�7+��rH��)�gp�Q �..�'#m�,&��́]�WȌp.�
�y��(�/�$�C�i��1㏛���4~(��A,1*����9���� ���O�$_z����Q*{3�О5:h��]![�!�M��g1���%R�\�sSg�/���AF��
�sӾ뮻N:)��{��Q=���u����=���I7��g�J�n�JH�4�͉M���y��ڲ@BM�;�U�g#�ӝ�� �5���~�<m����*xz&[P��ti�����A` �/lb���Q����F����*8{$�J*�R��6#�,��X�Z@ 9��x�����W�^�g�{�(�%�t���1Bp�9�d��v4z���"S�G�^I~�m�⭚5�͛7�램s�7�j��ZW͔�h6
���鑥��ࢡ+MQ`��oQ��๾�^R���Z�/�����Z�DJ:6�mz��Υ� � �h��5%>�
��мKW
KA�,ՈQQq�F*]���n���^]jR�I`dEzݙ�WHVQ9���K���4Ĺ�$�f��%"�Q����7<<L�H�w���^xA��
'��l���# BR6�
� H���W�k���kA2*�}Kw��Ε.�p��	�
#\�[��?���_y�m	=��
tڿ�f��>��쐨�8�����ʡC��Pw��A9��DТh��D���o߾e�z}B,��$�LK�]qἕ�j��t�_|Q��2U�w�>zɒ���t���3����9��ty�-s�	�y7��~���q7l�� ��ZJ����h,Ă����}뭷�[��&���b�b��7ހ�0w�����-��+���~�J
��T	�B �9��I�jY_�V�%�2�SC�=�ʕ�ϟ���h�4Z�18�u7:�<4f�{�Iq��o�!�ޙ3�33!��c�\�ߙ��E��aD�΅ʨZ*�xe�حz��lG����Zף������|a���J�����v2��;��SRh\8�H�=�S�YvU�f�Ϭ�h	qC|ryH]OB�𙡖��n?^s��V�����<��]w�eurժ���-���26&��dq?i���x��Y�Z#xM��O�R�1>��'Z	�bd+�u�&Y�T���d6�^��Y�@��ы��tʪ�s�����!hA$f��q����~!�����!]����=礕�oG���(�b�·nZxF�gU��K��K�� (i��z���@2�\h]5��ˡ��l��9�eu�CRU66K�|4�l��\hB$����/Pp��%��%~�QuR��uaA�b�B\f<-���M�OB�w���l��9�K�8�7	w�КA�mda/#lDq
�:��JxI��t�'g�k �>K�Z6��Z��f��K �!��ΠK=5T�K1���)\�Ԋ�ɂ��HSG�xWlb[�О�)fqU���yG�(D��"�̥쐔�M�k��& ���)j���kC���j7�EP )�p�K����.sN0@�d�^�YK����׺���j����%:eX8�D2}ݺ��M�q��*D�������$��u�F*�vi��`7�~�O8��G��ͩx�'���FN�^na�b60��"��ꫯj (k�^s���޽{uܷd�mڴ�p!Q򢀒zA�-7T)ZV^>?*�a�#�6&�)JdS(�yW��;�G�~���o���a����ϯ�XX	0�m��Rڂ5e��K#��I�M]huX��z��ukמ�y����\��B� �*�1�]�A�?N�6�Bz}����J+��D���믲4E,��T�۲e�^�dJI�z�}��xE���r�u1�z��Ç�.��S*[^=�K�ȒV$E.9U�;�C_͏vu�y�J��N$ H�rLy�6E3���?/�D�����\�fϞ=�
�ۆT��_���@�N�Ɂ�1��ᩢ�A��G�ۿ�[c��Pڱ��~�ӟ~�3�CA/{�x+����!��&���������j�
ʤA��;366��P�L %�'Uu��|����Go�z��s�Ɉ���C}z9�A���4t�6�v{�[��``�*�	�8Wl�uG���Z����7����ft��0���;)��%�`��_LD1�mI0����P��k�ʸ6H��9�,��@�~�@	�'!q�eJ��h�^�u���ԧ�E���C����2D񀒘ٌ!A���s�h�K�U۝��c��._F�W�³@]��J�؋m�>
��s�R/#M�ى��8��N��@X�tpnN�Cqzz��ޮ�dl|�E'c�IF�x�	���3l|�i�i_&�������s"�!���G���K�J��ō݄֠�ˬ���bh�J���/������,����B[�,�xJ��N۹�Z^�I��]]ƶ��I�o#m�hn6vX�\�|��a�I	$���x�-�GVB�M�a�Ĵ�ٷo�VWzTze����8=U4���W�~DV,�UP!�i�ξA���e�"<�l;���_}�)8Ð�����=ȱڡ���"@LIg��C��^O����3��X�ü��x�w������9�_�Z"_�0r��ubax��y�i�[�����{ ޤ�0��񩡥˩p�mG.��V�ڭ��������w{6t�t���^X��"^�= ̭���7�w�t&��)���e�/�]�`�D�:��j� ����,�?����䬤ˢ���j*d�������"�n���ik��R@3O'Э[�Jq�Y�|L��KA�"�m�XX�@_�Nb#���[�6��]A
]�}x���Gz�}�Ot#Y�`^:K�,U��2�]�O��כ�ט\H.T�k��E2�����VF�[Ӳ���}�s7�x�F"��Q���,�ZMj�롡BA#'+Qs�Ӂ#M�%�_H�����~>���������C	����\�{�ݷ�>�>Ywky�̀fF�׌	���dh�8vLDk��j��xǉ>S0%T��s5�x�0����� ����M�w����;�E��ϚS��=���w��N���B�S���L]%��buH����䦘m�<i��D}]�����(lM��/��S���R}���~�a!�W��#�Я�B���P/E�P�R]$߃(������7o���{���$މ�X�o�<y���Ի��6�i�J0�d�\�x�-�2mӰa�^:V$R{����NZ\9�����P P�A��G9�"̼.��o����wQ�\y��A݄�\�y�U$��.KK��ѫ?YϤ$m֛�r5){�%��:e��ZF��K��!M�L�)�g���VO�k���ed�t�.k���m�4�h��v�ʊ�����N��D��e�&o��b�q̕���2Li�[�B���F����:�5�21��&g�5���������7��*b�C����V��m�=��zCws��n��)7���\���bf�������s�+:�@���'T̉���B�#�>����	'f�����s�t
����׵/�{z{���/z�w�����ki��ٱb������tҴ*UՁ.�n�@y\tC	��S��MNN�n�8�^r`p'4Ώg(u�i%pdUJF���p{4��%���[L;�[���XM�~gɮ�u5�	 ��3f��Z&z��`��1:��==vPk�Fδ������ݻ��'�G�6��,�Iw�J��~������M�UzHC7e�i�jn|6��٢�.�L#�6
�I"d���J*
 >gt��M$N�xz�LL����PtV(8�^(�L�,�F~������i����	c��e���	��@mʣa���/N=��9�O�<��q~�|.t�"���7Kx�U%����Eu�o��6ݺ?�V$�_���z��W�isϔ�x���tFE:Nr�t59��͛7�R�BEX��-�Z��	�⍟��ȻԼ��F=4zM�+�*ȱ�5
:i��ꋚX�YXSs.���K/��;�S��z�eث���>}�za�5��`0����H�EX����"3�$�S���'�^#���t�P��:;3�dp�G%%�K����'q�3�
k?�S󃤆�F�Ҝh~���/ �x�l�,�,�B��,���>�+(�H�,�`/���^d���~hmq��fj�t)��.AbN�k<Իk�4W��	�h!�x��p����L�~��ZY�e�F8^3lg��%/���x�^D��O�Ј���O�_��.j`��c��
iaZM���T�Ӕ)v�����6�X�$��#I�ǭ�����.V�����+&�#��=��O�b��e(���M4Q o���hf4z)�)19�ˊ�ZmH����Y��C�B@�"t��u���Br4��h�zQ5o,��N��'�|R{r.4�$�+�TX�u��R<��e!�v��;��������;�}��
�YR�Q1(Z k7���f^�I�h�P&.}`TG�8~��ۣ	���W��1�)��u���KBl��K)w�O�V�Z����]r��~��̐��!S��G���B*��p�\�����&1]*�iVb���9#�$�ǌ��z�� ���pY�t!���)H'=�n�{�St�j���`0��$!���?��������%��$����Mt���ĵ	I��r�e��>>3TSp}=���(����-?r��%��.b��w�w%�w?�h|����4P�i��+�y��$~���U|f�86L+g�Q��W$AF�u�={�H�_�2|�ji*(u�%,��=s�,Y�z
�s��㻪R8g��]5@�Op�k�5��?��AJ�D�NHv��R����	���#h��hCH"�\U�*jx�����H�#lD�
�$œЃ0J�H��P�U\�%C�U�Z⑑f���¥X]�2XP195~i����Kԣ�a�r$��	�"�C�,�f"�q�LLП��#��;U����Y��Hb�Ż��%��,���Z�.tv"Ͻ��܇���,���h ��u�j�>6n lǎMO\��2�5H�$��I���F�8��][K�/~�����?d�i��1d�g�.��lY�P	�K���hbY�ZR�.�J@�z��/5��P;2r�XZp⺓��|/M��u��!JC L�Np�irt��㬢bC_��dƻ7
c}�ߴ)O� L��+��
�
�\���+Ć_MOѤ�-�@/8�*�z5	�[o������C]A(G�7��:��ִeMcOD/Z�qmA7�J5]�蝀l� �h�\A�!#��,�'q��YV��\p9��p����ft��wN�E�4��Η��I��m�������_�e�޽�CQ�Qg{��v��{�޽��lL2�� 6$:�$&�A�$��B"M��.0n��[�[m-i ��7�k��t"�J@|xxv%����a>�ǣ@	A4�N$^piI<s{u�uב���Y��_����r	�m�d;�a�IfbA��v�X�Cc-k�V
�d�Ԣvf���%}��aV���T2G}@�o,v��+����Ȕ��Uw��nGכׇ���@�	F�����ģui���ɒ<F�
i)	գ��U�	_/�`��!��-9�{��7�����ZJ�\��P.9�*����W�v�RiugVB�b�`6���;���C�R���kgV*V�o�s�]�IL���Xt��$%��ǘ (/~!4��]\�"�[�k5Y�u�l'�f���e;�K��V�%gڻ��bPA����N9�I0=�E��h����#���e21��k]�z��f�<�t[�p��ʑ�I���UX�/H2#*����fB��s��56o)�ټ�>��>:�X�؛F�L�io��h�u ]�T�s9N ����t,X�e-�$5�u8�u��Q6��
NrHm��	���9��5�jo�FB���t1����{�2�� 1Z�3�K�nh���6oެ�:u�~��]��j$�%�&�t7i0lԸ|%�c@��6�z�}������(T�1lw0+!B|���S#%�s(ݠ�P�=_�魫H�� u�X��u�WH3��/K�b� ?	j�L��%gcN�; ��H��i2�R��T����mz���h ����%����`�^F�	�$��ۢ$H�0P㑆���\+H�̂V�7xqR���)z�*�Da�3��p�am� 0�6�(��4W��>u��4t�O���i ��k1Lw��z�-�|�k_ӭ��]VU�o{'�sH��I�%�l�����C�ѣ=&?�k�.&p������~���8�l4��n��6�U�
�7<��F�ɭ��ٳ-od���ז޴i�����˓
:r��֭CK-_n^-$��UBU<at_%9=�D.͏v��=�}��"�krX��Ij,JHG����}��SWA�����E����8mKzDR���aȳ�ɀ6���$ŐP��a��_ܫ��>��[�O����y1m�)B	4���Kz\FS��qg�ōf�������Mn�����̣Y�H��a�깱Ȇ3�����	�"	5�A%\�Z�9����v>ԕk��>�����9rT�?&�`ic��6h��d�E=���U��.w�V]�e��@К��k0A. �&����4�$P[�+%LAr7�l������x��v�Np��r��,o�ֱ*�T^^/v1 [���>����C�{UJ�do�=*��8��B�zQR��W�+|�L;�B�}p{��^o�(8b�)w��p33� ���I	�|�3f���i{��6���:��5��2j��0v]I��*�������y�l%�M���D$��O�s�Ĺ�V����E��,��U�bM��$�B3����}�B��f1��?E`�_�J+��i�sIB�v �JC:Z�|3(ǎ����5�7;�ŧ�zze�V\��n��5�&�+m�W^yE��x��g��kא ���O��a�<�Fć�$M��V%�V��������.'���z� ���w�w�~{�Rk�<Ȳ���gG�M&E���"�TAQ'��7��{>p�uU�⒄{�.1�qL�Ǳcy���lɒe�CK=w������۝ Mp���������ֳ���7u��<C��amt?O>BH�0�ޑ��߂�E�����8<�s""�ym+T��ʇw����X�' 3�MO_ooŉ�VZ�tV�I&
S���VK�b[����I�$��X�\�p�����K�_�E� |�x⅛t2�q��	K���{��	}�s�D����+��]�q��4��+M����j���"�!-���
n-���P�uƃ�4.:�հ[�ܢ�E��4L�v�+�F�0!6�kh�
=h���d�1�B�]���u�)�� ��V"�	L�
��l(�v�H	Dn-_>N������#�biOa�����}����m��g�8��c{������G�J^rX�A�_q��U5�	S}5 �FS�cӻ�"M��N�<v�ؖ-[ீ�� O��`�X�����"��n��v��8@0]#{�ۯ]����6h�ǀ���7o�L|V��Y�PS5|�q߫�ԩ��肵kעЁ틆�w��U��z&��t��k�5�z��o��F
�\�v��2Ь^��oa8���5㓓sH�饄�9���ٽg��G���ZwW7���Z\�F�k�"uJE@��c���s5���E	��Q}�� ���9l(�@!�
����P&)�����S�k||���_��$v��N�DE
.p�-><5 I����U���� .�v�%�^�b!l����ip}s�94͈�y������)�Lgܡh�/�.̈́��a�2�*%��������1\V�L�\c�G\;��Cի��]D���Vum�Q��|�ei��$��`��#�� �^���N%�F�zg��⴫Xd���V�Ao�;*�B!��C���,���լ��]8?%�t
q&<��1GyYM��~M���	�L*A��Ys���X�u��B��u��L���*��_4g�H�ajbk��Y���;�+�c7�\�K2.�!9�2�8� i�=�^$���S�격 S��GS1V�	��I�v�+�L�CRɦ�O8F���0j�)ϲ�ͨۃ� #�X:h����Dq&i�$[�=g?����Ӂ�p]۵-�-���b�����H�"��%Z���e:��_�B���HJ�:Xd*	�X�c/�In<4(�d@���3���:q�9�\@(��\��v��p��c[*qf�ZY,�d\���`g�ڎ��ţ�T�&(�	�|�+.3�/��n.���}��u�|�=���m������U��h��l�@���t4�aS3CK&��;�Vj�Ww���ۑ��j�ز	���*izr����7ɽ%>W��3��CG�+�e�]����
�(�A#E,G+M��^J0Z�kt�lj�^G'>K��Ϝ�m|=v��ч��k^d,m**��/� ���܆���;D�t�U��N��^���A8@��z�Z��v�M�0��C�S�:�3^����Z�{j-R�[�t�j�hC��n�q���:���  A���-u�3)������W�Zq����)\�M�Jl_��6�r5IԙTo�'��01M}��ЭdUR�V�̧�z
��E�룏>*����
�脆r ,����[��N�b`��ڻ�Ν�iǎ�N�>��K/��B-z���,E�������.5I�ӽ���}������ݫ������nh���Kڣ���.��uib��r�a"����t����5�_|�E]FJ�ވ�_�W?���n��h��^;>1a�r�dZz����Jo���^��/�t��g�j��?P�/�!W���[^$ 5�GSNU�@#�[�'�
����Ш�C�m��?��t{Ml �2�l��j!��=~�}}H_�Պ^�Pm������1ۈ�8\%@v�T���:9JuG�m�n�lh�z��D��u{���ːrI�*2�6��C�tH��ގ�i���8V8�p�T,;�9�ʴ~�P����~ރ��+��5�U�Q��j��>�`���)j��B���x��7��@��drq�1�J!0^�`���2ӫlu���H�D`!k5z<��� ��l	~@� A�㝴���2~����'�j ���pR$wHŢt��P�]e����z0��� !A��3���F����tNGT��Ya�ݑs�}s29��ds�����0o�(��0�9Lk�� �(������/ ����3�c�b�G�Eo�Nq
^dMK]4�utt�bL�W�B��_�(�Q(�A�|16��4�����ݰ``B�Uk8� WJ7'�4A�0N���IE^$�(u�Yx�����~�+*�����>��^vZ��$y
�����wB{����eiO��D ���S�w�՟a�8$��J�����*���)%�����b�TYXyv��T'�.��I�W�}��u���cAp�҅�Df��5pڲ�^?��O�f:��zwTٴ��<e�eH�.&K;.�� c �h��.��Մ�B
���<Pc�ʘ�5����G���r5�3�����;���Y��w��K�|���&�իȲ��\c�ARD��s3����\&��eK����v�"gx^���+��z������Ò�4Dĕ�@�`q"�FP���Gw
[4�W�Za��7��G�v�PM6�țo�iۨ�h��\��ܹ�*b.�i�:'����]���_��jJ ^s��"���s�=�쳚��Y~�~K�_����O�B�le�����)&���O~n�~R�u]����D(*	R�/|���|E�z�ş���뫯���S���=�s�^C�������4ev S��_���_��OV�����뿂tO>�$į�'�Ջo�y3'�n��o��?�<?�)���ݻ���/�[��$�f����Qxے����)���7:��z�G���cc��[l݄<h�7�N����C� �D�����I���Y'�6S����z������o�M������s�)����D���������%�g�W�N��%˒�S��/ͨM�6!1�[외rªU+W�����	&A���Dd��3,�r�,�����B-p[1gޚZ��8Z�i��v��xxeV.�,<a�%54;�s���창D�*��B[�,.{\:�Vl3J�K�*H�̭��Q�*�qVDgC��	��YQ��{������ o7�N ��ɧ噊�oPb��J=�Y���(���SI���
�~~a�8���̈́/��}�Y�ʊ��66ȁ����
!���v��|�^���o���q�������.��;�e��������*-G�
&��1Oұ�I���,��$�?@�����jbc�@o�k�a��D����/ ���*\"��'M^�gKQвPo�r/�17)��Z[�F���3��)�MNM�Bt��!5R�XPӈ�h��ӞUk6�ӎ@U�D�t�Ri-�Hx:nR F�le5O{A�6 �RfJ�D�Q3y%jd���D��]��A��o��(�Z��M�XPB��Z������d�'�{v҄ܠ��ҥKM׉�IF��Z����g-�>5IMWB�A�K���u���)�d�"�v�Θ1�*U�F���< \�)]C�
���9��.8�+Շ�F]���J�p�ڞdN���E�5j���q��TA-�񅙭�[�z-*-�.�aR��y�6; �)�pz|<�O�冗��;�C��
:zrxU�h�N{B51#]���۷��7����{=zT�YB�UOꈟQ{[���"��a����x.WO����L9N5��]/H�k�8j���P����h��+���e��3s�y�(�ǃ>��u˖�%!!lT�ts��Ћ'�4�TmOJ"�X���*��-���oئzG��; ��\G��G?���/��;
��/���������g�7�AB�C�U�4px���_��_��O<�D����:W������^�<�2T;�{���}�{dE�R]N����zJ��˿�߮^��,�2����0���?/p�b|��9zQ5�Y'���_m0�Mieq�9s��8&9\ab�1H-B9M��R�.ӛj�d2k�lJ��742-�'�A�W3��򬬹c�re�˚�1\���>!Y��ZJ���V������=8ث����0	-�5�Cl�u�+��uC�L�S�IPő��t7}��c�����C��C5(�Ӡ�=�#t�=��k�.����~��&8v��e }�_�?�S��b왩��$Q�t�uj�d�����ިu�fȞ�Z0����>N6�z˶Ā� �wP�m
�ĩ� �%N��d��/�S��Z�.h$F�ow\DW53̑�h������Th5�E�� �y�Y��ꕫ�5��J:�Z�'J��u�OO� M��,[�	���J[����<�n;G�8��+n�,�X+�+���?].�6*��ؖ��F��[��t�&E�KŹ�S���	���>�%0�&�ԛ��F@�����K��h��q֒M�|������u�&#� $����NI~�Άd�]#�`E 59��<��b��{.Z�Ң������,J���օk�is��A����N�M.�jÅ�0�oEꗊ�Xi�248��?��W���#�	�Ȁy�yS4�3Nc��,���0���,F?�7�M.T.è��Io8�o���-�Ҽ����Ź�9��0Rv�VY\���]��r��h7Z���[\(-V���+�gg��H��KE�y��f�5��3�t��P��d��{�p�n�Lӝ�4�_$����r Sf�~4N B�"���g����>s���YS/��1<�F;�ׯN���~��Y�tm�D_�l@4�*t�W.]m4Lj|l�9o榁Gv�<����5|)�9Xcc+|;�w��+�b���ԩSgt�H*᭔�`B!�o;j^��lO׮��2 ^���&���Cu׈G;��,]0�:л0;5;e��1u�\�0�?�ja���Z�Z�Q^�z������ec#W�4�\5�RA����K�/`JN���	�z�JK������FRp�L7W��wީե>�?ե:<�'?ٌ�A) e��ӫq&a0�7t�:-�N߷�~�3U���I!�j��s:�G�}��r�u����+W��ӟ><�n�H��x���ɑ�!�!�y�\8`���G����)�VE��()��A�z_ �|�� S
�Re|'�*-wd~��W�<H�\����|�"�rإ?��دN Dۨ��ݽp�b���5Y}����[���imD��x�^G�����~��?�f�N:�����g�;{���binAGv_���M��R*�M,�Y�O|%02�5���ꕬ�sȉ����~���;w���?i5éɹֆHC��y�ͷ����/)��ѣGff�o�e����oہ�j��D6(�u;�����>�V��5�tk"A�|(Z ���m�V��j�je���F�99=����.�ڕZ�e"Yu�ͨ}��%$mɧ�N�G@o��1=9U��z���������t���e���K��b__o���p��rA�ic�f�V��k��\���˝w߮U��J�	��J��Ů�J�b/���i�N[����E�2���1}���k}��,Wj��^A0!Q�-����M��Gъ�����ٙi?�R]�]�Vuh�T]�j��Ҏ�z��% ���2Ҵ���䛁1���\��6j�t&W��s���.Wlδ<�� �9�xG�q۩�Z��-�H�[�V7Ч����
�|6��^k� �\�p	x�f�Vٌ����
�L�!l�5뭧����U����<��ݕ��J޺u��M���w/e��J��G�3��'p?
Ѡ�]q�Φ�t�ZiyY��O�D������Y�"  
�RAGw ��O8%a��\�Ӫ�Clq�����7B�׆쥕Fh�حd>�CPs�.�1p*���ȹ?m�EU�����J�mH�6j�fy����Z*iC��޸�W'R�$W��a�Q������z����3�t�MJ驧����M��Y�N4��߳��@�~�7��7ۼ-�%�'i�e��锧��{��kק= d�A��[
W*ZA�����U��2���C�Q�������G�4�����(�{�u�]����@XޖH�q�DO�yY�F��9�
 NM��f-!Fd�2֌�.�J;�*\����hY��c�J?��!3WD��GA7�t������\,�K&�8>0m��$5����ϙ�Y4y�+W&w����oB𮯃���Pu���Fg&�Ї�8nۜK�X�B���ws��)�9/�}��2�N�E����n�6Yof�dSI�@])�27� sK���'������j��I��L+<�StES����e��~�Uv��e\��2�$�!��an��h��W^yœ���n�x�^Rv?~S�HT:5��/�	8�A^�ӂj&ymؠ�A��Ҵ9w��~_���43w������`vGcXd;��!5�PA��2�U�S
^sI��i�&����D�(�4$��.�r����V�����t�M"/��r�'*���0N��#pl��G?����`M�2W��&����3g>�bY%nN��3"�V�\��D���C��q�>A�?OH�\���!x���1��s����bawy�����j����Vй'��a���[�7<�hX/�����ԇ� u2Tj��w�}��B�1�v�Xk�!ۆ��ɢSK J�ܹ�[-�z9y����E0Y�ҝ��ѣ�H�sSjN�g�u��f�X���Eí�c9�~=�6���K�<r��B.�A�K�]QE����=]@|� @-��E��{WW�ؖ{M�0 tP���R0=�� M3D
��G�Q;�&F����zeC�XbIZ]?�	���rlq�g�7	����2�6p�	����9"k\����YS8���= �J�uw*��Qss��Y�F�D�) թ׹�M�8� !*�+���U�)Hjuh���P	dh�Sʥ�-��R�_-�&X�o5��S�����؎@b����[e���gXh���cL�B\w''7�pغ�������S�jQ�㢙��ΝG� )�$�<�4=�<[LH b;��˨]y~~!��X��\�����^k��;��p�!T���w��<SՊ��BSDnuw�h�"��(�Bsm'�s������m�[��Tg1��@�����6q#�����u��}6�SqaZsr��jG��;Æ�.&p۶mD40��������I���O�������C�>��X���p����i�si&��ĳ���M �f�3�����َ��*���K��i	��'�2�k���XfI],<��ԴE�<�^"7�rU��R���D)��q�a֔���O������x��Ol�'����6w��P����n�A7Y�f�>$���w�=��t��'��mxA�7�xC[�pZ!.�7[�4]�lf���nQ�Q_(-�di�|����&���DE'�Fd�>�v������{�!0��y��3@F�ZIv1)�}`�Cp֙
Ƀ��A�&hUB��-�J�(���4(��N =�A�����0*ʠ�\�01q]o�H�ƞR��F��UJo��c1�`�&���}O�'�7oF�1ux�vu�p\��*qyi<	4�pѺ��f_dTtȀ�X���y5'��M?O5��]hj�Q+�e�Y���,,+�y-�F��9��������N�N B�P\�U'����!��8�9�4R��z�k��d;�M��,�㈟�"�.ض\wf"�M��b�\��E�6U�5I/8|�0�gl}h"F��`^�V���R�@�@�F�7�	��x��BE��I�@�[7a�
==�vc�9ռ�֋�nͮT��\Us��\&��]42��W��B@��ʆ��I�c'��N~���F����p����"A
V.RD+WCb+k��Fh�ph���b�Sss-υ2�V����i�i�X�5\B��a�*e�4	,s�'	�Z�A\���=����ŦD%���?��U[8"��N6��.�ؚ�d.�I`��6�u�ʜ&?��<00e�^�<�Q�x��/Q��b��q=o���%x��J²ǩx>5;d5�RxA��^�B�+� �ӱ K#���6���[��+��a�|��U*U2!���x����_Ɂ��B��]CH�']�o�XQ,�����N�
���*�{R��f��K��@�@:=g�/gsD��H8K��;;�3��|�C��+�����CDP�aք���	�p+.���������m!S=���λ�,�ҺX��0�d�-u_ǧU�mCb�%zt�X�����,�� @��a,y�����a��h�C����97?���w�x�G�p!A�Ȳ�ҩ=�f�I%.��F#w�u.�ďb%��B�ZX�*h�����|���]^��!B�S��0���gH�Ay �CoQ)[�U�ȱ�~o��j���a�����V�Yc|j��@�����Ar8���y����҈ד ZA��x�+΂�͆>.K�����b>�z��?j.s�쪛�:�׭[�v�(��>��dMrZ�!�� v)zMnv�Z��{��φ��)&����E���\��N������;��$�o6[��S�����JM{�"�fVlٲ��FE1�%�������gy�J}�]Ds@�mwsbVڊv>�zR������s�sڑo����ϝs/F����Z�Qۖ<Y��/_�����ʐ������4����˦4�Mkns���W4=�p����^b5Q���E�tsd�E8�:���0?��>���x��t-CXw��G���ƛ�ZC����"����ٟ��7���ᴨ���}�К���?�q[`��m{�6��ˊ
�p[50�0�+�>��'���mG5�βK�6�A@�ktxDw@H-�'��
�́�ߵ�R�L��<���!�Cy�3l�՚&�RA4!V�{��܆��`��i���D9A9I�Zm�
�$sO�2�3a��I��|�̃p����0�0��8�u\/㋀��W�0v�_�Mujb�'� v�%��ԏ�4��C<C�_L����k&~>,r:>���TC��!�
I��ڮH`	j�&0�Hf�Cl~��b&���dbَJ\ל0Y��xO��v�k�$�6�f\{�t���l����h�Je�TСꇸ�	L�5��;���Hm&�&��ê$�ܤKq!c h����j4��AԆ��S���t������TD��e&A=�N��#�@�}-5��eѢ%���(ӊ3�i���+,�߹�ف������,��BN^6
T%�J�i�:� �3A����hO���M^n��}R =۠'�'}��đ��e"^�f�Uw1������Y�##��3Q�Q7Y�_ [j��Ic�[����קO�������s�L�k�Z:c�Q��e�q�,Nn|�ԁ��!��	��Jz��𞧙�@�V��:�u�7�|S}�-���.5 dCq�\�kW�v�Q�ר1�5To���:���EW�^	Kp�jU���ؘ�s�i=��,�h�*�?j'�`}��7�:�_�	���ɔK��ƍ�$�DAP��]p�,�* �z�ȑ#: 5��'��z#}���^/k�d�w���D���j�v�� .w�H��zwb:$+Q�P�MyD'(�7M�g�/z/�9qRg]�d�r�-j����x������|��mj||�Q`W�Xˊ���7ٰ,��x=H:	SE�1+#Y�.�= 撗ǆ�b�E�/��2��.���E�Io'�a�N'%Zg��Ţ�� ",=��p�C�+�s���NI�ű|����ʯ��?����Ǫ��i)��s�t��H�����|��7G�P��ܳgϷ��-�b�x�i�Z�~Fv�q=j�.�9���̾�5O�G��u�ݟ������u�CHW�߰���^�~�����O�U��s�&�S}�r��~�wo����F��9ܬ7~�7?��|�k_{����A��&��LY�{e��Oak�����ǎ�1�����DX���?����D�l;?�C�&�v��s�m05"�`ǹ����6�D.�Z��k������i�����uu*}�����q�����'7n���ٳV��jm�J��N��Z�^�Өt�Ѡ��(�\�E�Z���s��-O�k����vo�!��������*�������E*h50l��5�G���������o2T_p�)�_~�y�%��Џ�x�� \�xN!��Dq�ʼ�AW:ұ�̦Q�� AT��!��ZR:K�gA��e�J,
*�%���."�ą�l�q0U��M�I���8�"���Qr`���I`:�l5��^�N
ܽ� شc�� �v�I@	F#e�!i�q�aff��=	{*��šC.-����Od�׉�P��"�Z�,���@UBf�ef����⳺�6� �o�by�N��Bj�M�b,��������<98�	��H��r_Z+�h�O&��+R�p�C�w`VaJ�V��`X���E.ju��tW���GxEj%S�+�mȡ�uzި.Cjrz��x�n�8�P'����KOZ&�E���"Dhr����c�ba޴�\��Qp�4�0"9wd���O���XI��N�J���q�o$S�@��u�i�� q=p�ײ��u�"J� �p��(�FLlgg:�h��?L��Pi��ڑIb:g��Y}���jod�2�(a���DY�ZKx���C
'Q��u�n�37�<t�Љ' ^��c��אP8�Oڅ�!�J�\Bە�=�'u�$1�H�~t6#gE.'�U ��� =��ol�h�
0�+�P,`�3U�"��P���q|�j'����U_� �a �PB�SBu��:��.Xn��Io�S�|),h��K��!�B6�-��zO���K/aC#��c>b��nxn�^�/�������o���9�a��S��ם;wRnAJ`��ѣ�G�r�b�����ӕo��'~�O��O��|����������'_lz��
g5��~��೎�܎R�$�\lL6����y�7��5����j��]*�h~�{��{}�c���Sf�i�pg9S7�5��'O��+_����zR#��OZ�i����8֦A�!��v�ڥ�}�g�K%(?~JO��`�ZCE�/i�~����~MSe�޽��W�&>�3lK:6�wd!ۗ<86w=�}�̙3z���&����)����+��}��218ô����f9)�s#��j��zU����)1�_�)�ej�F��z�-5��(׮]��X9�-��|[u��^p���$�Sf�.x�M�!����'~>����ug�mR&,�$K�c+9�x��"�h��D5�U�v�Z�I�+n��b����\�!�i�z���f;��ę�>ҭ�țgtd�p/�4g��=�UB�Ǐ���#�ǩg6X�anD�����r�B؝e���#Rίe�c�h�5�@J8�8p$�G~�g6�H����������a�F�m�5��E��n��8���K���)�]�fOJ]�t%����	�p|�Q�&N�3������oh�X|�a���~�f�WJ�X��������9!�@<�.�	�ڑ!7�;0����j�r:%�U��h{;V����S���>z�ё!�=�*	ׂ�'������~�>:�.^��1ڼ��gP=GF����?X(�i�Mv}j�	J�M�?_�y����٣
Ôv��-$��Áް+J�2;�Pl%��v�J�ٖ'a��$h�&ԂmM�2��p�`�O�hld�X4�eS����+
�io���lzttq@Խ�fT�
���nS��}��a*�W+�X�Z�n�f�NJ���f��u_�zYx���|U�Z/�e>��Q��K�:�%��duT*e?���ږk&��-�D2�^�bT67t�(�H�&��q�e �ϑ���K�wD�B}N�x}����r�彺��F�B�Ď�OU/~��"�X]LT��Ն�_���^�\��E$I�@+2t����׎85N���im��TH�/<��:VA���1��AK�إ�z7m�DXP����Mb(�T�Y�l�j���c���LR��FN>��8Z�z�4�v�ޭ���Jp� �3��_�������:�O���������Ο#�b�}��~Æ����'�Omڤ�i�;vl���h����/�<��|��$"�j������S?}��ɩ��+V�z!<�����q�Cx���j���*��:�z����%����P�\���x�V4�=��`�w���F�X���0}E [�yR{j݆��D'|�-^ky�e��@S��4+H�n��~/CE^5�7��j�>�eTz�{�d� @�Z#W ���ꫦ5�U�f�}�SSs�N�+�g���vj��h��2�ʳgϷ�t�&��MMi��<�xn�A��ux�j3;|��C�x��5��l,qn-=����
��z�� �]k�\"��&����I)̘�ŊfwZ���D��r��Nh8&��m������sY��0�p�95=[���wdb]
~db��jq�B�n�W���VK�����2��!�Ӎ���A�	��i.U,���B��'q:��0���f���%	k��8�ڝ�-��:h��:DC��*�b0�a�0�U/j�@��d�[.�
՘j��W��r�jB���'�a�G0q'�O�LI8�Gx�p��J��9<�Z�	k7|�?����B7A	d���X�X}��x��a�����l��	X>��%���B�F4�9��/@���[*������vI�6^M���r����S,?�HbR�A�fc��ukY-Z�W���?�	"8���r݄�Y��2�q5�_�"��T\~���}��}V�hȕ�ŤY�?��h�Z?V�Y��Z�O5e��/�T�dٴ��i�d�=qn!���E G�O}�S86�Է��UV�������U��ز���%47k�Edz����O�X0�,�ujr���GC,Y	���ӭ��� =N b߾}�j��@�d��[��Ǻ�{�C�8�!�A/�E�רE�����@m����,K�v��v"��)|��҃:\�ݰa��y�ur���Ĕ!��p�6ܨ����d\@A7a������F@�($�dY�������i�d<��9���i��LWB����qUi�82����@IAMU���O�<IS�����&DX1>�;�E�l*��zHX���:���R@�TOgA	C�����,���B�X���X�h~nndt���������-���[RuГyw��ׯ~�w�wu͟�94E�H��'>�rG��ԑ���Ow���?-ԫ�[�F������H2e�ؔ�^wE�ٵm��^xe���?��3��̗����~���2��eb�>ֈ���j�	oQ��}�ѽ����o��Հ��+��rO����c��f�D'|��L\3'������S�� �FV���Y�t��X�D�;2~��-� �4R�|��ɲeCڴ��
�xS3�nݪf���?�Kݥ����H�voM��%+ű����"%���\��>��̤����
�Q�`܌|μ�0�*�d+���c��?�T���}�ݧ�{��B�4�h���$GoKXq��;1]	���gG��;	��0�L���9�؂���LlP�v�7%�K��e��	�c�T� ��������c�w`0Gj�)Fђl�8� ̔��B�D�s��D2�	����:hx� �*K�o��\A���C��g���ш�o�X�wZ:'�-�)�]� ɐ]�- 7A�:<+1�^e�,Z�(�8�F��b	[gU�%�Ɗ`�%68��a�CP��������<����^<v��MK��L�Q Ӵ��B��05��0{]�l���=q�y㐙��͸�ȰSP�?.��'���&��S��\�����gRa�V.v����܌U��T���|$��c�V$���Q��!
�؈DQ��{&�ӧ��/�K���;�rՊkׯ��j�\�n�.�0�L��%���2����ӼW�4�\��c�q���=�d�i=EK�Yg�}ʳ�&djn�Zm�����{�)�Ѩ���p��A��ڀ�\�ds�+u���cQ�Y{�.&�H.�f$���e�!$�%:�H�Оp��N2Ȫ�����ޢ��P�[�W�����c�e�2� L8����C]���q��9�[����Xp�T-Mϙu;0<��u�Ŋ���nj1��-����&.�9�w���)	f�y�	�u�&�q����6�t�����9���)�(�s�[�ND�T��x��MD�06� �U
)D,-mn~�eM����~��K�ɍ�-Z�Z�ԫ5�|�FFS�Ҕ�$kAC����¤���H/bGH�E11а/N��O�z_S�J@\íFz�EK�zFST�������ꩧ8(C���f�:��ѣ����$aE߂����eV6y�=7=ۭ[o��;~��@�!�-凊�r�)�Mw�ܩ�~뭷�S��EI^�>ٶm%n��v�P;{������<�?������hN\���?���G���#�k��������[�H�:�(��G���������Cx�������_�mI�zz� ƃ	A{�ȳ:�qĒ�;>>N�ۑ��z[/Kr�Z��Ru�s����7��9u]�V�����ng�C��<��c �'NX���e��{NMڵk������C��@E
�,9���$�8�ۉ�����w�imvT|�q��k���C���5���+�t02:t��	���5+ϝ��6�l�UǪ[�մ�q��t��ժ��7v���hOO�y��ao�z�܌qT�c����7�T���F\$���$䃒���lO��s�)�_�ҭ0eg[�}�6�P_H;�b��L\ �{t[�=E�<� ��P��q�D;\��T�M	�Ȕ���SJ���.�ҦR��j�F����D픹��U�'s�0��^�B�S�2��J�@~����6X��~��=�QY�w���
P0���_\��e,	zT��͜8�j^�^li|=���|�c�\����^��L�ё��כ!������<�/����q��M��i�@p(s
��`ҟ�D�b��ɓ�����X�T�5��6�t��FD/&g�nN��n�E��%�NF� ����m��S4���+��	��D}X���fl5�Y�,)���(25�-���Z8�4�a���6������c:��J���;��Z�/�P�c��?���+m,Y�����	/��زeˊ�+"�RB��.n����K���8�7ǖ�����ǩ|��?x�(3��X�槅�]FѦl=��vf�w���t��)��'7!A����x��\Z��B�,pHIփ�-�S�PWh�pvB�ґ��_7�#e㄀��p�����Y���o%�][��S��:���g:��-=�T6O.�l��>� ������qn�IGmd#�
2ǡv� Э�=k5����Ņ�?b���	�� �4t䉼 ^����}qǎЫ��|�KwcF��a����R4-�ϋv[*����M�3�]t�h���¬�F��z����e7�*�cљC�ES�p��4ݙ�Nnͻ�;�$�u�f�Pއl�������:�"���1����n���w�^vp\���+��޽�YG�2Y�|ug�J�Au)]z�����Q��/��D�:���pj�����ANXJ����sR�@�Lg'��CD	V��6J��M���Z��_�|��]B����'>|��&������B5�7�xcN�9�`�~-g��Gfg�0".7�1�=	�ɪL0��	U� ׾}����GFص�Nrr1�2]�wѰ��t}ʅ�u4;�Ո�٭�i�����%]��3�Ï$9�z��.}Q����Z�s�����рe"Q#)Hz뭷��ZO���`O�j�
��j%;��=|��uj�M9���~��As���W�q�ϗ-�dd�KU��Ǳ����C^��CC(c�{D�W�+�%7ܰ�9ƃ�B5ێ�W��b���˚l�\ +���>C #�O�]L	�MBT'V�����4̄If(-�H��T�D�\<�u�e��t~u8p�%�l��RvZ:��Vk�W�Vy4����Zb����-�=�F�����@O�K��<:��E�!��2 ����,y:�]L�Q�u�	"j�0i���ϐ����H��,�E]q�+��b48�D|N?����l�4��	R,�S�b!l��C�0| _:N�`+ �ҍɟ�S��ە�pk�p܇��� ���/��X�{,�+����c�O�6?Kh��8�1J�A�?~��?�o.q��s]KE��\ �L�,�V
YG�#C����bIذ��%9u���)��@u
GR��s�Ozm�Hlh��\�۩7�^P��Ɔ�-ߧ�X �઒�u�ւ3<��5�fs�TJ�\��vD*q�����d%���X!�E"���XcLra�$��$�ug�;��Fۮ�I��ꞞV3�]�?�E� �լբ�I0?�8>��l�0HS��ki����2qM�-�!���Y����o��,�߫�I�\[kr���KP����UИ3� /#�~��A!��x��u��!=eӦM��Z� ?�^�7n���(>Κ�	�@��(�U�+�U�n��B�C/2꽤�ꌁ����蓊�r�+�k�ɹ5�/I����1s�[-�1�i7oތ#M�������U���ק=��%[?\CpP'7n��ш}���._�P��iW�4J{��m�:Si|��97��L�5kW�w�3�,�j��}�V\_-׼`B\FXG]���~���_��j�"�3�P�;a���s�?{�"�P%���� �ҶV
�tM��o������B*{�=���{��A:Xcꞕ:�s�|���$߿���w�9��nٲIgI��{���[�$�F��s�N�U�AT�Vz��"6%�Ϝ9�)qebb��oC�k���aM&�^AHB��V�𙐖i_��;~a~���_	v9�хB����.3��_ԁ�Z�#N*��>�|���-�/�Ũ���,�%�1�5�S��\T"f�g��'�E��#��G�j��*tR=l�`�\����'�|���75[��j����z��1L;]�����Y�Ic�r��L&LG5�_�|ｓ�]�AbFυ��X^X(aR����G�KL�#B���ɴW���!%zP���ÄG�$�gj;��bk�����f@*4^��0h�	m`  z"H�N�t����J-���;�С��DYǃ���a��Q�\5ԕ
5i���v*���Y��L���rqtB}^
���XƂM/q���$Q��M�5�����o��vu�����L����d�t�h�t"��h5qn�$v)�&�tھTO�� n����d�k���/>���u@���G�9|y_019��B�Y8ex`VۤA����Cr
ÜqO_
�	�N�ٚ�
)a���+"KFS1^g�����-�u�`��%g�T�5�T��1Wl�V���v�Z��X@�+��㩻q0��2v;�,�|�S��B�:�V,��e�س�kB ���Dŋ���:�G�`��+נ�@������ڱ���w�^��f��:�A�2���c�B�����_/�lm/��g\w4�
���t���Î̚ŀ�'��ru�>��Ո'/!wkY@����]_�V�-�1�<�I恰#�Xw]P�<�]{�P��Ήc���ʲ9R�w1V0=ɖ���>m�vKiax��q��no����ה�1�s�5��Rڝa��+��.	��@BcP2[M�
��Z���o۶-��}��������{L�ӳ֮ZC(p���TBt=�����of��\DT#%�r�d5����8`��2��ݓ���jǖ c��/i�xF��̣&!*5@@D�k�����y�ֆ-�C�@}E�9G�a���cQ����5E*����I�ܾ};�vI�3�
��1��vó��9�#A�����~�3�m:�5����]�����/���?���Y��:S�L�CVfq��]�o�:׊K�B �Gb�!���>���8]�6M!_�X �'��8+^�ESE0E`T�����gz��1(��R�A���4!�Bn��V݊�l��`����$-��o�����)^��X�Rlz5�yzj��+_�RU=��N6�W����������+�.�΄�g���[���cc��݂e�w�@� f�&���M'��y9���4�hė��}X�Q�C����P����[=z\����A��d�S������EJq�bW7��z�֝n��;�XڲS|@��F�'�nK��6�L�7ӑ�er�$� >��'�W!ѫ=Z���r���0LL�.�" s ɱ�ZB��z\5���uZ��:�-��%r� _�"�<|&�jR��
���Y��3K�cRq*�R,��]�ygqfΰnu��\�Rg���� �}������s�ַ���AU�N�>�%����?�svQ\SԹ&�Od���\D>�	�d�qުp��KJ��#	4ad�5�h$N���\�D�\���&�tE���~��݈�R  ��OM�� @?x1�J|�n!�� �k�f�Y�8ჃX���7���qq&'{&�7,Fd3|&�Yȃ^�[V0���2�j��<��J�Ȼ�c�Y2�_Z&��;hC�4ZK9+Hkɳ��l>ׂ3�+��x)��hG�}��P���hSPo���i�P���άM<���{w���|Zٔ�<��g{{�5��0X���!�(�45>�S8���'a\[6������I��q� ���È����������Œ���t$3�V��W`gT$5(��?A:�#�|-���������ޞ~��eu�s�c��'��x�u���3��Ԥ={,�`���z����Kn�z�SSe���}���ZE�C[9�r������c1����;)E����lV�up�T���R�:|���dc$L&MTܖ���wh�08ѨB���2ݦS�(U�3X��L̂�v�w��Ru�K��?Ӈ�EoA��j��(���X�я~�Rϋ�M�
����q �+)H�S.16�{�$���z���z����^�k��g�z�!�r�$�o~���_�mI�+�8�N�{��M��y��4�庛�H�LMHf�Z]��
��;h\ [m�"���1t;;;�qj���,�V<if� �K/�a��Ո�X��>} }��7iR����_=r����jP�X�ٳ��h~\=]�yc��=�$�,��2�vm���m;v�4�x}$�Uk����7u�;�d��1�!x衇�K�E�
�+��7�T�_-r8��~(Y ���^����p߾C�_��'Nj�Y8����h:��#
OHݸ�<�st[ݜozW�RcV�>!G��q��Ixƨe"M'l]=�+_��>�ޱw	�az�F��d��:�0��8��N,��w��NM���#ۉ�<�I�}8_��>q-hG�sW�j�kx����ڞW�;�4���	�-b"MhOq1� ����R�T�ȩ�́���� �U���F������;W�A���-m�bo�:`B�J�gQ,�8�R��$���l	>�ܥ���-q�d=c�AfI1%~��e|�t#.v��NQ��zvV����L#�z���ng�~mbr�d�"v��'��Ǘ�M(޽�!^�:鐄���Վ�H�!�_�����#7!!���$B�+$ԝ(��o������)q�p���#�+n �ht*���\\e�'���ә�&�5��[�3ђ�ޮ��v�0����2Q`D�q�H�՚^��(��!�$�RS�"��p �n�D^3`)n�$��`6�}ѠR�Pg�^A�����ȓ��|���A��������PK�4I���6�8�d��q�y��,��t.0"u7�k��˗.h\GXr6l:<�F64�1���ҥ+jj���8��]|�͸�q�bK����a'��8�گ5/<�*�$6��uݟ�'{b0�8�u$A�����;�����+��LM� c�5ې�������^��cbr�y��(������N����^��b+���?�t$���+�8#�n>~���恭����f.�>�8�|��������o�'b���g����e�r�c�0�X6-W� ND��6�$�Nr+�m�~�U���
���i�d��`��NJ}(�����N&V�	d�mGiK��5gI}����]�^7�<5��̄�ѥ5ь3��\��;���߰G#9��B`�<	Լ�Uw�.��w���Xr(���"0��:�AZ� �nK����z[���vs��Q�+i>���?=p���>S$����!��m�ݦ_֯_w��e�_@PP��b�l�i��Yk5��'�t�KQ�)��]�f��*W�z!3�[�d���;?jĵ%,�V��y�]?��࠱ЄP�_0=�z􆠏�H-�`���o�]���O��i�m��t��Z[j��ծL_M�S��֪=^�̳��oP�u��c���rsVU�װ2Rd��2�`�?��R��l����ʕc2!x��"*�2UHB�S���<��T^G�F�S�1�5�d&i..���y�P��S�HDq�!�B�6'!�hr�ȈҦ�3��nV7+�� N�K���b���(���l-�
��aX�~Y��f�a�c�rc+�k���Ř�j��h�P�Ӓf,�f�K�gəڎ�lJ��Y�k-Q8ðញ���c}��*�Y�f
�;��=�Ψ^ylٲ�력�HB�o�����F5s�"h D'��h"}���A�ƅa�P!�g>��j!����|��&�34�Tgb�	��'ľ3^x���[!"-����u�L�4Zq��l����/���M'A�"��!��pF.�lu�i�:��j��2S��;WK�D��o�m���Y��|M������:)���4��B�wӲ׎|��mɉ�5�E�f"^鬅-Ҿ�#g�*z�}��D��@N�.��K�j� ї�U���Z��'c��5 v��r���;����B�՝H;����JȌ}=�#� G�޽{���/�]��aSݻ���;S�g`�SŌa�i�hFD�/�;A;���a3a_j�e�?,���Cv�:Eڼv�؁=V,q:���Dt(j��������6�p���LA���W.^b�ck�|��C�YC�m]�(���w��i%m�[�S���SK�V�)�g�I�=7�ّ0�����V-Wj[���s3����b������:_׮[�B;.!:��ͲS	�[=���=��hF�C��4!ї�tw���Κ}S�u�p��ba^v+$3��Ig��T�$CZ�y���2^�}=��U�d�y��f-�K��v����u�n��,'Q9ݓ�`M�d��s�&�ƍQ��hꡤ& +��3it��7h}c{X�r&��`/��ҡC�ڱ�đE'�b��z�]�v	�$-	�.���'�x���<7}����n��,�H}`@�c�ٍ��ԧ~�W��`��H�%ŗ��4e>�y˖G}*��6�g��Zn�
E��LT�4#o�e�ͷV�-x~�x6<��)ՒR��:%N�0����R�lT���6��nnڔ����0`%GsV}�V!A����?A^-�}���r�5�u$,Fߘ���8�*��_��_�!�##27WB^+eܹ(����H|z���/���1��[c���	C�;�S�=�)�A�X�纈���ª�Ԇ���x���\�P�Q��]���Qz���XX\(v�0��0�?�D%���XQ,9��ƪ:q�L����G����L��� zH~X�H�*��/Zy_�߄];��r���+���l|�Ɋ�+jv�����:�|ZK
�����f.C焥�a.���N���@7Լ6My�E���7t5[�m������}/��+j�:����=�)�n3�^�
��==�o�b�j�%�8�Ø?�_�K4�8j�$���t�#���m�T���s7c�qgLŅ�����X��i=�mt<%��� ���U�1��It��z�2B�+�:ө�l��`I���T�Ij��$+����N���t�ez�t� �Ӈ����L:V� �T�`�l������ A=¶8�jÆ�˗����-�r�T�:���g�%� �$��l��)���-:� M-/����9�(���"�M>�pԹmgӞ!��o�  -�h�)<w��C��&�o�[�z���'�Y}N���c�p1f]UU���8��`�`8cI�$���\�l�Ɛ�?hy�`��Ex�e4:=�i���蒧�sh޹A"����5�swI��3>66Fp�F�w��׮<���.p��d��j���fu�+�9c����¼�?�2"-��_�����a��bQ���5�k���4�l����dg��#�˺=�͐�{Ѵa��K~qMj?�Z�N�����/w;�O�V�cu�_�́@ɶ��T�ĜJCγ}!c��Λ�q7�r��O�l��u��Y�Ӊ`�Z���'la�&�M(Lf2����sO�:�1m;��&�`@�V)Q�8 ������|%Gq���<�6���Q]m�p��x1�>� z]�Fd4�ockص�W_}}Ϟ=&10@ ��V�"�X3ua�K�.i|�\���'pᆃ���tݾ}�f���V�+��"��re��&�b����O\G�WK�jUe2h�!jB.zJ����8W	�1}�z�j��\r��Y��X���g�}�^�r��cL-d3Ѻ;{�L��˪W�Һ뮻z,���V,m%��L6���.H������x@�;w)��ޑ��7�p���<����k�\I��j�/��/�|��3g.�����?�C�"��b��чZ ��l��ꍇܭ�i���?�#}���~������׾�!����{�6AF����7�H�ui7m;j�>����8k��֫	ejj�<y��ѣ�`���D����>���q��u�������@��� r�j�#G��8��89�4��ا��i�S��I<R ���5��]�\���k ��>s�/8f������G�cQ�.�RL��ǭ����+hsĆ�
~�`&~ǹk�¿�؁��(g*�K�H�Qm�R;�����կ~U���7�	�����Ǐ�[m�th�Xa��'��D�����J����C�א`�㔂��?�e\��N?v�~�7�/7�d]�NҼBc��A�ǿ���q�h���#�*Wz	P���l����$�#����\:N�j�:��C�>q�Jp�-н�1E�͠h�i!�����/�{yn�A�=a���]q-����A*�TA�;�9�Y�m�2[�U�.�
�]6�[AT�֋�CC�S�R�f��|!JE�׭^�f�L��W�Ԫ�rܦ�ͳ�צ�J���f��5C,,�b�
�I���lu��t~h�`z%�؛n���VkN粫,�	�j��LOW��ך�G� u��9����l�ˊ)�Of��8�O����GG���.���N۫;���R�U+��c㰂��*�F�53=�kƖ�0ў~
�����#�	�V�����C�}��7���Aؾv��m�.]��[bf2_�^�r����=�{VmjFA�:O @(Ah&O��a#���p�N��ۮ�4l�'&�*���&ғק|)��ͽFˤ�k����c�L�1�,����1�,��<�o�ަ4��̤���iY��j#��np���Gr��#�
κ��}�]�ߪ�M����#[�3R_�馛X��g��� }�w�^���ZȪ�95CäݟD`����~�v����ڤ�B��]��\?�1Dl�!��y����t���O���ć6X`�����[�\3��L9�]�v]�vMmF�^�h�߱m��I&~��~���^��ɤ(d�~�듚�s���\�Т��g�U�E!���X�j�:���3~�EnUO��s�O��իW���*�+��������u5I��&&e�G�Tm�5p�
�4]dtt����w?�I~���F���G\,�..X���[o�U��Zuǝ;��	i��ʢK�h�]��n�l�[�����]3~����C��Ϝ��u�����'�m=w�ネ����׮>��ӿ��1?�����wY�����y�;�<w�6A�D��H������]}(�q�w���?F�s���;v<���<�f:�SWL.�:S�mۦ�g�f1��)S�.b�_��h��\r��ͫ;�3�Ԫoׯ_Ӊ��'�'��޽k�0�Fs��-B�z�&�֭[o�m˯<������=�ܣ�)���#Mg�Z����5ٮMY���᡹�ų�m	�[���wߕm����ً�'qΙp�F1gf��믿��u��'O}F�ܗ�p�����o#!�/����U��V/�z����e�|��|r����-+��2�r6�i���f��j���j��\=j����e3�FՆ�j��F��S2��|�ڥr�U�[�וF�k���9}E��FP�X��^
�X>V&]�iJ67Y�{e�-$o@r��X�7΂%�ٷ7A�Zn��U[�#ۥ�lf��kjE�\!���0:�Ӄ�8�4~����hiȿ�_��R��NM}��v����G��������ukљ����G�����}Q�s�#�M����c�քA�H�z�D �pHh�:]�@�1qb���E0�]�y@�x�f-��@kWS+��7c�Ғ�6RP1�� &.+\�8��I`���Q����|U��������xX�f�ʪa:��e�ڣYȪ����xH����mKϤ u>�M�2m>�i��j�J��)D屸|i����ٚ7B3۲-RO��hD��_pz����[�ڊ-�[n��Ź� �Ln�h����o_'�ƞ 6>�4DQ��I{q�U��j�k�TP���N��~Nx����HB�Y��m,�Xu��#��H�ʺ�B II�}*�8���߳.��X9��%)Q�	�O"o��uR��g��@~-�1_�����+��vڽ�ޫ3�d4�PO���[���6;<��]�|���6b}���S>��O�'O L! 0�s���t@*S����+u	��:�����7���iIﾫ��$�1Z��{ɪC��F�,��:tH����"a,Ѯn߾���8�úF/�m]��뮻�$���6m�� �Ĵ��ս�+ɼ��n�.ҝ�6\KE����������H��닰>pTp*�#�/r�"�&}�+_2c
m޼Y'��s笪����6��ӂ�������5[�U���[�^�׎��i"�[e2)�%��,��	����]����,=J�Ix!Hm�8qv<��3=˦�a�#�}�ٻ�[M�B�M&�n��|�I����v�DM �*�M8��O�z�:_�~��K��U���	��o��t�;���멓��u��:P�W�W]�I���ׯ_��O
�8p@�E�#L�]n��}��i�rl4�R�������~�W�NQ��.�ƨϵ����_z�a��l#_����XJ;�'�©�'�`˵�S����ϱC�%b7�a<6����c���7ݴA<������������[53��^�D��wEP�4��W����?��n�ݱcG(ͮ����~�:M�(*��l�@��F);3�Ǐ�Z(-"���$�[m�<�'Y_Z��g�Ϋ�IpxY���~�e�Q�t7���?��@���('�xP:D1��_m��x8�d�|A�J����&Q�+� ŏ�Z�Ҥ�mϞ=�YPkv�.���`�s�c-=��j��O���?���a6�Jr�A���q�q%."����+���1K��7N�Q8���o�/�?k���	����B^��؀+Q�F^$~�v�����E�J&�rշt+0S��Y�@K�:|	�\c�aG�M�<�'���y�������B-��|\�*�s,@鸘f#��c��$p֎ӴA�pW�����n��T����05	^��"��A�%NV�άK�A2I���Ǫ����\�!C��A��A�l�ӧO�)��=γ��Qg�$�t�����mb��P�/2)��L���@�_�*���.�O(�s&�g�p^6��#�M��Ѯ�ŅĤ�H�E��о׊xd��Uύ9�J�]>Gi]�Cy���u2�p]9�+�S�ޔ�����k_��N�Ȕx�ƴCQ��5/�B�Fe�M�����T؀�B�ڦ�&S�-F�,ݝ���ә9�X�V���z`Í7D��X�W��a��i�L�^����v�������ۺe3����}�s:0t+�I��|�;BFٽ{7�Y=�L��,��[���z�;hvi�����5Ԛ��#B�WFY@ç;���	޹�����ѣj���Ձ�KQ\�_w�}n��v c�K8`_���Xc�Q'���a�KTv}5^��P/�P��4�W�by�:�u��/��Q](�N��Ѡ�[a�j>���;o��_s?���X'����X.�9rGt��u�7"떹��
�S��ω�C'G2C��.5����(�jL[��
I(S��Ⱦ�꫑��s��W��d{��և�i����~7�%D5"�^z��u;^~�eԪ#_5H�Ѧ��h��@4`���Wo�\�b�[o����`<�B��L+%�H���,Q?񤄵t��qxm%J�w{�,�r��Ԕ�v4��-���ȩLy�U�~�=�$�uus��UZ,ť]�M�˗����<�f�c�a�ԃ�Ԍ��P?����� L�daD�RM]��mg�C��vmB7ѻ J�jWGs�3
a�����a�v�����u���u��I�և��k�s�k�}��*h;\N��u���p��[G�I��b'�gF���q�E�d�d��e����_��_	�Z����b!q���/��K=�t�8}?�k�k�@(�l��pr$$�0�ӂ9M����x:�S^X@�o��T\�vҘċ�;���c9��p�>wgs&Le�α-�B�W��شa��?��?$�ݨ�����F����h�eq�9���W7�\BO��F��H'透�kƚ�$B�v�VhB��i)d$�Hz'8Pfi���v�7�␸$��}�o����Pi�9���a�@*㒉{ z��`��݇,�l\+Da��e��f�*��k`4��C$jQH4����E���-�cL�4�)�ש�iA���4vC��ߵ��={^�z��+�'��Ը�;w�D��/�(� �r��;�v`'��u�%�Wۍ6�G�B`�!�Z ?,u�9
D�����Yu�z8��k:�����	%��Q�OϜ���AB�D*�ש����'�4s�u�9����P���8�F�Q_�������C��fa�u�L�$�;r��e��?]�$�y���ݹ{f0"�3�	(��)��L�Ȗx�T.Q��C�t}��\>�#��-�.�t�p�@uD*�2I� @ D&Adf&wOO������a�5�ٽ����ֻһ� ���`"�+�2�������-���Ly�}Q��{��x@�Y0ejv�@a��Ո-<�#�0��.�*!+��u�փ�a��ԝ�µp�ZS(:	d��-��� ꕥ��$�F��D��(��&���^<�����L����#kPwЃ�J[�PEø��L��H}Du�6���x�o@␎
�t�N!t'�l�?p�S��������ժ�9�����B������q+e��ܰU�'���В%��
��i-�.�]�R-A�[�}o�r\���I�Ԁ�,���
y���f �?����DpK����c��_�~�G��3����],/_�x��Hd����$�[5_H�֡�\_O=������1�|��1�.u����Y�\�F�F7xz�7J�
Dn�_M,� �@(��x����w�]ccW���р�g��Ġ��B���F�����G?Ҝ`�c�i���m���ر�h�N*i�z�^�c� ՞i�B�?<C�A�R&DE4�@O�{�T�?�m"=Ks�ұD�Մ����F�!��{�[dJ�	>�-:�� �vv�Mw2Y�q�p��}2�mX�
��A�=|���54������akx���z{�K�?������H�%S�w�ߕ��-��TA�RA�3Q�;>A3�L<k��fTi�S!�h[�Z#�����B�퇆3]�ǖ�vsJ"
�d���G$�v�3�g1�=:A��+_GoI
d���]��p�h��mۖ8��fx�B6Gݮ�UM�j?[����Q�D�&�F`k����\]w
t|��;%��4Ҕ�C���!A6h/���)R�B�����8�0�ٓ(p��҉	�<l!`9S<"Jv�����q� FH��y(�(qB[I�H�V q�t�J��č��I�����R��q�t�vr��,�]_`�`�����g�b]+�,����ٿ�n��`��S��W	��+W���3r��f�5�K��ɻ��=�'����!�	�w�y�J
�����q�l�e�'?�4hl0)P k��h�v�M�(w�h��;��ĉ�ӱ��j�-\�z4�k�5b�@�@��ӤYx6&F����ڑ���խ��
	�y=[S��[���ka�����2֒l�4(kC�֕p��![�F�5z���͍���M�j������si.+Ȣ��u�=ܥ���u+z(u���]O���֕P}j��F,(.Cxn�:Ri�gti��RX3z}!���f"1[^��PR�Qt� i#�P��>���Pi��w�6S�6!�N�����V��&�-�e�͏`"�Kj�5��b�C��U*"�AA+���7-���c��JC#;�9�
f|-��c�@9����s����'x��cl����AͳΝ4�v�Ǆ�U�.�]������k��+и�j��<�vA̿��cҒ��L��V��s9m�ROw�l?��CHRM�ǟyb��sV�ԡ�(K^`�7�M��}�v�%~e��c�.��Ѫi��=��C�-^7��פi�4'Z��;w~��@���;����j����I��4�8��O�8�G����P1:zI���߆���t�AR�E��K/���޽C�����[	�k���t�>Y�ve�٢��j���\un��駟&�Z��hѳ�oZ}3�ƂS�����ne��0@òK�.�u�t�v/����Eb�ƀ�X��8�u��^f�V�|���D����v���;�A��C=��Yk12��W'�<q���v�F���d�>}�uӦ����B�eˆ��o���3'OQơ��ܹ=��m��LN�pXR���A!Lb$1��׊��\e��u�@�JԞX����XsG<G�!{��Xk{&4��q�б�"B�W���'���z�;��]���l����T&!�-�<R��A�������K��r,
��r%�q%���I9��N�� �a=��0.�+Ќ� r�>��3 śH����L�a�K�Ϗjb��0��4{U%Ү�S�"L5���Y��4B��z��[x�<��T�^C�(#@��i ��-�(]y�'��OLZ6j>�o͐}�[�a�gE�~�Hy��K6nѰ��c���'B�/���|ہ��X�M�Ц��m�ƕ$�D���M�}�W�܉�S����_$!_pHJfA(|���T�7��p��&��y��Z20Ļ��KXoʒ����ޡ�M3ы�j�08�T�OMY�>Tp���� e��+%��Vټe;�۱�t���I}N[q�$0�A2�%�%^A���Ÿ5�Hһ������H�a��ڬ������E������Du���2l��Lw���6�;$�&��n���w�"g�գ5<�u�D�ȳ��C�K��+����z�%셺��~ٸq���K	�Li&)t���#��ס=���/�d��*�;jY!b��;��)�@�I�H4�4L�5�3k�Y�� ]�BH����.�4=H��g��KJ��N��Y�R�<�3P�Z�����Ϩ.��M?R����t0<}�4�\7wAd���T�@@�j�����$I-��F�3���^Y�z�������#p����zG���g?�ٚ����H�"z��6��f�E�=�\��5'�7opF�@(:�;z��W^��N+�' V���p 5��{zz�}�Ym�m۶�����ק>�)=���_{׮e�]W����9�%(]�����ab-��x��c%F�"� ����:�>�����������۷֍��17����^�M*B�RZk�m��$&�ϴ�������{Oh�p�bEJ��M#��3�bF�;�:��I�C5��Ý�d�8������ۢpRK�}�f������Â�[/8Z�zu�ʥe#�R�� +W�z��={�譭�*�$�>�hڽ{��g3���a!�o�%d=�R�fRJ�t�S�n"�91$ /:�m!�>���:�����v��P�����#r���M���7���L`)[l�_K&�G'ɢ6���$�@6�{�HY��"���nX3����P�A�Z���1�U,�EGU/528Dk�Vݞ�5�VD�֩$k�+i���\�	8x_���8��>�8�
�@!��B ���j�J��Mp[��T(ޒ� ��l��`k��FT��ӆ����x˖�1N�L9Q�;�\:���z������Pi*X1w��k;~�*9�lO!I{�Т�ӹ���ao]����5�ɤ^��i��9��Y_��̖{󂄤o�gu���g ���5�K�C��nGf�6�Ec�U��@T�9�;S��h@�ZĆ��&`��ON~��h�%�F���)�=M&޾�15XA��U!��m{�J��WM�%ac�Yd�{��x�-��)�z}�&)�Ao��ni���t��Ԇ��;����,A�ӿ4�7�|�pO��
ґM�V��A<nۂǓ�����h|�'��9��z��Ԝs%Ć�&6*�3�1���II�˱c��QcO��R=]Ӣ�����������4!0a�p����Ѭ���u���̍�7>�J�6ڴi*����댐�,R�h��7��<���g��[O�U%%�7=��Dr�[������Ib���^ib�*B��#g�1��ɧN٫���ZDZNY�v3�慳���5�P?s�,|�Q�]�!�t�p9|��U+IQ"�*���ZrW�����0(KӠ��?��SF�u���5+ex�9gHWX�K%0P�ZS=E�I�^��O�5��CZE� @F=�裐�&��QP����z��H�?�sg�j�~��|��'�{�bQȯ��w���7���!���J�����q��y'�ki)-��V�vq �����sZ�IE9���/���R	]���67EKh)�P��u����FP�V�`ƪ���&azݤ�}��_k�����4����K�I��|�����K;v�<y�֌h��Y��]�vF��&V�z�k[��ZC�l��3h�I%(�+83��	s3g�,�ͯ_���:z���7;z��̤O}���;�T��v�ET	m7���ّw�k�����' ��7�Ď���U�4�t��:Y��|�Mӧ@T�Ѝ FHq$N'��Y�ط{q�X'�.ɤ�ԋ]eѥ����33W
Eu65oM1_hy����D�����Л�4�����l.���;k�s�N.�0�N�~��QQ�q�l1�if�xZ!�@Y�O�E��~��F�՗�/a	W�K;�K'C� xHHM�l���l}���p��#�4`!�e7Vy.^g��I���U�����=Q�MBk��*��� �� Z'1��H�g��A�?yBl�L�������$t��4T���`v��`Zh��E�˙k}�|;��6L������z���d�B�O�X4Cс�=��y睛��*Po+!ⶬ��n�^��NQQŊ�� ��v�rzƔ��fh��.u�u�>�˅�.:�P&�X�;ġ
�� b�Q���M��6����S�<'�[I{ѽ�I�hQF�Ɂz���:���2urt[8�(>�LK2vI'uCoq�]w������A[k������lD�\O���>&�"�@~�
��ŚL�-i��JSO]G ���/Y�"qG���[�ԋ<y�P%ib���!�����2�Ic�5!��5��Xӣ׬YCG#��50	t��4������]��9Z��'�s=WST�x�D�s'$�$�k>I%�L�c��,	Cho�]�J�4ҝ�(Z�x�;es��z�u�䫑'�����n*��^�"M�z$\����i�#��a�JN��t���Mu�^p~�����!���7�x��U�Zm?"�o���'?�I
�2�(�]��LuޛzF}]��O<�������|P������w��^3��]`��#~�ӫ�w�!�%0E��^����A-6�f��^�Pй\/5:�����������?��^z������C�����d���B�oi>��#&�FJ�-*��m۶GyD����H���c��1��5�Ȉ�/�haG�?P�P`�f�/��/~���y	�坿:���C��v/.p�0�o���H'��[͕^6�5::�	T���x`�%��[z],;J�%�w߻�æMw?�>u��U���H��S�^�^;mժ5̪��79-���� �)�-+4����J�+����w"�H�cҹ�]Z@\��P��ȚM��F�)�.Q���)y����.���+f��'&b@�+!�"�ؾ�Z��$T�v�]F�ť �EL��40w�X;!�j�I�����_�ic�v+)sfgfd�<���ر��9[�j������]�b|�VQ��J�qU��}{���:+V\w���Rh��s�~���ʢa8}�\�w=����eί�n�ʕ	TO6�rB�08�uEȕ��x*}:==��)p����v�'�&�;�HK�M�4�K�T0X�R)y��3=ZB��ŅF=�]���촍�9�͓��(��������l�Н+��N�t\�<T��+��,S�#�������}�\ZTh���zm��e3����9���Q9����0����������@W+�" j��YCr�_�k�����p�W.˶9.M�fĪ}Õ1+�@ȒbL.��;�'�� 9��Nk�;v��li`�)	d�̢$Uk�gix$���h�0H�Cɦ/!b��7����.mG/�c(x���h)H�Td�������$�䙕n���ɉ.Q>.7sU���x��ΓЭˤ��jXwJL��,c�,������ّE�����eCpN0�ZY2��[�n�:�g�!�&��N*����j{1=b�3��8��g@L��<��\j�n��s9���O�>��5�[�h:0&�ͭ���B�	a��*,亞<6�/#!�	�1G
2�c�u���C��00M4B^���vݹs'>�$��l����W�B��	�s�w�^)6�\{ijz�=og����B���io�LLLj;<���d�hlڨZM��4z6���&�����l����z;}��5;������{{�34�.��������:ź�o����WQuW�.���
M����������vP̀!=���*�w���~�[����CC "Q�l-���{i;0�d` ���k��'�'��R>�j�����|׮�����.�r�c(]mm?�$��WZɰ�oho|l��U��������x�F��_�fx��8�@9��c�]�i� Y&��l9��;�C�w���<���|^���@ɧ6�U��C��[;I�L�u��YԘP�Ă��w�٫Y҉��|�b�N����"�I����w�!�V���Z��s������MG���tg�GӢ_�|��
 �)��/~���4�㐂z��9���#%�"*	�m�@��U�V��cl�e^��Y��>�x�玫��xy#�\(�I9z�lA���f���{D@6͹#�Z����_�'v�4<
�Kْ!)�d,|�α"�Ŭb
���_}��k;���u���_P�щ����C�7�om������@K�qXꮬ��3�&%���@SA�eȕ�ű1s�:y��y������GF,�7I�NL�x"��S�,4Z=��&&'�8�f�}�L!8lذZ">���Yeg"���GFd�7H��{�H⤅�j�ݭ��
��lul���{ĳCX9�V��1.�=I�0}h�&¾-�5��Ԥ��L?N_�e�m�iN:-J_��)P�a۵έ��=��.���1���瘂v�M\�;�F,�<�ljP��_n�������]���w�#���D�[�`��g])E�[��=%�Y�P����ź��-m���q*�w,d_o�[�uo� ���I@G��X�NRCc��I{i �V�����)�X���+�Z�8�	��$�(�#>x��� 
�QM�q��󒶺 &��s�Y]p��!�r¤������=-㼕��y��Pi�����8�'��PKON(�e�g�z�)�����Scӻ�A�ّ�Fn/
szW��v�I���k�q���իWG�!�-�>�;	�'VY��킌h��mBT=^�Jg@��F�_�D���ظ؇#W
�N`GP���t����ڋ��~�zR�A��n��-�>2B�̒�^40�.���^ᨯoܸQ���n�',�� ӡ�۝=}* I{ð`�.`w�-7�w�}Z,�Ib�m�qa�Ÿ0M5$�56��_��fj�Q�����O<A�0!6���{�ܹ��A����3�*.=�_�{���-[���ز�&L$�r:�4��'O�E0�����$wo���ЧF�5�[mo/����D������jA5�^�رc�Xâg@%���([zZN�á�:?5:�Wh�8�+ut�F������u��E	�z��K+@����~�3���>�i��p�&�C$rAB�8?�dw���b���w�{耖�¾�ر� i=H��iH���ݢy�u'[�Z&�֎[��ӗ䪹�'��Wi{L^�@��\�d������Bc2���OfI����@H��iQT+!�{��{�Z��կ��o:] �`_+0#$����0�ِ�~ynK�QⅢR��TĿ����O�p�X��=��@�@���_�"�Ґ�Fd��O������߅�zt���c��o��w~�w����<�[ƿ]*9z�֛�.آU_ TW���&'��9��ڏ�'�Hr���֋�� i]"��Q�y�$�?�jz#���[�.!ĩ��|��ҥC���$�^bP�Eg?e�Iq�T��$�k{��f��&SDc���#� À��ؘ���S��i(P���dig� %��x}���P�e�E=ʸO�[���Ṟ��q�d.�m�$�Vhv2��˥ݞVv�$-K:ew�	���N�d���	 �������D�ҥ#�r����, � _�z��Ի��G�o¡�q�$U!k��/H�G$�Ȉ������Jk�1��q����5
��x##����0��ȈNr�D�!O>
�KPκ��������gƆ��j��ۅÏ:�Z��4��> �&ℌ5)
p���%��h\S3չ�˗�'(��&��T��p�z#���6]�{�j\���&,H��櫒�R-�2i�|�5���D ��K�e)��fy5Gbл�Is�9����g[��O!!�K���&_c �P�pV	�P��vR% D�O�^@I�s)���@
X�Z^��i<z�(1Y�U�������x��0}�tv��tjd�`�?��X�c�v䋅F˚p�b8kts}K��po�l
�E���$�L�������shƽ5��-��	�����N��@���SZ�G}���߾}�Vh<d�[M�]���&�g��l�ڮ]�4W�?��w����A&���sd�	�h<Br�dt����v ��wE�Z_�J�d�P��K�U󩛿���0��[�n�xf�|��	R�����.`���UmY������͛7_3�cy�ؗ�[͹Ď�T.�u:܂�x��^"Ye���	M��A�	�w8���5�a᤼s�k�V�X~�����qH�u'}��<������B4��@ B���+���+���W�%�ǀZ�d�ƠwO���ΈF"4���#p�67z�\�����*]�q)��ɈE]I��o9[�g��͝�L �7� 7-���(RtJ�;	N�k�y{k���(Z� %]w{�6��R�9�Nh"�f�D��	-Ѣn��k�{M���S���X��"?;]�����:ۨ/Hۖ
b��V���*��� .��˗[�~�`�ݸ0z��d|�"�Z�:��4i8_P;���>�xtѹ�Q��W&��b�ŗq�v(�#��!|E Tc�u&�� z��`c�)Y�htk�u��c��ܹ�	����XC�S�	M���\�$�|�Lh���������td�b�?܁!u��,L_ș���5�'��ްe]����\�&�$���@下�C4�g&ךr�s�W����, o��?�X�~x�\��0%�N<	�
7dbJ4�ănF#����"�3sv�����g	
�;��,k̾i���lA��� 봜˵o�3�[�,���Lj3����Ř��o��F
��7t*Z+�ṪQpѿ��|�L,�b#kވ@�-�7�=%^)o���v�e�s����>����h��Ѣ���E��S��k��=I)��9Lxά��EW�YF�4�I����S����p�S���ǲ�s*�p�f�	@��ܗ��BɃ���I�P	�O�#�qIH5��%���j�䘦3��.T�8p@�U�!��|f ��hq���,Q�.]�O�N_o;k+&� ��߿�T������7��<��$��Pq	F'^ꂚ�r�$��n(��i���ۥ}�U�|��ꋂzS�J��z�t�z��C��P��D �:���)P�x�Y^�dELNLc:�&U�$����1����R�%����y��'?����?�X~����g!�p��L�r�U&I@i�N  ��IDAT�����o��$�Ic����#��Jo�j�2#��� �^}�U\�Ȣl`�&��"
FV%b���S�
����]�B���C�N�,L�0��]4*����4-�J���p�Ӻ��4�ޏX����ԏR�y =�&�g@�~��4us�p=����$QH�DM)��s�d=KxKB݌���$ɩ����?"{K}��y�5����=#�j7�< h`�W��o�شE%<�$ �6%��.�EN^�k*c�X+�Dt���[����h�X"0�����v3!1��z�'�� ��
e�<}��#Ɗ���N>�{�����(-���2�I<��� �X�i��i��c��[�F�B/�r�f;���<T���:�L�>�!�f`k#ٮ:�0`K�*�`f X�چ�����
lQ\Ok>�2�ؤ��-XL_�Ke^�!��dn�l +�EG�ƚ2ueo�B䗨]1�%���ę	<&܁�ے�#*91�0.n=t�L�R���5�nj}�\��;���[��
��ª�5.�ŦEw���6�2��Q��sI&m[�M۝���B�	�N���l����P�� ��
r��	;��`c�i����@U#Xr`S�D�'ה���#�bYM#4���0��㊀��
����+^.���a�[-��9��j* �
s�Ҥ�ES0HWDX�$=1[)��r�� jC�,�*��+u~����w�k��^��П�~�l���7����%ʑ;�H��Ǚ��d}~���t��ARP�����
�����Hd�q�7}H�>�{/���M�#J�ȉE�!���<F���H�8�>�U�σ��,ţr�@������p�z�s"'�e����0f�Iq\Vt1�^d(��mI��Ŏ%��,�S��ʏ��_�K�E������Y��Pl��>6�lx�w���G>B���d�궺��Ѩ,���\�Zt�M OS�Ug�Q!��Y�# ���d����_�86:zQo��J F=�߷��w�|��o�U�k���ţG� &4��e��.g��������{o�ȁ��e.x���={,#���2�Mr�5<���?���޽[/B�4/�����>��p���x�=�m#�X�J8�
�Μ>m�7���׿�я~bޤ�9n���R4�_����^�u,�c��M���Y�z�SO=�?}����)�"%�[o�mӦM؇�5ږ�]�O�Ҩ�y����wϝ?'y�-�ߑT�|Z-Ԣ�a��*i�3���NL�X�_���������f}��T
I>݊�*�����s'2$���?8�9wz)Ɂ�+�b8��m��v���s�ϐ�o����d�jib�O���5HIQ����HR堷 ���f�2!謀�,v����M�9��0���1�#�~���x�Pv<g��f�Į@[��p~4J����V�E�.���O!�}�t|�Ҝ��So��+�V�\7g��	�+8�d&c!h^������Z���c(�{$�z˕�zH��ɩ�g�V�g���)�����A�1C<����di�M� ֓jfg���W�hVurq9S��^#���J�ݛ�	�8�<L8׃�ځ���~tt;P�_�K'�F�,g��5���oN�;Ơ�K�i�yP3M����f��b���,:���.�����ٙ��y��0������!�2���M��=���@Fܐ�E�C٠:���r���^I����>:iZ-I�.-�׋$TAHt�r�(� 0��;CG����_��5���Kנ���a���QE���/F�Q~�,K���q��gR�2U��Wt�� �Jy���ƍi��hv��*PR�NB��^�4�,�b���l������D��g�#�8��V��ȑ#`D- ���5-d���1�9�AЌI����yg�I��cT5jq!Lj��8<LWR6��WWB�	eҐ]Qe&I��2�[�G��`��/�E���6����1�
Jޒ�$!���}F7�!��sl>H.��BƫGP��E�p1����0����bW�(jz?V��(��BS36?��?�E�h��s�<�Ľ�,���QT{��*�CrǤ~�Ӓq�F:k��)@���(d�k�W�jr��ܱ���k���	v�H��G�տ���z�٧����sڇ�(�����D�XD��w��;v�|�СC�Ր9�:�Сx���?��k�zǶW���?�=W�Z�D$&m��r����Oo߾�����=z�H�s��f�2�TC3���|E�	��%#�N��'_��8`2�р�c�����h�4��o6vV� }�{�ۻgO�['��گ��o��<xT;\{OPت��9�J�e�}�I��aW�l�8�Z���n�]mY��S	�9@t,����e�8}}[�l!�V��J��D�=orH۲��1�4���K@Pʗ�~�r�|���O�&��}W�y���+�C���(l�f$$��R��Yw��0A�^Ad� �IKū�5����ç�C� w�R��s�=����o}bȜS5�2D�򓄲 �fI$P�1�
��}�~x4�$���bD�q b�O%U����f}��c^Qh�<��-��ĽeCr�.-(.�4��WNp~뻟��g��>9�D�6W�.�ǟjҲl���\b�Z���� �SpЍ�YL�4�҅
�K��b4��rYGڳ-��配>��ێ=x��K�a�iǸl�~r���[p��S)>rJ��b�d.����(�V(�u,�����Ȅ�x1��!�`A�� ͜W�&�(�K�+kc�wϤ���H��j'"đw���.��b�ֽ55����G��f��������Ip�at��n�����zgC�W�`Hꚏ�v4%!g2��ۡY��FT�X-�$M�
 �6-%|x�RO��<���p��0�;iH^Ƃ���*^�}��ު7��pM�4^Dbҹ�N����8J��>����M	IӋk���>qD�߿_J�DK41"^�D�;?:693M��*�Nn�.�2q���K�,��a�>+x�>K�Sg��Z�_4G�u���d�K���(��=J�X�ę�Ⱥ3F�xL3��H��1�!ACz,$2M�5���Ljo��ό{�W�V��K}�v���ԳR�]MK�6�K��<� 2z]F=#V/ٖzЦM��+���mԌ�/����Ѱ7lؠ��|Y�B�W��I�21�L��[R��B�t�c��=d�8y����gT/j� g�CiP�gm!>r����6�&pŊ���<�.���1���P� �,>l9��������������ҟ�}�]}Q��Ebs�SO=��O���/m*�MU��]8�^X��Ś�RM� �F�j�����?�����.�z�r��vц���o�V_��}�۷�0����g?��7��.����^[3�J�EG��}�c/���믿���Ϟ=��i$z��~��_��W7o�\�Y�oM��>��O����+l�����"RL-l�lH�D E_�P�P�jP�����'�mN��HH<^�i�p��FL?6�N�[C�O������l{�	A+/��J��$pc3���(����в���e�_8���N�9��O�5cfrJ���b�m��E��+GN��&�n�7\�.LON�I�u��$9-p��-#�l�pjr�Xeŋ/�����D��@D�?�&DeD�*)��P1��������sc�X���(����}}C��W����B��i3�uJE�=��n��:�C�!��M�$�K(�N(u�e���㳿�/}�R${*(�|����ԩ;�#�It�y�	Z���6���#D �J���Wç�	�ks_y&S'+;�h��]��D�漢+~�b�9�f�I���:���UV؜,@<N �kAp_c��q$�2.zy�_�>�r�!N�(�!ݙr\�F�B���$�/P:q�'�� ��c��b/@aH�v�t��X�#����?Qlt��cI$��[��E/���M�����&����=C�41y��I>�ݲ����{�EL��t؋�V���|�sG�M��
R+˨.��"���B��sw)g�n�xp	e}�b ���l��_?�i<sB��v~7n��� X�4Ӎp���AH�yJp�<*t1�)�yo���u�ɓ'AZ�����;Ӈ[H�M�^ǃA=�R��IF�)4�c��s��DN�ꕫ�Т¿�ۿA3�c� (~��Q�j���$��I����X׀�� ���5xj���(D�鴑�Rf(u���G*��Қ '-�'�Q�	��ժ����C����nZ&)��ЍΆ����¬�L/�Q�ߵ"|�yK�|P���$N�~���W�a(t���:ߺu��	��4Ia7�.��>>񠰞���_͞�Q_���z���I��Bӥ�D k-���+Vk�����?��/�AG��G>��gx��x�	���&����'>��&�s��R��rf�[o��{��􎂆z�0�}���Ε	�D�M���/Y'����G����%�ī����o����7�7-�8zI�c�b���s�Ʃ��#��x�����4~��M�Ʃ�k·l����~���~�7t���0�t�P��$��P���p�<xPo��m۶M甽���sϝzGM��O�����'O�ȣ�|@O�μ��[����1J��ح���*@��p����h�bv��eM�]����s4��&�"rj�̙���	��1	@vnZ���;6ݩ����YZ�fM�h*�-�!Ū�f�S:'y��eK�K��#������T�.�Ǌ7hџ �%���5�Q@�����i�(,���0�i5;DbH���P��a'"�$
�
l�T����	IK�5}��x�yV�3��.�f��(��k�%��#:j�ϴ�ٙ�wa�/��>�Vg��!�^:�/�1��u��c��]#�b�T!m��M��6�-�j�Q�ӈ5���/^}�т�/
>&��V]t!�:��.�^v��#��]�a�拔aiOFn����/���#@��<W��5y�pP6�nc���a��2�����]�ݿ�����e�CSGb���<oay-���GKA�,�K}ڶ%|���΢�E���'��
A��2�^嵓�K�s�L����5�Ӎ����X�\���wrRg�F��Ȱ%����y����kT>#E��|m&��m߷&'�(�]DM�'i��Yc]԰%�NNtIe�e#+�f���i{����r��fc��TR[p�{*F����?�8\�g롵���ڐ+�2\b��%�
�g�����Z����)��������K)	|?z5�E�<X��qðK�\���%���+���߷D����I���[�����_�$T��9�& ��I����b^=��lA2k�pfzN�[(=f�n꿴��s3�7�[+���عsg�n�?��S�+4#
|�7H �����$�v.]��r�M���ţ��u@��Q��N�H��^��3
;0�ug3��T�n�&]F_V#*
9u��I�.�1�?K����W���3i��Yy)Gǅ�9�m��Jْ���.�?7[��Ѻ3�6� �D�F�Vx�
�e;�;6O:�<b��d����]"�ƛ�+ñc�Щ�t`�y��p�X���2>���� C���%|��-���Μy`˖[n���������eP��^� 3:u���g�ޡ�Ę&Q{�ZSH7反}��һz��+W=~\@j��z�ro���SV�R�9qT���w:rD����1� 0�=��3?��3��ӧϮX�J�[f��9��uso�V�Q�/��̮\�J�|���Z��n�M߅XDb�ҥ�ރa�1w��Ȳ���I��F���}Ng�Vm�͛�z�_h�i��w�����5>s�=�t	��Hm�<-�/�����Ѱl =0}V�ϓ0���]ᘌ�,�2*j�k�Ϟ����[��>|�H�a�v�����=7�[����+?ћ����
��g��B[Bg����w�Ǣ�jd�p_�ej�ͽ��$Xr��{�#efs��B1o�v�U�͗{*k֭I�����B]��/#��� �����o�Vѳ���bijvN2�T��j���<~�豃G5*�yۖ���G�;����`tO����/���5f� �(� ���V�u���m��z��N9c6��B����Q~��jYa"�/G����O����;��x��fL7�t���m���i�۬�;�xYb&~n,��{zzM�fR��z���rͶ&�1D>_�\1c�+T����BG(�#�5!��Œ��͛�U��Ss�d;������ނ�5}�+���z�ҥ��f�*��7�$#K���%i�+�f�z{����h�v�:7�偭��VCk�ڶ����J�	�'-��$i{�:3�'��!�Z0�] +��8p�7��A���X�w� ]�Ew��iIHxE��_G���8!��'�=O��d�7<�@�2I�fS�`�Z]д��Ɛ:�����a��Zc��16JL�L�5ѱʖ Qe='� �\B$�~����8��^���Ysyo7���F�[�C�
��4ҖJ��.
�l3����V39�p5�N&�v����lg�!�p-E����4[L���9t'&>\\��;2�y����	��lt��)5��+Wƹ�S��Y�',.A�YS0?0xMu�d��|^II�g�-�>���D�uH��C+�0�/8Q1b�^)���t7��n������.�P#��6f8�����K㢶��Eh�"�yy���@�k;= ���B�2'xk����[��HU!P�%��Bk�47/UW|?���YRq�W�y���#T�	X��z:��#�N��� _�B���&A����ċ8 ��w��������+<x%�A$����8#_A�F-��'h{�7����}����Ϙ)q�����4{%�p��a�����{���(�)ѱ!K��ZP}P�`M)4P�<x&}�'�NPI�HZ���]8�5}i'�K�H��W�����O���w�;�̻��=5�A�r��9�3ރ�yGF�ZP��=��O�|�Mmx�%o*J��^ةz�5k���Ǐ���N��/�R�e'N�&uA��,���� �u=YGZ|���c�=�����<�۾w� ':��o�>'V��,�k�O�������n�k��G}T���I4��N.@͕��*`�ۀmP�Y�j�ԊC���k�W
ʴ�z��SO=E*�Hf�V� 8�Z<����g?�Y�ѧ�q?C~��`)�o?.#��f+�2�%�3]�u�I!�4�Tz���3?]�0�
�ɾB��ڕ,zpi�=�O�z��[�{�ܿ�Il{o�0B�%F�'E��@nki��%��_w��!�ѿ4�ןV�^u��1���s���y{׮�^j��EȘ�2[�b5!��P1M-��-��4]��s�hSF�i�0�	�TB�H<��`�TD�uS6����|P�qp�n�t��MӳT��)p2�|�px<�kĠ�}��q��'>�	iC6g��̣ݖ-���*�N�)�r���2����o��M���X{0ΐ	s��e�!5��+�:�&�wG�Eb�j^[�zN'��bD��ďzFw�<�Upg,5K��0�`!axHi�1��HÏXJ�2��⽲�ǧ�y":4��!��,���%���u�}��1��󆧙no��{2�5a�⩵?e�Hr2�d��M�Vz����L6�/t�ҡl.O��Ь-���������n�&ֆ����V�h�L2��R��u�yܧ�@N��h/�8����S�D�^�'�����W��k�ۺż!&����K�_̅D�h��U��~��q<�T�!�����߳��/Ғ�`���x}I�M��&�������w2��x�l��&�1�I�a�_��&�~���F9 �:\�9��B�Y�� K,��@dc����+����^
Q0E+��؀ʏ�[��u���%&t�[n�����`b��0� �ω2����(IC�u�X��C�;c�a�ZO���qxw8E�N�";a���wn���$ؚx�*�E�~��V���������J s�<��s)0ieDLtw��CtK�.�4X���p��S�z�/*�EU�k�Q9$2r� �R����߶m�K/���_w޻w/^�J�����2��}�1P*j�wq��%����dǎ����eȇ�y��U-�",~����^���,uv�rYF�[Q�K*!��+X��C|��9�@+ ����) ��v�m�ë��J>���ظq����5��۷�\�bϞ�d��԰&�B��	���f�����kHZ#�=�.�Y}Es+�Ly��z�ҁju9�LԒ��t�D�	�	~�{�Ѐ[�K�����4<a_�� ],4��ӿA�T�Dj�i`[�n�V�Z�V*���AARBc����&'4g��a��bF/���ٳgbzJ�/C5���'_����ؒA:U�Y��E��\�}�7�S9&�T�pÒ��f�Ո�k���h�skk+<A�>��4n�0�h� C�3j5��3�b�Zꘟ2�j�v9�<5�=3�-��g�K3��BylE��6�!�/s��<��ti�Ɉ"��.����H%��L�v�]l���ߕ��������eg$1��j �=�&3lz�;����\�T�2�˛+YΙ5c���6C�M\ki�� =�<G�4iyW��T\n�!�_-��3NS��c@���vh�@um#4S���֩����Hv�k�., ��W�$E�1��� ⇋��l�O@c�@)�D�I6�;:�����u-�_��֪�[�8(�YD� ڵ��O۳��i㤕u���%u����u�d�Ȧ�����&A��	q8xt ,�PsP��9��r�Q��ƅ㳜�%� �ӳ�'d������
Af:en$@�419�=}�皁�SC�Y�#�K�0��L���n�R��Qժe�K�J��ʨ����S�a�`?��ga13��G�~��f3]�L�>���'�S�67��=*ߺ/]&Y��'���J����"`=���	A�V0p �������@��R���N:����%�����^����k���}�x!�h$�O�5�\�{4�.%�Iw�2��M��͛���$�j���[$����1�O(G�Ꝥ�9�L��J-y��
�����E� ����ʜhJ)�����]�mCh�����O��&��q���v$�2�����{���s�i�
��S�44���_�ҥ�"�
E�����do������z��󺹃�
���.�	��Y���`�a�5!�֭դi��}��"$>��BVo�I�M�g7R���dx�����=�h��C��s:��?��O�	�BpF�9�ÜYЏv��D��Wc�|+�/�����:���_����}��Ma,�=ܖ�AƴZ���K�k�������v�M�σ�O���ꯂe��w����C��&f�&�|G�	��HU$����ĉMg�,�-�Ln	�L�7��h���-@��n9���=���C�,�,�Cih.L�V��O^!c�~��|Զn����Ͽ�� ��w��U�UC�''1��2��}���ڦL�hY<^-7'&�Pj&�ZY�w7���>i,dC��3����U�T��U���n\2̢�A����C�j��Mu���vl���?M��K���Ǥe=�_^�������tF��2%;��=�t�6�P2dj��o�I���[`YL��|����T��Rkv���hC�Z���e`���%>Z n��褆��k@��a���@RӒP���2��!���.���@�ǇU3GT��\���f���li�UM�x3�K��������!��J^�7��E//'(��F���>kf�Z/�.�e'�)�c ��3�Z���w%}�X�#��q�Yv��ҋ�h�ĢE"��2L#�ٸy��x�aА1$!tX�[�5[�W�o\�~�&7g���%�v���HT���e+[�Ǟ��C��F_^�h�LVz���;[!|fĂ	��X/ #��$/Ñ,u&�h/����n�4D�P��Ǚ u��x��+���������kV����܀S3�A�`��5���iף����5�k�i�7N&����l��!%�� �G�ԓ����B �9Z�~2| ��Ԏ`!��'��'�R�0��sZ�K��h#�C�ih� ��1�ˇ'?��%R�0��q�˴��[CbK�k9vs�4TI�bx�t� �f���_�[�t�$�)�j|NRf����SE��۷o�#H�JQzz��ݒ_�?��MYb;�4�'�hEȲ҃�&x�'5=�'��a`&ZA�T�UHB�^��>�������ߺu+�oݙ����㳳���e��t�s�=��m۶Z��{�k������{{�d}�sf�߿_3�~�z`1@6�M���/��6l���E[-�g����~X#��७�u��n�mϞ=zM;Kü�=G���7o;����.��1��E�E�>�S�(�"�GMK��k��)o����ٳ������^�	�饀错S�
4�{k��;���5��"�^ҏ�D�W�"����50����H��:i��>�1m�%C��Pȥ�k�)L�D�GSW��y�G�LN���`emvΚ��+�Eݓ�mÍ:�DǣW����uj
)�'�,=�ΰ3ag({5 H.6`�����.O��j?���j���կ�>uj�w΅.j$'q�v+ƿ L1{	�j��[r�8���MT�9����u.�UJ�i ���l��s��&�R9$�CK��8ɋ~Lv%:��:���2OJɹW"�� 4= l�b�����֧8�B(߻w�����g�y��uQ�G7��oO��l��k*C���b�ݱ%Z!4�MB�ZH7������Sw�|T9�F�[-:�c�+�y��Ϻu �����*4�G�e���]ʺ��y�a�B!�zUr�H�j���pP�i��!�����i��<��8�΢��1��OC��d;%�n�ڋ4tR�Qʊ����l&I�iF��C��k�$�.���o���}�����+Wq�x�j����2 ��NCE>�x�*m�I�P��t���J=�����Pg�l��Z��.	 h,H6"E�<$*FIt��`��C�m�L��ј�ds�Y8I[G�Ay�H|"x����_�x��;{	I`xV�y
��
[ֆBaV]�s��O]��
�Z��)\"[��{�4W@ѻ�B-�v��1�^�����eˮ�(^k�u[
e@m)�q����}��o�})�����g ̮�)�%���C�W ����3O�I(AV8���!�tu�TWj�`��W�I.G�Ť[�6��㤔^�ݍnx�7��;wZvEO��|=B7��9|����K<W�r�-����!����iO
F+ι..�L���W*j5~�"�{�A���;i���2��(i�]/�u�eC��%�r�E{��&j46m�m۶	�Qq�G���;�6m�>�u��7����H�G�+�m�46]0[����w�-���&�H��9"Űz��D= 7�����uM,a���C�e-٨�Bu�+-=�:_�mH�ky�f�\(�K䌋B\z�A�'�|�B���M���a����
��醄��Θ���}N�.\� s����S��q�d�4��9����kF?��E�9���ݴ�d���M��!P�ԙ��hII�����>O�YF��} �� LU���-C�SC��h��G��|�2���/�����,�_���[�b���qJ��P~a����G��O�|�u�-��LG{���/ڢ�J�s�Cm#"h��ӽ��ts���"�� 4�����!��#��;���������ߐsF�� n�)��i.*�\�����8�ȴ_��!��,�k�2���-9D`�@�_�>T��� r��\��rY���g�w��1��O�Eɘ�fU�w��Gup�{̭5ۥI�W�,��|dv�N7����NNYԫ� �r��W&^�s�H�'آ��� �[͗�W
<p��KF�9Cl�T���=��A �M�]g\�PL<��.��|��g�{�?[�	#�1i�a�A����@m���X�'@���X)�~ao�Cɰ��2s�k�~Z�P����f����]�뺷��� �V!��8L�k�]|��YAg��b�\*ۮVr�b&��L�N����9*tMG�|�&�����B��[��Q*v7ktb粅j����Y���̲Yd���Dh�:<�ErEcӐP �˒4;�S�.�F{>Y�i�,8�$�H501!^ b��l2}���D�%ΤS/���E�oP<TU$����|�x�'� ��@^6(��=Tk[X��H���5�0N�������e}3t���eQ��%�O #@�P�����鶙��?�^GҐ�г����T,8@#����V/R��K�G;3������vg<�,��rR70��p�� QW?3=Wȗ�kV�059����$�_�ފ�e��,���Pkw�D�xe���Dp�#��K���u��B�{��?ϟE�Wn0�#� ��e��-���D�c�/��&���M7ݤ�׃4�$��bN+%Eo-
R׌1�9�AmN�i+h��������ߵk��?��F�-&u�(-��B*KtB��L�QWx�l6W�X��9����.N�����믟�reͺ��fp���8v���|��Ϗ�;wa����*��1�cu�w6Ն,�S��\�;]4�B�6l�m��4!�V	��GG�Έ!@�?d�t�Z�ά��mxw,�ƴ������G>���R_�75uDU�Z����%Ŷ}�v�i::�E��`���
�f�lx����\Oφ*�f(���ID>�6�v&����vz#�U��Y�!�l����f�u�W_}Ub
s\"�k_��6�&shx)���z}	U"E難��,g1_��&���l@��
��5M_�i����+?������%�4uT�j��K�Vy��t�c�/�:��+��pE�=Fbb�ePC�0Q�?z�����������+ɬX��;�i	�����@c�	-���C�B��u�H�F���s��(_BIc�������䉈9�Q��Ѱm�L��i���^�F&����S��bT��
�{��O�������j팻*_j��I�]�|%���,�o��7�U��
��ѹ��!U�8Yuj��V=_�Ip0�����Ej�$p[�Lh�V�cm'����$����/0�����J+F�-��S�h�	ٸ�����4��ֈn�NH�F_��v�7�$�'F9x��o�$�lhE�8m�3���8ёY�
��&!�-n��oꎲ���Y� �Ś3Z������j�J�~7��*E�~j|Z6�K-��ʵh_��p
�~z-k����W&	ٰ/!��1g��[R�:�Rrd�X��X�[�8��ܴe���x > f�x	�ڻ�a�
���J�7�M	Q;_�h ZMOO���S���0P�3�Ɔ�r��%�B�(|o ���	8F�Va&Ia�s�5<|��zk&>t�⨖B�[&&�z�+�Db��l$-�:��\�}I��2-!)Q]��H�3!hb��P���6�_�$�"���K�8�D<��!�����J�ar����_Өw�b�`.Xf58~bƏ��yF��7=����'�j�@r�Tڱ����F4(|��D�m������W�w!���Ɣv\���n��bcd��^"tu��w77J��j�p@��Vƫ*}I�1=�|���/�EY�ʙ3��bqI��{4 !!�@$��u}W�׷4	�i�[�
!�hc��ѴZ�=����CB��v�;���G�g߾}�F'BXmǎ�.+������>���^{M#)��͚�,c�9�ll�'N�2ݙ�-�&���Lۡ��H��v�-^(
J�N˼84|��2Kؐ���qB$�!�&���1�4�@Rs����IHQг4N�D�M7j:�>�Qj�#�x�钠�������z'�V���w������������>cؤp�؁˖U�7�I�h��9�N�!o����u�͛�;u�����y��V�LH�����ѳ2�(ՆD_r�H3"EL����f��#Ѻ�a%����/��"{��[��F�9I�O��O46�c�ykb�=,^�]BD4H1��#��E����Eln�0�zz��������a�@�bX����N�:�%�j�((�$���,צ:v��}�7�ٟ��K�Uˡ�t�-�h��8��;�O�O�w).��H��A�~��շ�ڽ$ؠ�4�����5*d��#>F�\Ż�u��HS�R��B�+\��xP�-�q(����0��L�4I��-9�-ۀ�P�wI������"R�v�BKC�(�$�	��� ;$F6[�[��N2m���-u'H��H��&����na�r%�xae�����w�m:L\�P����.��Qo�V���f�I2���h���\�JOͩ��-]���zlbҵڠ���I��o�+ט���nU�zks��$���!�?�
�ӑz��6��wG�{���%�i�8�֮[ח�:�y��;ֈ�+e4tmQ�?�����3��.�bWN��)���{Z�w��ԽU��6��0�k��C}̈́�,�w�����t:��M���㧽����,�3�㩿��� J��|��yw���";::�;cq����	l�%%�$)�ؒ<�;e�,l��{ｗ���h��+z��3�/�_���_�z�匸8<B�^�z�gC�Yb�o�F<��T�N])�
\�<@�j5��J� ��"���q<7�������ZoD�5��ĳx����E'�jJ)j0�?A����[�&Ӻ�r��٪W��u:7l�M#�{e�6�r]��P�I�8G4����C��Rj8�I� ����ģ�-@:�e�N�v44,0`Ě�c�<�����#�fl4��=���O?���3��kڱ�sxi��a���,�pX��+ԽS*tޒΘ:�7aL�E2����6�<���әŵ��n��FzWc�DqZ�z�!=�#�U,�����(�Ɏ�Ck��ڢ�-�~���^�l��˗ud��������m��%K���={��O������ן<��ۼ��>8�gg���4'�yoo�>�E�5%_~�֭��޺뮻0Q�D��z�@��	�zMJ��7bw�=E(Ԏ'��1��_p�R�,�܋�(w0�M�Зϝ<}J�����?�߫�KG����=�%کC}�G����V��}�{��d��	�1V����S�wJ#}�I���}�f`Ӧ;f�ǭD`bz����{���7�xCK�p��7mԊ�n@��gMh5ёX�ԏ/_�����.�?��1r��nh���6m��7��կ~U��F7x�.2���(���ϹZ��j#��I-1c�����$�I����d�'�v1_�NC�ZH�N�m�X�L�LX �(�	�3j�E��������y�f�  G2!�k��fZ�ϟ?sÍ���_7ݼ�O;��[oeW�K=XnP����i��r�MG����uPBZ~H�C�k+�����@[��zM���u8���<�x�8z�I_�ip8Yn����N��<�	$�	B��v��Ck�9H�վܰǛ�j��@8L��{�']G g����l.�!jT�����1g�m$py�!�E?�<~Ǒ���<��f����슒�K������p#X�A�M����B!�G�%��0>�;,d��r֘5�"G��Mz�A� ��ڰ��$�đ��-5�X�ғB{�R�� ���~�{���%$��z:���}�W�&�7cy`�#�Q<�`��X��%O@�E�)�̺��
��%\�~
��������P�G�`-��@ၥ���3c%d�/��y���3��".���8U��%���.��U���;�7�?�(kW�B���u+�������. �f�<$��;^�����?2�t��w�M�����z�ԌF�w*�m�Q��~��Z_}x���ՇE���)"U��n����z������P3���n���h"��ڜ�R��Ki�h=������4* pJ��"�,�DF�G�e=t/���j�rN2��x�����j*4�d���
a2��$^�]D0�:xg�j x����� �%���\7��~��9r��_��_��L��}���� w�
�5���u�j�4�i.ܣ�A��VV�M�'�c����_h�<Nz�,���Z*ȥ� �� �ff��"oU�L�u��^{mӦMR�z"�?H�����J�V���GS�qj't��*lg���
�̆��7�|S3{"���2y����\��<s��,ݣ�Ut���u�mr�(�`��ڵ�01��*i��B�'z��7ꂝ;w��x�S��Z��ѩ'i��UH��#��}��	��ֲjɾ��������>��_��WFG/�[��{��yg[�Gkb53d֒-���}4?����^�Fɔ�Ûu'P�^o�F&Pv�,[:L�3��:�j�����K�4���5��MN.\0y�/��t����z������~������E=��GO�kg\&�-FƉ�H�?q�Lh��/3�j�5jx+��jW���F��3g��@��p�A,��l�ѹ|��+9y~��i�d���R��l��̨��/}I�S7��
�= &�a`����l!��iM���qR���d�$ͮ��h�r%Me��^8��n��"�,�Et+��-e︊�Z�#�km0��^�]}N]K�2R��y���%x���6eu�r�́z�K]��.U
rl��
�1�Ȣƽ�K���+�A�7|t3�@eC/�V(k��$M�PIV��2ZV`l�[ׯ����,(��o��ʦ��Z�=]�
�a�sƏ��tM��i�W��lNщ��eSsK
f-��8�Ѷː.@�b�$6��uщ�����!�>4�'�,�nIׁ�-���kW[����d-4&����U�bm+d��8q"mw�WI��y7Je��W����y�<�B�)�W�+��b{�d���q�0H<��aL��PG"I�����~�NE�!��L"�"�I���G�P/Fւ�׆��5z�;w�L[��sm�4���\�@�Ж�%f}�Z�YoL�uD��m���b֐%�Τ���guJ����f<ǘuxtY�:�(Ү���[�B�T�)������=q�sw�i����ޑW^�5"d�[�{�����,lw\>x7	w��=�Œ���9�d�P��p�o*8I(��c�]Z�8�	�8Wݓ�QD��WRp(���,�}N>���0%��tHD�%�����KB�HO��^}�U�ڗ��z�'�dD�ｧ�{3�[OM�+aT6�B9�P��K�M�P�5�G��[��T��I՞?V�_���Y:� W�����5�m۶�R�O?��n������?��VD�&���}O/H���fphH��cU�6n�e��s�E^;\�vq|\� ��S�yz�����K�i��Wz��η�g�x"���R�@��_"��d���b����N�t,���$hӎ����Cb�������0�tU-����<+H�EH�^A�=p���,�����ӄl޼��ױ�x�	�Q�;h��E��Z��z�Pҭ�j�:��N`��n4�ظ�䊅4���0``P��g�ܤ�\ L�'�R�	��@���j�t��G��s���E�������?��i��}�~��?��?��?�C2\��A���]�9'`&ۡs�h��@O
�S�i�O�Q܋a�e���W�J�N�ղZ��mH=�1ϝ9��2� ��,�R�XbI���\�,[j=����3�
��׿�u�0�9�֧N֔�*:�noO�kɡRE���qs�d�T%qB��æ�׬��[7۰5Ռix7n� �_���<c%�m�+Iv~nl�B�g��TH�� �K�S��:4�j���Ʃ�"�8����R 4qa���\»F������8����r�*������v8����b�'���c<��`���D�-}�Q>��+�Q-|�u�ɢ���lFGH,c����7=C8�Z�ɵ'[�Z;XS3i.Ù�xq�{�[�1�o1Y?>>�U�x_h9��fC	R����T�ndBg�*9G�w�{��E;{��3����5ICi�b.���M�n,�z�o������[Ed��t�O�	�	���n���4$*��C&�cFsC,�3�����O^-�W�[e���Ȏ��({;����=��3�����v�x�q�l&;��H��Du/%T���{�"ݶ�!UB�(�h+�B��@)RXJI�؎ǎ��$��2�ǳ�}�������!m����t|�=��{˳~��[��C�������W� Z�"�Q���k��&�V��kH��� b�I��bΞ����� &�Y���3���j[<�#��Gk�%��<L8�A8Q���{��f��e$IO�'&0�҇?�aN`қ��*apC`�5�]���}@~ԅ���+V��Ux,1�v�Vt� jf���_���-�;+1�����̗���h�����h� �11)C��2}��5B�rE3)����hb�& H�,.`��ޤ�u+�W�'�A#�#�M�[�x�o}�[� S��_����K�p�=�h��!�4{���'��t�\L�
�Ę�n�u��i93��J�b� pyHԜ���|3�tG��;��]9�]ԧ��2q�Р�)O��'J��S�J8f���U�۷o�ץ�5$�gz���l>�h2�1���3�<�oi�� rĘw6 �I|ie b�r�V��5��ҥ��fL[���6�_�	,���O
V��r ��yw
��F*SWʚ�Ɯ��{�m� Q=���/�=��r���@�;���7��4�q�ML,[��w�w�'=W���QKSGhӾz9`FT/A.�l_Jtu�. \T������C�e�q.0�5�2��r�#���#��5�[o���cK�B���B«a�I�k�¨"�v߾}>���^;�K�|�3��v�׾��C���*�4����%�+p'1�T�Ң(���"�݋�h#�B�|;���
0�oG��Z1�--Ќ�t;�J�~�sJm͍+nJ�JFɒ���>�����b����.���t �h���3�*���$,kֈ�e��m�~0��.�.xf��{�1D���^[���R�b�*�*�C�{��@PmBk�Τ�=P+`a�eli[5$>G��Mr�&��dFv"�1�h�f�QS[M��E2�\{9�f�He�C(��Ią(5�8�E�'08������zIy1e�H63��wD���a\�Z���"��w>׳���Q+�9�A��h씖��]=KW,7�sVOd��F�\*�<
b�߻j����:B�=݃�C�Z����2m��%��B4hð�	�ږ�5W\�zmj��{��N�U�%��F<]kw:�ջ��N���T���\#P�� �$!�ߥ	4 	mSH<X��u=n��PX�(��[��,����
�x�g�I4�uؒ=�WD�7-���g�.].�~��qJ4*mD�ۺ��{Y>Qr37������{ ��Q%�	���
�]�kڨ��+43̿furr��2z��D��k�-pέ
ġ֑�h��h�p��Á���t��]I%�ȁ~K�LLLbk;|��[r����h�d/�r ����C��\-�M��	F�y���zM*K�$���!ɕ�k~��'V�\MY������.)4JH��&�?L��u�c3΄��~A�d��>���l�@�1w`�عs'`,R!���O���[O?�4�����5�z��~��[�n%I�����Á��
�N7
�3xڱ\�(T�Z�$�Ǥ۴im�-O�:q�w�څ���� 5�l��G鯲��\��4��M4�Q�	�g>�}�����o��v@���(l)��q�wv��L�v�]w�Κ�GV���fO3��h�i�!SI7��e7l���믓D����8�P�:��!z���Ѻ��C�����r�cp���i�\w��w�4Qē��ƀ����f;u�m]������|�ߔ�MA�v�����?��?��?H,D� �/� U��$+J�n�(xY ��֭טϾm5�K�/�߬��܅������o������'�"(xc�"g� ��=����_��/7�@�YW {@^v:b �Z�(}E/���V�"�>�W��:����/~Q��'�'�.^�~�ZC����F���P��KHJ����gs&Ѓ��̳�杖���(�fLo*@Wk>��M��U>���<&W����vF��n�52p�FN7�,q����?����/�@��zci9qb����<�y��GL��y��j�Ij��T�t�{���d:���غw��LR������txg��W�j1`9��R�!���_@��Bc�@�	�*�8�ZN����%��I����%Fh�/b��J�'�cB!��ŐJ:GU�פ`":7�"n��3�Gq�ps�o#��g�AY�hb6݆�Y���l}jq�R
����l%����L
d<�;��Ycq��9��-��3��Wj
���l�{��П��g[��T#���p��b�Nۅ�j��J�<����bQ�\����Ѧ��������n��v@!g\hIߎ�&���p�K��1M��d=:��t�T��I蛀�^D�'�DhA<0y��$"� Sq�:�B��Ct�5Rl�q(o�*w�J^�ݚ@���fg�=f��s٬2n E����q%�꧱�aq�!��RԈ�1�qꕯ��ioĦ?I�Ip��Ff*bp�Iӎ�L|TÃ$ D��E��.fR���SO=�ρ"�	�a
�$I`�V� �d��� Te�Z<9����- B���-[�d����OSvr�[�-,̑gt�a�_������Pm{�.�)@b��� �QBD.��G�ٱc�^p	�R�V��(�ǚ�;�r�@0d����me� RI|�;��P{�1��f^W�����4R�@�������7�׺�ݽ�$�)-�M�z�����_�|{�:|�nAC���hdy� �/8��s��/t6�zW���4"���ڜ{̓���ի3�$K���i�L���R�Z��ee�a��߶m���,[�T��b� Q��Yt��2o�[08�%�E��T�c:��|��j����O@k���-[р�����4�z��'OR��1��g�������i͚�D֑��:H>�J}�		>O�FoM�z��$vSNȇ\�h�n�ݬ��Y7X-��h�R����"�%�~͚52�����<�>Ѵ��^ �8uF�G�
V�$��A.�S�&f����tL���/��曩t�1�{f���=35�k�cE��G�wx+9�h`:��uv��Y<b!����h�ٴXQ��f��p�	�p	oqҠ:#���k��8���?}�u����Hk�_}�U�E�6AU̆��]r{�f�����H#�Vu$܁�D	��ψ/p$9�C\	�%7_"���A0�7�R̠�������W��ZǢ�]�v(�u��T��ɉ}Ff�����	�U�I�h1Z�C$�fVH�50/�I��X~��-�̢���Y�i;�^�d#Y�*���d�2�BL�mٿ��lG�ڿG�D��o7+�V��h���*���<V�10S<�j�R3Կ�Q2W�����B��h�����@3i��[��i�L:���q\�d��uØ����̞�|Fd�٨ҶZ}�$����8��:�fgee����Bwp`���^��y��K�G[������"�ٓhWu�Д�4�#n��BK"�cX� <�Z��X���5c��� ��(��"�;]]=R�WqeS�;���j�id������s�>t �0\� ����c��6nܨ�8p NƩ��%�w뭷"G���3rٴ����?'E%MFÜ�s��W^yE�w�M7�;}��.x��5����3�^���a
A����EX���T˙3o�o4k ��Sã2~�Z�H5<�R �"�J���9��iPY�^�=�$[����J��~&m�  .���[2�\B����xl3
��b�Ľv�� ��߯��u8I
�ݾ}�d~I=��Ym9�K�kj��ɣ�>��O|B���424|��5����T���BP~ˎ��$ъV,[�����=ٰa=��2J,�4;�8�u�xnq���L�j���?�f���]��6 ����=��������_�R��������8�"�TDꗛn����޽{���l?��uOLX$F��Jg�	�H�K|�._���0R����F(���s����W�^.5DM[�<�VVGP��n����o�_"^�éO`�X��V�&=>�_.Wx�\.%�Q���/x�e��?��?�I��T��pl�G�G��"݄X8$R�:��t�(A�A-��鼬x��W��0�.��z�IO�YH��*�t��o�ASH�,����X��r:zQ0���j
�$���a�J5 y:,Ē�15~m��+�����cգ_�җ���oz��g�c�x�e�v�L����\@b����I���<�e�dRi�M�PX�bN-Q#�������e�ӎbZ(7�S�*��LgϜ��}��|�+_цoy�fR�K�\�����0�Kqdҩ�@�(�L� $���3	�%�FS1_+�&�3�O0����&3F���5>j��0����Z�(�2\8/�뜝��EERZ�?��%�~��>-�3F!ˇ�@�`a�]��/_J|��N0A�'���8��*[�(>J����f��|�T��!�on�[&��4�lU��x������ͣE��C�GK��Ƿ�l|Q�*�	C����&�A���Mŷr�@�zãt�J&@or�՞�L1}$%^u�ݭW�Ƌ�Rk�Ȑ�jKX�렎:Fxdp��Is�I��0Swv��2��r͐"�CиcK��$��� �C��(I��`25����i����ҋ�
��<&���(�Y���t%�C7߼�~D�����,�
�E���]rmbb\����$�fH���C�8�C%L�O�I�ɯ�] ~D��u�Y�$\@GE�"�Ř�J	V���QO���J�|!����%���Le)�p�f}A����vT }(�� ^����st*�6�rx_��=��-�==�I�[QQ/0��ݖ�W�� �&8��j������W�8C��g��ZR�tg*(5	j�]NS$��P�|+V���[R	-@�z퉻w�Gϥ�F��~X�o|C7џμ�v�79�}����䥗^y��4K�=p<��N}W��W���ۻw/�����R�/�����i�=Eb.��e�^���tI�]��K爥Y�z`@�B�ִk���qY:n�����nAv�^A��su�={(��M���*����{r�I[azܳ�>����? ��웑�!�����g?[�n���۵�6<���.�,�n/v�رCv��}����x���F�e�;��O�S]������O�O��k�qj��VaD��U��ґ6�cǎ1hq��
���St���Q=*1�������Im9��V=[d2��uَz�f����ܙ��[�=�������}�:�,�h�5�f�U�������e�[`�Mo��6i̚�vgD����E�)E�L�h���Qha	��K�W׌&w�狯!��i�>��Oj2��~�{����"Q�5�rK�8�66r�t�T�J��*NfM˪���,-[1j�@��y&�Ią|HP��5~2np'R��A'!��|�����d���~'�P����t��*c&���y*���AP@Ub6���.X�T�CZddHB:�_hv�`p�A��jظf��JCC���Q%��0Ԋ�"� ��s(xǂ`���)M���d�c�~��8��A������8�seT!���v�� �eb`� '͖ðN�ܮ���ǀ�{&�>?�t�Ix�'��	����kU����;13~i�ۮ�;r��8�n�r����Ȼ�7�F6��&ӄg+�d}an��#;4��V}=�N4��K�/�?{n��Mݝ=F%Ҫ.Y��F:���f�je�;4l�J���6�o�y�Q󅡡�&��n5�ٞ�����Z�657E:���t:[����Z�o��&I���*L^�tc��]�DH+YM��&�x��_ 8��3o9��m��Nǲh�Y?��4�e��c�Q�`m^++�YV�D���F���]j��^���$�T���gg,l`�(��7�I���׃pO����%�9ݼ%G(��S�6�H�fF�)W���R	Eޯ�!9�� ����q֮KT�D���z�|G��Yћ��XkR3548�u�6=E��0�i��|[Aӹs�=�aA,M�ԛ��ؾ�%�����B92�bZ�Љ�֬�>j%���g�b�j�v������)�8��)+��q�p�d�䤕�/]:,��4%ɢry^V��]o!m�[Y�fw�=�i���������T��>�r���]�z�J%�I"��'W��\�:4���e��l0	�ȡ�z�BGכ���Ӝ�-&ġ���^e�>[�Q�{�
�)�vD^��{���Ov���"h'�� ,�ze+��zC|����>��s����+���p�%�}-��.��ئ��4�R�F��?��(&���Ch�׮Nk_��{uU�!iz����N���J.O��j�Z�N%��D�͘�;킻"���,���D׈��c{{�<�K�ݘ�L͸�&�uK���!b���h����%�fmdģ�z�d ��&&.wzbK���g�dC=��0��@�
F:$�ie'2��=󋧭6Ы�l���;��Y��v���Y\���[|\\V��Q]?~�"�%L�ޚ�+��C}��������G>"���%�O�J3O����;�A���k�m�Yr���
V��r��*�Oǐ
�'-��:|�O��yi~A�'�L�tt�ՅJG�cۖ-G��QgOWWs͚뵂o�u��y��ʕڵ�K^K��V��X�|��{���M�@2�ڵ��aY�W�|�6Ɔ7"��s&i?�EI��3���<��}��w�u�����_�h��~�9&}_�p��򽀢�bmVo6��b��BT���6MڨUKu7�<��聖zia�]oszKOU�]c�I�	hRk*?��ZE�!kϓ�\�T���'����ٟe3Y�8��]]=^��-�Q����̌Q�n�;5�s��*E0SW�Xe^�d����e#�޳�{������\G_!�_�W'9#Q�a��l5�}���z������?,`r,Na��-�L�HGc]�"��P�V'Q�21)�D2w��5���?R#X5���l%\�H4���,j�M�� �Nٗ�.]Fa-Y2,U�X	�\/]/ǀ���!��ʋ���{�R�\n���\6�W��n]�`����"�9H��	�A��s�7�f�\�ؑZזk�әF�|$�&_����j*��kF�����$LV�O���c�I�ʈSq��L��FV�
�D\;�n�V+��~ԍ�Q����Ү:Y�!h�� �O�B��y���X#nK��o�,���]�%?�F��rk�.�싹ݿFb�]�W�s�@r�M�6��L�`�����mI"i)0pz��� �`1����v��|d�U\�$�@ܘ�+�ꩱv�>��U򂌟b� �o�#%=M�͉'`f���>hՄW�B������|�M�Kbz���:�m��t���FQݡ���'YZOA݂;$���Hn_�6�B �"CS��^Q�ԇ�W۝�^����.YTP�8�	����+�%�Պ��C6So$��T)�`�%�p�u��j�ҙ���m �'-Aف4�$��Wӳ��"����<�2=��kC���.�uZ�;^蹍������.)X���p�H�ux~���#�CT�@fQ�gy�[n�D�뮻����~�޽_ě^�[Iw�O� ��z#���Ӆ�Ν3X�Uk}�y�y<@�;K&"��WK�̭�� At�E�)�]���q�>��2F�h-"�,��ݗ�?wN�%D����KO�]�DO�����$Y�ú]����!�3�5���O@�S��S�����5r�Bu�u�8�¨P�B���xf���s�mz��[8)��TW�X��t�h�s��n��{�w׮]2��N��ԧ��G��b��+�`@��q�y��i2��W���ohf�`A"�åM(Y�g��m۶��O`7C# �]F���<q�6ώ�Ϝ9G�r��s�S%G(ՋX&��72�/ɞI/�ע�ŉ�����G}�[�������"Bu��.�����!����D)�q�2����Y-� Q\����T\�G�0��(�K:(����3�"-��1}���oÆ��������G���C�V��� �к�b��G��1�u�#ݖ�� ^�e�o�e��Y���D*NBF��N����rIK&��ǎ�'�x�(n�@��4��S�	_\����c�������req�*d�I� �"OVj���r�*� ��F��K/I h6���S�Dӈ��e�3����EK��n��V��E��PL��u&�>F�Y��x>oz�0���N24j[{���� C\�<}W�,����v�hQ
�m��X���hw�b[q[7�H���0��|��V������R��3�'�.'����q��/�.�[�t�A��5ᤠ?Cŉ�	�Z�u2���e��`�f�x2�XQ-�[��%��z]����y�fK�3��Lc��
��!���&��5}����U���l��HƳ�PN�_!XҞs��������AT��N�Bl_ȜR�6��33����	/��D�I������v(7"��G �����e]IJnݺP�ٳo�)�_�|�n�!���3)Yȁ�"��vvv�us�k>n,���]�,Q@R�X{� A���MC�#�ϩ>cc���;X{�4�R^�b��@u�9W�<z��7߬O*1w6���Λؾ��߿�&BXi#u�/~��s��w�+�����iO�t�,�i�s����ؾ};� �LЌ���C׭R{�'>�;w~��������ɤ& ���d�P5��������f3�;I$�Kݍ��#&������H �wt��(j���8\���t�"&/��Zn�L���v���?�~R!〻U*��Z�Yt�.M�FH�qR�f3Um���4,�,+v+��JU��&��)�]' ��.�S�4�m�T�f��K�������v��y�đ�����t�T����.d�&�Spp`p���ŦdP�tɩ�k��@���eˇ�I�c�=��O~�V�T�-_�FB��]P��Ly�EH�0�:�&��Y��KY�����SH�Ԗx��߯e:x�v�����\�-��"�G�6p�Tiq� �Ŝº�S�D�hHb� 8~���ӧt��R�v2�z��!��L�C?b�DC}��'uB������_���'d1���8��%�E-;�e��-�O~0�Pj(G��7�{�9@%��"%ba����|�+_����9?~☶+x֖��㵒����n�LfXԝ��sx1;<�U�%����SB���0�Ѓy�u�+c  �I�;;���e3�c�nC����Ta#�(���7��A��f������D#FLf �����&�&�C�C~��<xP��Y�ԏZ`ޜ,9�����t0�~KV�l
��0Ytt"�!�8�Y��sdW-��l�uR�4X���g;(3H�m���޵��'������ߵ��e�a8#%�߯Yu����[��╕�]����^k_��D�F�iď��h5D-v�.�.$�Ū����.�hʛ���ӶXq}�1�/XT?�x/u�o��v���;%��@J���N�@�5I���yLFj�3rW��Ǩk�7�_��h�N��|M"����)Pʑ1!�4��c�ӻ��b0�d�tc ���)�ʡ�z�7$%���j 搤>�o��5��X-�X��\�߈N�fh2t<�	�%�ł�����>�h�9�U8���*�Qɹu'��k���d�h��$1�ױP�J�<��
��|$���_���5�{��N
��V �]�Z�{�an޼Y������W^oW����(�Wk�P�q�:u��ѣ�3��������0�^wr�9bz�����ݻw���'�6�	��-��'8П �ý�w�%����β���f�;����$d:�;�-�q��E�Ϭ��!hC�.�-$`�F�!�2���w�K��Ѭ����!�����DI�ӯYߥ����D�����^����n�I�OƼ����j$���q��ÔăB{��H�0���3#�It�}%3����Z���ZSWg$�i��TI��*bK�N[_��kS�+���i$��k�l��r9T7��57t�رc���v�㩥Z�1ɧn"P�p�0u*Ĝ>��~�C���"�!����{��o���J�t�Mb$Eq��P�} ��8 ��/���'�L���q# D��t@V�]X�P3�G+��'}��d�Wn����-
��ߠ3�5�,���#r��Ź��|������K�m۶W���������?��W>"!}�7bJ��D���Ƌ���uN��%��0�Rqu<ζ��*n��HhR����?���G����%�����ի}{��.��x�uk�;��V�����#(��"$6&Zɋ�OmY�2\0��8�/Vtx�8�Y� �9G�a	i>�j��F�(�ja��ʁ�D59P�U�!`����]�CG:��@���<g�j(�$79��B�/����~�3<X�;��{h��8�I�A2D/�W����:�Ǐ��2�~o�7��;SGqzһfܧ���40㒇�L�qj��(�b����F��-�[Q̔���Y�D[���}#{�`�Q�\����xhx�����S'��f����v�Ʌ���a��L�صR}~����{����c�e���	��q#K�*N�D����O��0 *�o�d/���w�����+��ƒ��X�F�W¾�δYw���!�z�A��G��)�Àճ#��*Pۗ�A�]C�
8j����`_���D�}b���/�,�H�&��/�G�z�B,��ǧ�#�A���9���<4�]M��w��%B�PY�, ���<0`�e������2GhpN:X_�C��8�s]�6�9�"��d\�;��,�>�!X�,@`>����#ͤ��K��P� �z��k� i��c�	� ��_ƻ�:Z�tS�t�����gqo���^{\*�����g��A(J�aVˡ�Mv�\"Xc��!�ِ���`C����pH�h0T�Ҟ��`�YBt���']��i�J?��'?�խ4$�� (&
N��{��H�"%�+c������k׭{衇����2xR�D����ґ���=O=��ƣ�����}q�֭X�z5��������[�n��ԋ�w�}z�β�nǎ��R6���_�2[����ׯ[G�8�[�m[��[�ZS����?�m��{�{5WXs!��#ã��7m��4*��?��?�.��{�6A������O�%~�;�'J�Xu��~�Idd������������?��?�Фi����G�/�Z�ТW� ��v�&j�ڵ�x�@7ٳg���I���^Y����ؔ�������M4��ä	�j�BX�WƩע\�p��z[�$1��"^�<��G[<�����屮�rs``�?�>��}��k��`�z�$���NՙҴ���+8���կ~U;��?�ѿ���#�Kz��em!�����X_�H��kϠ�[q�p����Q���Z��?w���v��_������R`�����WX:���V�����"�O�K������r6�����W���\�_s���>���,�Hmc�v-��9<N����h�5�H�h=��t�����Bn��	PI�(4#a9�;�R�,'�DW��!�Ap"MaM�˿�˧�~�SS�vs�
N	���#5��H�{�9yښ�wҷ���$.V#$�F�31T��K9�Z�ZM��U�&S�Q���d㱴v���Bj�Z�?������FK���w~�E�E�vI� ~ h"�dtTB���֮΂��^�ڙ���F}�hm[Ʃ� �K�6Jo��˳�?8<�v�:��$(�!u�Z'	�}��}��t��~mP�B�dW���ēh�T��Ι�,;Ku�)�X������&��CH6����U%ڢ\.xҤ���l����B�w�6�OEM����ír},���7�=Jsk�=�fiN@�Q[��bQ�V��{��Tj��n�fVL}S�4�.C���N%M�o�}}Fi�tl�d���'�F��>�dS�q艜�kS3�x$8e|�����7�"��w8`#��x�i�#�;lܸ��a�e�9�7L� �\ét��@T�+��'�,-m=!n����<�$$���D���.x�S�4�S�1���GjI�e׮]�����H�����ג[�E)�e {������ug���]w�e�T��35������[o}�C��q�&����_o��%K���O=t�����ҕ���p`�ug����e�p�fz�'~��_j�ᬁ�C��z����-�c�=��-B/��艿���/	����W_���^�~}�e�@�_�F���&�R����5<@�\�^|��'�u�p��Q%�e5��μ�Hk!3��[o�Z�}%�_��N���ο2����ܹ���7ܠJ���(th���w6��K����>���s̜.Ӌ������,�
r
�%�@H�R^x�-�n�����5��[��|�|^��:M͞�B�Ңc�M;�n�������=d�nK�6�f����� ��Ѱ�l�aS_��,y��_B5t�K�T�8Z�K�� �$%t�6��BQi1�DzM\,t��)H	ݐ��]{I�����S헿|���������NN��E��6s:@����!��$��pZ�@�n�+ǜ����Zh�A?��
2���(�W��p�С�k�[�l>�l�M�+$��!BD{h)��CB 8|�X|��H6����lj{�a%�V����=�B$� ��~xF'�4�՜_{�K"&+!����)�\
dK���L�(�^>�܉�ńs����u���޽{�~�R��jJ
i���5�C�׶��v�3�<�|ddDNr����X��#F��h1�Q�D��0i�n��'g�O%�)�℩MṆQ��A����t�sQ�k��k�F��ޱ�����9�F}xt���z�J�Bu6�z��r�j�4�M��^)�yO͠� �l���j���Zm��¬1�{�mX`��X�:�����|քx/�*�I��/�}	�b#z�׫&�U������@�G���c�Ce{��l�=��n�N���U���ĖB�*B�������f��!ȿ�~n�$���>��N߅ԭ�l������9�%SY�6p,t�um5�P#�A���zo�D��m�M[֖y����#����C��6�#�P������c02����B�2L_G�Oz)(�"x�0
�fr��,�VԠ�.��w������

�@�f�u6�$�x�\6��I�-"
Y�i:cx�DM��&�x�%�J��G�A�k׮�[#�^�#��H#��I�!�u��jS:���]����c>�a)*�M�(#U/ՖLOYH��9k�[ۦ*��^k�貯���u��/��$e�A��q��ѽ{��p���sd7�݁��%ņí��U��O�jK�<x�����G�h��Q�g��1�D�<h��gɋ^�ٯj �����PK��ؾ}��Р�-�ʦ3��|�[v�U���2~�:�1G�Ԁhys�d�h��9�[�ʄ;�ص��<<���'}C����~�"���鞮d�����8kG�J8�֯��R:����VM����~(��/j6��Lo�tY�4D^6��<:��CT�@_G2h��Q%l��
�Qk@N!!��L��p���S���;�C,����B�rg�H��������p�����X�t����-�@�����}��LЅV���>�m`e�*���-��P�����a��> �$�����o��}�ݧO����ӧ��N'�桰��p�,�b͉E5��e@1��R�r�xႶ�)���.�b
��{�'�L��(/[�tj��s�+�!#I=���>~>ؘr��0�I���k�8~P��b�^3G@�-��p0��I��Z��5kVi^������_�5��rz�����O>��m��&E��Rh��/k�5	��n�������;�Z����/��D2*�a�	����$��,�M��n*4����L�>k[~�4cn��6�Eѻ̷�5��Cʘ�=a�s�W"��JgF6��y�'���J=n�Z�*WK�W��q�� jcQgP*[��d��5����֜e&H��Y�KK%׼����P�&�j"
�vu�P�IK�-_&)�Gh��0������Æ�����#�#��	�D�s��D,��
$~�j��͚R��iW�D)6�W�
G���ցѩ�m�D��FG�!�y�V�:�u��A���!�O�\+��}F̜Vk <�c��YA���A'4�T�RMJW{�h�G�g5����:�Rj��<�zݐ����	-zOݙ�B�K��O�h�j���`t�ӳ��0�d��49|���ؘ���c7�sY}��^"��敳�]���.��|&�&O��رc�$�O.;�NÎIyWJ�zq	P�"�A��F�&���xÄ)�V-*7k��l�mh9SZU)�a[��ؕ�T_���I�s�W~��6o�,�'�����@	i&��S�Of�� e��"ܫ�jV����� |��Ԁ5EL��������.�������Ʉj�4���6nܸiӦ�'OV�}��{��As����Э�.l��˷t��: Kb]n$4	�a���$_�u�n��e��w��lz4�����?yB��[�N�Ʊc���5 �.:R?�l�Y:X�l�t�ŋ�9CK���>a	@�*oRw��F��bl;vRs"3Z���/��@�%�ʕ�O���i#��
9@Y�<p� �MM����+� �ԶL�@��T��w�����5�~t�p�ɕ�lb�'�:t�)�Q1Ȕ�r%n� �^pjE��瀺E�Դ�0V"��ߏ�?��<����={�ho<��SZ����ΨI#[�PA��E��1!A�ƀ3ch����֜C���/���
{d���P��>��'i�Y3����k	 �-+.^��h��Z�%)�a[RR@o	=NA�W�O�XNO���T���p���'�C�^ˌ�! �H�L�K���
�Z�ǥC�� ���z@.���u��r���im<� ���_gv����׾�548����T�������W���^X�HRH"�MH�Yiz-�}�c -w�l�V�����ˏ� m5���\!ΚJ��
���/X�w�j�2ۥ�2�d�F�MG�>�X����#
- y���o���X �B��P�����m4�����.��ڎ͞ޮj��_R� �f��'�QN���XJ�ᬆD������.#�@�	2-���@�:{ʠ�30(b�^C���!���M����:������sM�0锑�T��;Q*�b��D�Q�'�6����PSb�ƇgY�D��Uɘh4@S�9��~$���e��r�P�׽��3=�EhS�I�K)��;���� b�b����� ���P���SR�����d���9����e�D����L�U�����_����a0�x	ナK�mX9��$7��R:���	�jSiצ��(�n����T=	�e��#�'l/b]�jI�wdS�Ė��̑������7H�fs�e=��mZ�U	����}z�)<$��1s�~�}I.����s��[�cc{kbu�}�����6� ��$��d@t���ʧ�BC�"���єY ���c2gm^�F��9,N9eL�#=|�ᇌ�R���Je���_;t�p���7n ��?R.W��Ug��K���ay����7
;z�����% �ZQ��E�����U�}n��&����jS���E�%��>Y*zY��viO	�Le��K�]���gp�2�:�%�>�lU�vׯy�yan��!�+B���o��TLg�,tuF�DW�[b�X.���a�tIo�ln�W��O�X�������ֿ��K�yK �~�-�f��K�j��%cfIe3]�=)FuV�b�B���_',��,��c�{�~ۢw����x�F ��6��W]�_n��6M�擪m�M]������h21�d�Z�tZ
b�Xss���D�k���J :h��mɆ�e�kځ[>'���u׭�d�w/+gl��MXj�_��V�e���.��&n
-%����&���r�v��'������oy���Ûn��/Z,�t^2&�㸕J��.M�֬y��C�������,��ۿ��ڍ����,��J%��N:��l���%C/�<+������X�@�/�T*���ZD9�Q�_�������Bn!I����8¨zIK
3aK�z#���33�M%g̎���m*+��_�����(z�>	� ���f���+hꖗ�V�)����r$v�#�D�ǻw�~�7,�����_�B[�K_��^��e��-=����˿0Hj�@�V�/_��`��Ã�ӳ�~��2rJ��LL���(t䴲�N�<n�O�-x��F���(o�o�D�0�����n�X�a�I`���b��E����C�e0���  X*�`P>W��xȗ��l�rH2�c%��NE�fa�����\4_ld=�=�#Z&�^y�g� Y6͹�2Θ��8�z +b�t�ɉ+����M���c~�t�˜�#�!w+�qB��� \cҩ�#~�e�	^E���e\%�O�r�F\U
�QN�6�d��.��?����?��O��0�nŁ	�`��^�v�'.,����7��6.�_�+-��Ŭ��OOĤ�N�T�Oک�AI�H�����ݷ���� �<yό���H�#�c�Z�����u���b���@g[s���׍��#��
;�_Z��t]X$C�������)|�-[�8i��=��!�����H��$%�CeTAo�r�	e�V2kpQt�I��BN��D��.���t�f��9 [yY�"=K3 ��Pj���x_Ҧ�F0v���/�,���ʸ�	�=5T�������
�%�]W�G���tvߕݠw�H$N� \�n��4�&^q�C��Y'�Ӱ��1]�U��K�^x��%JB�@;A�iC��zir����h��|i�;�۷O��c�}�˛5@�����yɃt�N��N�Ӕ[�+�n� �ꤻy�x{M��֝�WC�H�F����yC�S�_3	�����Sj�����h]����A������q��s�Q
;=p[d��"����L���G�J����5	�M[�L�7�|(T/!X����6��i�C�H2:f.x�X}����"�q������)]�$#V�$�*�jm$�[*��kQ40�4���:$z��}e���GE605�&���?�o=�쳚ɫi�����Oy��٩��He�.��}�ݧ���,^��?R�(��ų���<����1���h��<ڀjv�X�;
0Ʒ�i��Cmi&�R��&���N(b��>]ME�[l�^����� Q{A0bKh
��ӂ�P��,P���h�@��IK9+�6'Dl���e
���=j��{�nh1�U�%��������u�lz�'9�d��Ǚ��P2�GGG�G9�^�P��0,P�����F��[y�UG'�/Zb�bP�n5YP�ܪ��i����"ϸ���f���|�3y��4Q6d���1އe��o�I;Ղ����%��P��#@�n�T:��]��i��gZ`#Ԧ4oҋ��h�=-���?|��\mJp(�|��r�,���,�d�\r���W��X�\-�5�J�"�� �B��\ �{w���Q�M,r�J|bWIƂ@��r
N%��:[a��`����ef�HI&��3�\���$�I�(u������P�I؁����%�4{�������oa�k�ҔZK��p!�K@��_#�F^��F��D��Y������ ,v!�3ɾj�	�qϞ=&��$�`[�Sx_�+�5zؔp#�A҅�3a�c�D��)�CB�{�7^�B�P��D����Hײ��1	��p�Nf��n�L#|����t�[l���F���Ws"P/�F��d��ì&�7��U��Lw#�����n�g�9Y�o����3��R�ͮ`��c5Țuµ�t R�M���/���!�m9��24���uk',=���89���˼{y�wܑ����a�������T������S�4*?�Oʺu�ӥ���|����B��_A�Ў��D�f"���H��h�,4�jDb����kӹtfn�L��ٹ�gϙ�M�����9~��uK/}��םwz4�MOLL�w:% ��G(���W���JI�>ab�zY]	������>�,�R� �VͰ.��ǦM�dɵ���3�YlC�"��l��r�c38���GIҸ����&, J<U.Yr[TWj{������HA�^��J$`[%;�41���F7�mÍ�D�x㍃��z)Z��@*��X�~���*v�c�UyV�����{�Jy5�@���^�t��=�/.4�59!������	_��@��eSɌRDΠwLl�wG4�oґ��ˡ2,r�K�k��N�׊b��Nx"�\I�"*iWp�)'P$��)�EDkPV���lw#8Ĝ0$�$E�A�PX�ID	B [H�S����޽�$�����}�ӟ���̜��&�~�Ok�������x�;�d��&w@yK�PC$Q�Eq'~r��L�D�^k"Z�n�9�	���j�kG�qׯ�&W�_��-��]��^|E��͂��v@#�ă���9s�r����[f�h�\ϖ2_��D2T����10@���+tM%nD�M4�BD�����4T�v�k'm�tt1�Qc�0�[�I�
�6�|�+�$$	�L�2�K�� *�$�MT�DU�/��xG�F1Ů��c�If��5ڔ5nyi$hJ��pR�����[�ߥ��{x�	�Jg&�@���`t�h�S"&f�$�~��5`�NP�&����D���s�Fd��w_/�I���B�(�%Au��A�!{�_#�7e��B��(!.$���$h$�,��6�n�1�E��VpW�*��~X)�:0w&*]��B�$���A� �4��W4>Q�H"T|R��v 9@�і��u�M�D�a��H�
zA����Q0���O58h��	+�Nz(�诚gݜL����#���1����3��]f(rJDu�P�dJƓn��{CJ8R� &xd5����r�ʕ�|����L�j�i��5Ҭ�
�i����)�� �R��I�U��ZH�蚫SW����a]�`�t�"L��p~W�������0?GQ��Fn+�g���Fj��p9/2������:�Nz��Ν;�"�䆖a+A���3��'���u��Aw�/�C���&Y<1?�D?�T�gΜћ��(�E���{�LЭp���w^s"Q�W�qRd�J7�Ew�~�9*cZΆ�r,7�-��s�ApC��rBn��[�]X~d]���:��1q��@eV��?qbL����v�=����SB�^�[M������h�
��ݿ�.�H��L��i�`lڼ�%�i�pJ6�ǟz��dvW�Ѱ�i�,W�(2��-B��O��ɻ9J�80 ����-@Nk62,ϐz'���[˫���`�-� �B���@"5&�M�+I4�ĥ-�Q��A���Q����Jh�rc�5J�b��ю�ܐ���P(���t��I�1�$n�V��PqdB��U��8	�7�Xc��m��歏�m���s��,�L�5���?z"�yW�[˕��Yb���=�g�i�-�I��.hV-��y���\�Q/�K$����t񵳴Vq�t�&]"'c�e���� r����^�V :���LG��/G�y�W��y��y��B��I'�F�$�6���f�h�5'��;;Ζ-[�Wݿ��_V� ��L��d�cS��0@Ҡh���%�b�F̉���`�Iq��-��J��g [�E�;D1	;���h�`� +f�� eΩ���:�q�o}��;B���Z�D$8��`�-]������:�@ !���9^W�a��uO"�Ơx�!F])=M	~p��Eo7���' ��O�/o��$cH���D�{=9V�$, V�S'_��[�N~��!^\�˩]Z�4ˡ͉��K黴�H;?a<)��4+�Q��Bt!r4f�
ll"4X��v��&v-Ur��v����C7���4iI� a�Ɩ�/2J�]2����!}��������Cϟj�.� �e`��b�k!�n�JBg���l��;v���n������v2v	Qk��Cr�ƶ�'�f��c��{� �B�epd�����/�HQ�~g�p`�z5{L�Z*sf��6��+W&����z�U+G��j!��q`vʵ��իʥ˓:Y��	d[�����D3W��/j4s����r�[h�5ՈV}֚��8�+�``��b�s��3��sTy���1��dC�-��zҢ�HSA) XOB˜/@���S�NADH����Z����X'
�4���$cl�C��(�S�x�԰����VV�FF?zy��? z	�S�O�6	�,�'(i�[��\0	$dP�8B�i���=�I���u�I`��^zG\A{��si� R��U*���������;��v��1%�R��ֆ	%P��יnbA�^�����N@4w����bx����EЈ`�đ�>�p&�{�P���C�:��Р������Q�F9Ԓ%Är�*b� �����}_�lR����Ŭ�c�-�И��ޞ�_�p��"�^PwqR^Ř"�3������M�!jC�5T��U��:���uZ�f��T�!���:���y� ��,���P�[�%�w?܈��XTWL@H���ls��Ճ��\�&�6E"��L3��`mp©�"���E%
ϐ|T�e_|�E	�[K�q7�|.O��o��F�CTM!'�cX?�:[_F�H�Y��ٳ�ppd8d尽���Oz�Q���.�*jU؎T���O�2��!!����+x]D��CMg�`PD�J%�(9^�ZhO��q�����y�wo�ߣ�� �EXXo!*1�i� � ����.��G"@�k�굹�1���Oh�b$#+�n1�P.�'8%c$_��	5l����OR9��o�n�"���$�n+y3o��V�o �266��Gꙸ <]#Z"���-����b4�ys=�)��+o�o�-�.��D(%%ɖ����Ç�R�l�Y{�P;���7:�&�!��3A�a�Z����ӧ�М�;�� ����[�� l�/`"?~�@K��-8Z@�!�[��3o����C6�9qB�����/����^�Z8tuQ��~�[n�Ee�-x��7�I:���0X4∶��5t�><u��L���*|�X������?ń-+�n2���tM�����%���O����R*2�]7!\��P2	D�R@;-8`VhTb�@�Y=y򤶴1��L�:�w����@�a�k����� �����o�N V�m�Mq�u�i
*1e��2��;�z�J3��hf���l8h�?[�Gqh�vj��iy��)� /Z�����Y�)�L�=)r���she�t��G�.'Þp�]Z�%�D�^�4�%�ʄk�:�0��.H:Ǉ,�J�Ѓ�g��������9���?��P�OM��3����}���u��Q��4htM0��
M�5ufu�4���b�4�n#�lĭ0SNLqO�:B�B��1G�3�>Ъ.�I�;�_`��-�;t(�d/�7�B���Q�-�>�%2���?6�'s#��Yҍ��)do�A���G���Z���`4�
z1bk�Cqm�86	pC�V��ά�.�6#�V����t��2k�e��k�,ѻ�g�E}=��g:��(}�Z��+�V"Z(�Ua&m:��ӓ��P���ڀ��˗.����m�:����Aą+Ctό/���� ��84@�� �ͥؑ�Ih��7n�H}\c+4!�B�B4�:M�Y����I�=2�Td`V� 0�ԫ8�?�['S2r7�I!e���ױ#/�������LRSI��:���c���p.V�m�V���)���Vp!�8d��C�x굘��d_)f�ǣm9���00�#��l#�!\g�C����b���7�+�C܂ �:�8I���p8Y���TZ�fQ)It08���dĨ�Œt^hI��)�q�!�?�.T��P0�	�b�~�����9�;��=�@%]��x��?��q{�I�L��>i���k�2hx(���a�!���L������ӴS�Iϥ7N.k��?���jw_/�8�	����xlsN[GjsO��<�Gh�|�kQ��l*���[YW]�IлP����#$�ml����s�UY�a4iF3�κl�g�yf���RJ�\ư�ʾ�<꟭��:S�PH2�V����E�%�<0<����z�c�dt�0'~��n��z��4	ւtU���_�d��Ȱ�U����>�q�	���0�u0^�����2���@��)׭[���u�P�Fje�B�AA��[]��'І����<A���߽��O��O�:���j����H�V̘@�7���r͒�R-l/ A� ��~M��0����k8u��̱�)��9=�n�e�$�"��zw�!�P���3@�@�"�_Oqv�u�!P��F��~'
��_�d4���W'\������7E"1�\4Ӗ 4�d�Z��#\Ԋ�$d��H]k��GX�o�ҝ�qD�B+�g�A(S�
)�H�nI�:KĐ�^�"����{�ې8��JLD+ԧ`ih�'�U�Å��"�˹`�I��EQ��g���(����?>::27�@�w�MB���<W,Z5���ڵK�2�'hm�F3F��]��$ʶ!�a) ���I}�'�ƹ�,d�ި5����0v�f�E��5P���N�l1f�,�?y�1NH�jL�L} 8�:ߟ0|���/{�Q7�OK��o ���x��'N���d��o	��*}��帣e5����&?�B#	�g�7o�=���H��J��H"d�=�{0;(j�/���� b �C��\#�-�4���V�3���l/�)s���s�ƭ���Q�LVpq@�������# �/�h�Y��ɔ���_��-�i�2��Ǣq\I�M�/U-����N�j�Mڱ�ɱðV5�yv-��ە&�"e\���
@���8�������L;��E�pDW��)�qʦOH\jI�q= �\�E,<dB3G=]�B�����b���*�]��3�c*pb�_���>�^��;����Z)�I�"�F»?�#��E���.^�V�8�dKq��L��jK#/��'�3�.�����j���%��ҿ?�=�l�`KA��~�� ���o��u�V�M&���ز��Ν3=���عs���Kw�u�ƣI����SOU����ݨUq342�P:�ӁS��5�E�nH˭i�~߀��R>r��k �@�'��Rd��i��D�����E0�ĕ~���9��\�r�6�����H%�^ɸk��0�*���+�_{U'T�Hc��	IrNu���]g@�3gq���!cy,�	�ȑ#�<�ell���n�"���g��������tutd^{툮�^�j�P�#�k�'��!s���h7N*[��%1 6!_׬���\�ap�`�E$���g�X\����!�Q��\n���g�0�I��R \O%Vӡ�x�z���>���Th��wd�eg��F��u��f�Q�S�@g06 �U
��%�5N0y���ox��2���Kl�|�ĕ	��I2�Z���>����\21uunӦ��/\��.����o�i�B�D$�>��l�曰GIOC��Gc���rK=zrr*��mٲ���(z�p}�*��d�@���a�0z#|���s�"�hD
�<{�{�2�r"f��9�����L5t͚P]�eP�"�<�6��\��Uضm����W���/�+�c����2�6?��� `�����}�Q���O�.|i� PSEfB��~p�ݖ�459����U��X3�H���x����1����v�(Qk& � �faIk�5�F6e�J���ȶz�z��2�"�J^�r��w\������|W�<��hVnܴq���M�[o[��u�_s�*g�j��$K�	4rK��ˀb��9}��6�����/��z�Hn孷���k�]����/���74|���lqa�T����DOL�~-t�TToUQ-�KV���VRo]Yba�Ju����:�:���z�m�t"Y,3�BMO��S����<nP�Z5��g��$�̩�̦�����犚|����f����-[6�Y��a�@�D��4����>��W�A�C��V%���Bi�4ɘY$�.\���!UA5z�3�L�%?�ΥS�Z��N�$��W͹F;��@��;=�B�l��s�7� �P�z�t��4�j���1�.;>>/F��l�y�\,�ԕ��6�&jH<K�W&/�Kq�\)�v�����Zˌu������X$�R�U�-�l�I�"K��v� Ka?�5Z Xܚ����E-$��VG�g�;=k��
���4����¼��藍6�s�s�'����w�F�����d�C���]��R�M��]�z��t4׭py;�)-録86���\�j�L_� 5~}������#���:~�8��V�TN�E?P�e���;&+D�떭��[*��驨<?7~���-�j>���t/�?g�l�/%�)+���{�j$2�4���J�v�mmҔ�68p@�h $��,�@����=�%����'���8#�و����	�ƶ�߅��fޫV��첧��Q<�^�r����=��%z�#.�t��EmB햍�7��O���̥��҂���ݠETi��e]�m�6+�r�O�ҥ�y7�%EӞ��_�n�\���@׍����$��z�le0�Z�;vH!�&4�׿t����D��A}dJ���z/�2-Z�$Ss3�_6��t[&+��}k^��Op�I�SΩu��a"�2�4�,:~5�� �P����uOIr}��/���!�Zg�� \���3�{-�}�\�d��Z�ƇjT��f�V:��kr�؂8��En��v����On�h��l.�}���F'�s�¹��>��Ȓ��k�O�ܾ}{W���Ϝy���Ņ�4Z�~-u?6�/{SH�."��TJG[�\2b���B�#L֣y���+������E�h2H�c�X�/WX�b���CUw�^��r��?������Ͻ`ެ.�螜5�����"�S�_���(�M���vW��F�hެ��\�e�3�ټxႡ��^�(�F�n��s������Q�Ԭ�L�	
��qC���S�Q�Ҭ���0�Ë �@��\M�z{�g�˯<��:L�֪�W|�Od3�Zݲ|@��
K���?��HV&Q�4J�%U����|qt~6ْ�T�T���ӬW��B�ڨ�+�z��+5[�T�R)���$���V��7<��IO��Q4d4��,`k��i��Q�ԝ�����!�t,�^�9"4-�zcwvh��k��wwZl@&ީS�4��H�������7sͱ� � `����utu>��:r#/�������cȞ��w�կ��UJE|�Z�MǱV��}����$����!(<AH�a#�����:m���k�,�LZf(�Ƞ鞺�#�� )�e5�TK���(�
O'O����0���.�T��2��gI�h޻wtt>L�7z��0*�Y,@�जd�b�2�Y�b�m3_�I�e��P{F�����~aS%ģi�ԏD0�%��M�w��QxD7�_�Z�NpJ�$+��5���PZ�V�=.D�@�	�P�4�f0+�Fjb� ��a�a�I-��cٛ�x�����l�h]�+u������ǉ(�A
㏂"����|Q)(@u��*�@���R�+�N�2�5���������t�okF��~�*��G��`
�9	/}���͹������;�7���%VM��N�/T`�e��
����ʘӀ5Q��\������F���,N��uKmx�K�k?`�<x���ѣGo��f]������^�w�9`Gj��>�Z3�XKGk�>�/Z=�fգGN��j�����K�Ѡ��;@m�VyϞ=�mFZF�/�U�RC�vFK����p�IL:�:1K�Y[N�@�Ф���8%�c�� ���,�B���3��^�p>$�[^PΝU����>�ʺu���^�q�ӔFEpqÆ�S�+9A#<�īBV������e����P�\[Q����[ �hW�~A��d�d�Ak8���P��u�8�;�K;Ę͞f�0$�7����C� 5��V�x'o�3KE�Fw�C����d��` .��3
KqsҌg�QX<^��/z���И"��!����4Q�V�W5>�1� 8 ˆ}�۲R���T�{�}�j8)��tH�C`؎�L�X,�~4�fW8���P0j*kN��Ў�GGZ�����y��Ww����O�]�Z_���hH$�,:�4b���,TׁK��_�f�|	v]@o�kG�+J��y��%Cw��!�Ph�f�%���c	��jPS�3�օ�(`Jt��-(A�3)��0�R+��@?��X]���_��MД���?�я���q�����=x��wcxi�id�#����3�W���X�n��m�v�Ȋw���q���-4! �\���&�0(�8���9H"\d�k\1��AIT��^x�[�9�����A���#L@­$�#�`V�З�K�E�8��l��`8��-��XW�0�CMj�$}x�:1<p j���ړw�W�%h��Rz�6���;��P~wy��^f�;�1��d�;I��$F'Ө_��PB�(��Z逐WŜ
!�G瓲�J<�pb�p�+h���Da"J���GS�Bn�	Lg�XAvŝ!�^U C�>�:>�6H��J	:�E��%e��)��Y��kl�6%U����A�YĄrN_N<R�"��^��J|Y�U�V��=��#���1��7�$YO$�v����Du7�-[���#�G �o��V�ח���HS:rm�� f�w5i����ԕ� �X �Vײr��G]ƹМc;ʦ��R!|� � �C�#����oz}���]=r�Cx��ug�Ād[h-N�8���/�>�.�=���+ӈ���pX�F,C1E�^���w����^���|���Ή&�z����C3�tܕ����p�j��pr�z�V"�e��{�Gmll,�,_T���_h�H�c�hLK,d�ꕺ?�'͎e�>���O�q;�0�B���船L��4���@�YR���.-g��v���_�r/.37 g.slG�8�ߴBuW3&�ƞABV�_|I^4�J�����8E��MuR�#".�1�?�|E���R�;0�A����4�Z������7[���������3�����<]��˦�tc���J�c8�@��r�E���E��# �4b�@t"���F��G�j�O�<���~WJ`۶����S'�l���C��C�� ��c��`��MļZ��?�t'��N$=>�:ŔQ*��YbQ+0��P���\\�h7�q�H¶���6߱���w~�	��hց{ЗF��c��+lI�f�z� +�K�5B�42b�:��]^2GB�&A�F���=`*�9�����#�I
�СC���S���-�F�[�b���{�"�n�b
c�3o#�&#�,�B�r��x�P�� �*:��;�#GA�' �Gj@OE���\IƇ���ֲ00�haA��G�{ �u�w���^uԫ-[�$w�Vq/��!څ!&$�&!�I�drI2�@&��;� 	$7@Hb��	�6�w˖mY�eI�lY��~ή��}~{-$g<��}�^�]oy����O�b|G��$�O9#�aD�L[A_�	4�補�a3疰�c0����f�= �J+!�����ݬn��HQ���n�޾������rh�� �d�˧s�@1YN,�L�*�mna2��_~��(������09ZWs-x�7l���r�Z��̶2T��ep�Oa�k�������g3&!��/�`3nf���]r�% &�a�jƌ��H]���r[�c�@�u�]�\�ر�o�EA��nعs�D��c�@:���P$(�������>�^7�J��	5OEbK26	2��$����Z)R��K�:�7JsYf��X\pߕ��/Z�����[�P�Q^�F�!��ʕ˥۰���
>�S���O<��{��<�~PVS
(�����@S��y�y:c�&��5L��A�ǥ�Z��P�]�P����>Yԡ!���/k
�e��<�H�r_�TH3a�, ���gv<����7�k�M������\�}R�jM!i����&o.3�����)W�ktIM�G$D�ܐU���>O��ߺ%/�˚�r=WFC�C�_{�è��cn���ul�S�h��R��>�ԗ����Y�tٺC [��	M�W9�x��f�g$@<� [n5n�P��֬fQ)�����y��2�S��5�Vje�Y�@��L���I�g̗�úL�MI��"|qZs�]�1�,]�ּ���ų\VySξ}�i23B���
n����s�V0�y��D*&Vd�<��Y�uX�l!�ֻ�+�R#+4T�*iuS���K�='��@>���S�����M�����l�֭����|��G+$%��3�`����uZMQA�j��,%oNM1(�����/��vBm��1_)+�)�9f�o���V��ߌ����p\�Ъ5�BY���bI#C�%B��ή�g�͕BQ6:�z�TR3��Q.�JөM��{Z�0me�ӓSCX*_�җ�F���V_s�5f��!j�R��/]62<�鶈�����VJ�z$�"D��әς��������r�mOj����2���@���\�u���U��ɳ�g2�%�+f��4�æ�J��hFt��QS/=c���ZuW}]�(�d2B��O�<����2Q���ln��uuzi�[˦v�E��jf����Sr(�����V���FOt�&�V��_�9!�)�n$$�����S^!�|�+�%�:󦿊�;
G��}�fV�kD��ua��m:�����E�����|�]��h��z恵�>q���"�L�#>�O�]x�YQXS_&؝13��ȁ-�%����mj���E�2`7m9u?���ؽf�����^&���Y�[hݺu�W-b2o�$+-Dr�z=e�|2�G!=yw^(�.���b�n�#g"�E]�/�Ad@dB8�7oN
>��D��V�*!�K��nD��ʡӜ�_N�x���& 2*���u��s7x�[����}��a������O%�F\��s�=���/_��V˗.�q`nǬ��N ��}�����_���g����?���W_�8��˒<�~PN�Yዩ��H��g �@���S'GM 3 ����Q�+D�V��w��]� "1��+�����!�������<�뮻���o���/6EL��ٸq#w�z��h��5A�R_&��K��͛�X���F)������~Q�r�B�>���>��߉�����-��\�-��dl]e�D��#R��sx�C�,#7�!�^��dMyA3�D$�l��E�#0z�;O(�Ѻ
�FV!�-��JH�i?9�\F��E��٫]ѣ��;���Y1/ud���*M��f�_�6�����͌g?�a0��N�Z��*]KY��<��w�{�JF�)�r�δ��G��?�!S�{�ÕrvG'8��Ѿ��o���?�u��2����|�G,e�_�����Ӯ�,F%M�.xHx�:=)��Sg�y!�WX�zҵ�e�1Q��Friя�v�s�j�V���<�����R��l�P�M7���j����Q,��Ɣh��dSZ����$7Ƨ,�ѡ�R��$$��O:91Q����E�!��X��~�i$8&X9����$ӊ�\�К�$��,7�}WWw9뺭H�ךVQ��8QC)@��Hot���Xt)A�d����pz���
�$j%�}�_���,*$~A��֪inM�n���o�X�P�Ua�xNK�F�<T�V����Ϥo�����`�5JڎV$"E�6}��e����ckE{ ���I��غ�M^nd�j@O��#Z�K�ў(�E��f��͒:ʐ�6��`���������.=,L�-[��ň+��B�@+�kˬ�$m,ð�	7�jݙ�S����	���`#��Tk�V��mAN�K֣/Ŧھ};�p�78���X���kO[v��P����A��H>^�[Kk�<3+�L�ŭNCݰaVl=���<�Si�2����4s!��bT�+��KD͠��˕�C.�"����C�ua�{-��IvT���x���y�D�)Y��^
���1H*v�'���W�P���2�"QF�'����>&�(��9��^WŲ��`,�'�`\g4��C��0��:l�ڵk�&�hi�O������9obc��uv,�˵�^�Pm�'�-w6��p���󆆵��fH~�`I�B���n~�ܬ%���BRv�կ�+迴T�awD;���ߠ�	�9r䘦E�d�D~т�9����t�Q͗͝.:5�mI1cR�6�P��Y�)[pJ|�K�^}FC3���4Q$&,����jz�@}۶��8�|]�>��si|��Tf�鏘����<�U?�h&ky�q^D�q��!W
�)����amf+hMRFo�`�T�?5�C(�<L�ˬ;�M�0�r��\}b��']�b6� ˘�>$��HT��B���7�Hx*<е�"S;�~��V�
�#�W���9e�6mr����L��0�Z��q���#bӡ�
���7D��b?s�ه/g< :�2��jC�B�����K���?׷�g��V�UiK��Ͼ���1�;*�Bkrzjl�ݩ:%��n]ݝ��)Ϯ+�������?u*u����V���K�	aU{7q�ety 3!�z�F>��c,hN��_��I���AH�D�!��3V����zb�c�4��e��C�_0�?Ph&'��=;7͋����Ȭ�vy�_�����\-͈\��p�1�8�֍�c��}���� ]Ħ�����V�7��5�̯� ��XpA�8o^u������b�RƓ"-������y\__?¥�(H=

�<��u�Ί��h��;t��
�S�ޚ���i�A)��U���u�O
5	5�7��%w���(��I�����e���ON&��si$�W��	��s\Nt}S��P�V`#��E���?_-��N>|�m#�߼yC���]]��U��?����-K�6"���}�\���/���
ѦI��lt��Lr�q�X��M��C57��
�i ˙��Tk|k��ݻ�v�<K���sٓO>�ZS��*�W�G�Y��xO� �=�$�c�F�3���@2�o�_�+���_��ԃ<ԃ��L��S�_d)���Gartm޼���bxLBg��f�:�G�#� =�G��\�����e��cq�q=���cѢ����<�虽�ԁ�$7�pf�U�C]S|��r&Ź��ez[�o�/����:e����/��GE8��h�V	Bi�<=�2���;�-��v�M
}	�wU��$�%��Ν/aՠ�c�������ʋ.�(%�����{�l�_ϥ6ުU���<�Z��0�s�+e��V��x���\\S)L��a[65�V��̀��h?=�r%{f�}�JXyRȘ��Q5ɼue=���b̢C�R-��	m=�f/Ԃ^��5�`h��9���a�A�T���f�Jē��}���:P�2��{hf�9T,�l!��Zwo���ؓ�\-y���FQxY媉ba8yB��[�:�q�J�@�9s���I=@����ya~��W��S1$�f�� � ��`'h!8���g�yz����މ�1�{LȨ�%g�W����ܤVF-�ʊ�;�:ó0�h�*l¬�#W����F��&���Bﴪ��0MQh ���rn������o�?�P�U3��b�Ϊ/'ŉ���tY�y����R��HIļ,���S�|J(5����'w����hb�&���s��x�	���>�:~R�\�㥌�,��i]�v���eN++��kj�gL�Bgנ\��`Z�b�tZt/��E���==�s��B&@�[�,�SD?00��ڞ0��b��0��w#�q5Ӎ�����зU��\�q��$�g<6�3Y��Ō�ǹ��y":ԃ�c�sR
r3笖E1��*��RI��k� iY8�	��3���'*M"��h�\0M��;�OÝ�H3->K�Q�yx��J���&V��#cka��u ���	���[^`_�*��n�W�d`���Z��=L�v�J�+�b60::&O�����
b,Sj�-�F��oI����!�[��MLd |�d4n2K��������� 9^�T'v�
��B,�5�n���-���dl�%�B���Jc�0F�;?f�YH(�=�����Q}�ՂL�y�����o��L�vǞw�yz�%��L!
LX)Da&�=�8Y�2Gc�#p�W����+�
��y�Td<W��z�|O�t�M��fԤ�GCF�=�_����L	����g�ur�⌓�B�C~N;�q��H�0�'$I�p]]�`�q<=����cc)r�̘�hdmݺu��̪����,�����n�e�8��-��j	U�9�S�d��)����KqL� �d����v��AV�ߴn����I!����O?��Y���y����3�\Q	�3�pty���7�(眳v :vxT�M�ʆ�EX�"�~
Y48��^~yO$����Ә�֮r(*��y�"����J5GXF\�`�X�K����Qg�3i�
ywZ��au����f#/��T�
�<ՉG���H�6�F�ȭFF�8���x$~*�v���.3�##�&�����BaD�#��[6V5�F�gZ�"ӀWmq���rP[��t���]]��v�J�T?Պ��k�L����@�EF穻.O��g?;��֬Y��Q/�L���@�E6ڎ���E��j��L�@x"N�B�>�yLVT��<~*���Y�������6>+�K�����m�;�m���'��,Z�l��F3��Ug�/\Tk���{ub:��,6��Ɲ�L����>Ѯ)Z��Z}Z�f%K�����ֈ�#���e+9�K��4Yoy���Ёߑ�Z�ޮ��d���kBzu��n�R��+��G�6mD���ט���
�=�Gr�)����F�t2��;6�N�?.�8)�'�PM)c��x��'�������+�Tԋ�R�u�nG��3	Iך�mfԂV��&�����(���ywx��h*>50��Eu2q���&OXmv鲤�k�� ���E�dǶm�
��C��:BI�lB�lt;�N5yΨ
���m��K�yd���RZEV���h��m�X6���zC��U~�r�,O���;: Y��w����+�3a�Є�d��Z��]6v^�Ld��Z,L�s,��mD�/&�(�Eo�3*(%z��c�Y�<z�@��.��S8e�u��J��z�4HY̝y.��&��۲4�����C�����2BYs��7��](�Rl�B�ͨ��"�&L��
(�yiiy4X�����O<��/�F4�J��9en~��V�2`p��իo���g��	�idt�L`;;���oF@S2{sA1���k����n*7D�R":>�}�W��{v���k���c�N!�x�+W�l6���y��Q0��-��yDW��׬��-����[���O�L댕��+�������y���	���y��_z��ʹZUݧ�~��_J[E�����3�QT��F	��R���ܔMJ��Z<6	sr�78Hk�y�c�$e�y�t�n���?(�M�bl&B��t[@-�<��s�s��?k�0��6�̍dE�)%�bV�ԈR-�"�\_�ϤbX�ͨq��}��OB�\�k�z��,	��`t���}�|�٩�;��D�i��(%���/X��I��Bf,_�"��:5��E
E����Tta������B���v�?H�=JJki�?ojw1YM/D��iJK�����h]�,�3��9֨=r���/����C%"�JWt�(Z��c���׿z�-�Ȑb�՝)�芒�Z�>��3�Ɉ�\�*1(�w�65U�іZH��VSbAU^jP?��xJQI��Xj5��~	�f)�Eo֣0���p��ֽ���PL��J�r�V�~�8_ƣ��!M��iEoo����֚���.�O���9�BT��M)��5�2 s�EV�V�^w�u���뱣�boiJ��+�4�*q�ȝ�IP�K��Z
Y��/2���%<����2��c�P�M/�]�F�E�۲x�Zֿ�y3�B���[� ���j_B�h�d��ŉ�N6��X�.Z5,�>X�nK<�����L�qV���`���Z=d�Yg5��)5g�`kn�E�h��Ԝ���'S��4��~x�\G�I�\���̘�$pѱ*5���h�`�t�y�<1�WM�����A2	�ėj���P��ۙi'af�^	�@�X-��1=5�/�f��W�hN�M��%�\�q��tI��ޝ�;4���DI��d�=�"�b�����-ʚ�8t���3�xMū2��C��r��4��͏<�z��؝Sv4��A�%���@�2g�s���I`��K���a��L]�>���\�!#�m����}���0�x�#*�����7�����y���������o����4y�������~�Wr��ۿ����d�-]�!��7����^fםy��)�ާ?��fp>����}�{o��&��l��s�=��b����/���������q�7o�ʬnڴ�O��y�����Q$�����'L���&��>�%x׻މ�Ci�2Q �ħ��u�\�Oɥ�m�U,V䰯Xʟ��'�l��uv2z�`�fi�쪫������עz����7>���fU:���7Ēq��ے}Gm�b%
�}u�Nн��H�a� !�Ƙ6�+<�]EE�?-��SO=�9���;���Qp��	��Y&.І1gm�}���պ�� �Ճk�P���PsN�ժ��>���s�^�����7�L�ߚf�����:�u�Q#��X���bԼי�x:���Q3��ѵ�1o�"��Q_z�m��Ԃ}S�Ä 5��'U����Z�3j��?�J�/"8�ف��!�b̏�v)I�ʨ�uG՟��Y"j�I��a��b�@f֏���19��/7R�[�S�R��9���_�󎟰mX)�xb��oFX��SʚQ8��=��/D�Z3�L��C�Z�[1k�S<��2A�B9��
a�{�E񧽯�(b��\mr��,�`���
�pa'��F�S�ͺ����F�g����S��:���]^g��U��ȫ�dL���aP���DR6P/�Y�ӟ�T)6a���}�C���SSa���5ϣс�a��ާ�O�2�FL\G�bF��E��ݥC�]�|ԧ=004�5��x�:�����z%+ʨg�'��WV_g��B\X���k�a�#T���[�C��6���36e�����Zt��]��K�YV��f�C{&�����"<�=�5�ۊM�sØ���:���G�_3�QG!$wDÖRo/�p6Ϡ䆊��U�&�W�]����Po�-xs�x/�	xqy>��.�'\yW������^f��T̂7�Tf�tE1'�XF�~;�j\1�+��#�j�;�5��b�J4�*D�0��dɢݻ�G���DW)S�&��_=�������c&-K��"H%RX]h��yx�����u��0����T���F�ݨ:�4y:����:.*CM�24��v������za`k֜�w�k�"�>i�o��C�x6��W_mm��1E�''�"��L �]�v}�k_���g��@�H��뮻�򖷠�/��Bcx���^M 5|�'�hn�;��A� �؟� |�u錦��:.Ĥ4�ϘQ�S�S��/ޟ ]r�+���M_|��'�x��ھ}V��ը0y�2 ��Y���կ~�	a}��w��؄ZzR9�Ř͠.ѫ��������7D������'��g�:j���Y7�� N�8�g�>>g�H�j�k�>�c���֧"y�����F�'�������ڸ|4G?!�g�JjS�vI�.���^{m��CF ��C��6��C�ذ܏G���A3RT�v�Mx�U7�L\ȇ�c[��wfU&���t��g�F���%7Qbh��4O�5�������;Z���������0�M?�,؍�ՌB恰^���<�͛/�[ڥ����l��A�cWb����٩�ɷ�����L`qՏ�n��㔹��e:sߞ8���R3B�I9k#�cB;<_,��F󌳙��ŚV�7׬9	���7n��w�������#��R��7��=�Ɏ��
�tUֳ��Hj���zp���C�<��'uWL�q�^�,%��VV��N��Um��r��s�g�r� �k5�-�<�M݃r����MGE��i�yثu����=�S-z�	�m���ݤfA�{�y5 �~5���}���?��3SӒ`z���o/D��Ρ#��')
�:~<Q2�MOL��Y�Uu��:�(��r�]+e�.�����N�xq���Lp+�*A�ᥲ�`-gŭ�i��X��SÔ�#q�e�6�Ό���A�tY��s��[��#WW�}$��]��i��w�3N}wts3�U��C^�f�Mr&.v�>6�rdR��#?�Y��ok�d�DB��)G��Ƭ��GRUO��2SX���P=��|��Ï�C"r�����'�W��=U��5�%��k�'V"�_��][�܌jӔ�e^�J��A�KA�? Y�c6���F�U���K������'?ٽgW!k��%�1�l�2�\~��8��.��x��N�4�ǀ�ؤ�;������f�t��(]��~3���k�'� ��$�AL�:�Q��gJ�[q&�#d��ٲe��t>�������Ӻ��V��i� n�K1�M2�M�.ݹ����a�/w��Q�T�a &=(i������я~�c��J{Cː��먉�Q��s��w��a$(cd��`�Le�Q��'H-=ЭHO�+��z-�Q:�ݍa<���V�L��>��1���k�M�cc��}�Y�Ʈ��*)"�sU��K����
���7��N�[���-1�Gլ����Ƴ���aي�\r�I{�`��,�i ��g��i*������ ��,�u,a)��|�9dg^p���^z���F_�IX2d���-+G�{5��LP�Vz�mo^9�`��	Yg �"Vבv������6΅a&#!S����٘��zT�L9C��o1l)�̚W���! /�d�>��t�Β}.�w3�B���G�k�l�<�=l�<"��y�Xd�
M���*O�W�iz�D��Uu=8�V��ZޛR}2�smHNG�:E�f��G�a_�n(Ƒ�����JX�k:��~�5�`�w�БH7_2>>i��w~��l��~������0^�;
ԦO��띝��/��csV�7L��>)p���1�1{�M��Il�H;���H j���>Fx
�B
Ow��p�O*m�v�G��(	�b�F�kMLLU:�6#Jc��+y��G굦f�/�N.�p<b\�ɒ�t<z����^�����m޲a*�szj4jS�3�o�@��:�}`�+��M�8c)�!��fb��)�g���Q�������#�'14��e�%(�VC�5LR����G�A���3�uDo�ي5�F��&�����̆1}g&(ak�Edh̴!���	�rjk6X?����b\þ&9js��@�ǆ�m��@͂���GD��f|����_�C�x�L"�׫yn~gW(�^�9ި<::Y�]@�H��������<0σxW@�	,D��Mv-9#h�[���v#�5�k΁�>�{�&&�0'�!���b�`9���a���<q��ݍ�����Q?FX"a��?:��7��5���)R����c���?�cJ���й+�1Й z�[��{�n�
VS��w�y��ʙ��	T�ͪ��DC4���;sJq�������W^ٰa�~۶m��t$�~�p�ક���<ר���ñU�s�QT������J�,Ms�`���,�ɺ�p�?��?��]�� ㋺Ā;��(�( ���/k��>�˖����K�����żԛ��&��D���#�<�rr�M���ƈE2i�֒�ĉ��3�w�1z"!���I	Qo����ַڨm"�I��8�)%4���F���M�4���T�a*��o���������o���u��1�1Y5�dw��-L��tf|�.��)^S������?�O`�ڵkIt@6�.�ӡбjS	ZE:τ���D��8�,����ƘKA6�f^q���tn��T�>b/����7�x#c�H� ̀���V�m�t�0!�,��mm�V��nk� �R,����)ߚױ~E�s쬸�_>L+&`�4f�v��$��PIG,%.f�\�V��IG����}�����Io�3I�PC�8$��sqx~ʓ�y�Y㣧��Z)a�p��F�o9_*��5bGF��|2�V���6Q�Q�`r�d�r��!�3:�J�;�3��jI_]#kP�6z�j:;�5����bV��2BvP�ҥ�1(#|��DNZ�fx*����zsO���CW3��	!?��,�3�k#ŋ*�V��UrJ�R�TlE׏�ij�Ӵ^�t��W��t��?�U氋�ZI~;�yz�A�W#�r��hח:�:�R�eO���qX�O���Оv����`b��CץI�t�S)k�����b۷oek%%]��^�w�o���G�J��#h~z�[y��Q��(Uf��#�m*V`kZ�R͸��*H��g�C��vw7u4�Z�K��s������BךeA�=�P�+Y�`'�ȑ)�)�|��ܘT��͝�<�r��J
�1-i��S�N�)�������WC��bu�c)e�;���nYI���$̭�������ɍ�!�=�I�
,��JՆ6@�!����(P˵���(Dɕ�B������%� t*�YM7��\!%j��~M=ϳ4v�1��\hF�E=���;	<ne�R@Bv�����o|��6[u�C����/���_���x"�L��=��s��Ul:i��*9����R��b4֦M�3`Q���'�f��f���t{��1���Z?��Oy
�VDr����z�`�����N��y;�Fye[ �W��f���T��Tɀ�r�֮�dᓟ��W��%&3����[�����T�5�V����g�g쫷��-"f5��[*`7|���6�j�Έ�{��������?�� 2<�)K��@�13���򃔕��gդ�}3��ʚ�`ƪA����\|��v�4Q�~��.��/~�@F&
���۠i�������7<σ��WL_�X�'b\s��I"2��C����TV����v�Yb���^k�D�G����xl`�~��*�A=+�ϒq޼��{�G�h�_٨<�lE��)�O�s�G^Cco_�v�!�s�~ʘ��ꍦ�@[� ^�B)�ͬ{b�O���MM��Sn mx��+Y]T�zo�n�s�J�a�4or�Vt6���k,<O0��=���f�
Dn�շr�����FG���:{�FΌ~��5���G��,h��tZ�J�Y�F��1kOww�YDѭ
�Cf8EͨkW	��9V�*��]?���:(�ܰa�o��oq���*�F!kta�[9k`ӌ\)7��Q��D�����CG�����`�Oz���f���pMB>�d`�r�z"�W.���i����N�Ζ\hL�g�5���B�h���I�F��l�m�YX������M�ˣDS�J�K[&"HTъB���^l��{lfz����Ս 5��=�yHt����yjT�R�42x��E�[���m�������Sc��3��$C��.����q�Tզ,(���ofM�E��<eq9kf�c�h��N��i��EՉ���VʻX��ң�V0>�P�5M��A�C?�33���nE� �Ք7���	����5�̪�j9~�rz\eQ�ԨZ^f��Zɶ�2u$$��IV��KP����A�?�'���Wl1~3]�f��2���pN�h�f3�QϚ1𡳪��˺��
{-d�Q��Ϣ� ��"��.���ȡER �XG��8|䠎�F��lUff�N��-^�x�B�R��ȣ����Z���Ը��N���i�Ze��ɮ_�B6�y�7�|���Z������#�<�ibHg�y&Z�|;Myn;����g�~y�	&YJ-��~�z�m���@�]kAdl,��=V�iDe��mo��B�5� <Hw����\��m�2.��h�dK�V�HɛY��B���6 m޼�w�hdL���7�y��ѕA ��ph)�w��R)c�3����r�*��c0�^�9y����d����4~gB��^��a$B�	��_�����#;<8t��ᙨIںyK�X|����koQ%�X��۪�H�ss�N=4�.�椝��h� =�M����y뭷�<��=�&�7�p�l���4=����ͮZ��:D㹇���nf��=ɤ���LW]u��#�U�lFb_Q����7�����P�&�ӂ ޅ�0	�v~O2�AK��8�٠�Ӎ�5˗/3�%�����?x�N)�F��]1���OI�n���S��"A	@�?Z�1�g�y��t��|�ɶ�f�{�+Z�T�iXS�i�4���0c�d'�*��U�fR�/l�+� ��P�bG�ɇR�(���y�&�t�cV�X��+ˠ������nHp�\4>p��f��%`��e��DPyc"X�bd��nE�R���b�NGFW�: ըIۚ��=9�P�	r>9�Q���R��1E�y"{O�x,��,���B��_��M���g"�jBKQ�q�fTn��� �t���J��.�tq�hT-r� ��=��(�di���z0��@EYJ�~��tp��������oM����%��I�ߚ�4�R�rѡ�}e���ćy���]��3�qx8�"�,�*7稼�o�@�����/P� �LE��b�����Z!H�����)�4۝R�Pg���oFN"����8F���B$�&O�M�é+##Ջ���k�Ra�%G؈���Z����2�V�&��eԹ����mĔr� ݙ5��Y2@�_��gY^ZA�y� �tT���s�4��	�ˉ��������?�瘁����;��u�5o��eJi��C>d�T߆��Χ�όQ~��^�0jt�ɇ�B~:�"�@=���L�C(_������&;��=�hv[�CM�O�]�w°���R֚-a������كAQb�\�+\���)�lŖF���~���û>��ϩ	�z��bw�)b�p�0*�L)�~�d��h2�M�.����۶mW^y%�4�P�= ���%�����[Q���|�I�[5�Q:�Zsv�aN�Y�`�K.�D���_~߾};�V�c���wo����g5{1�o��nW�-���6�ɩ�Q4[����K��uG>�?��ĥ^�	�}=z�h��|��JW�@$�4�)��{�-��Z�
l�M6n�hӍQ��4u]��l�K/���������O+@���[�3SʓȊ�9����2���T�E��bnn㥗�y�}��1��_ւ���9ԗ�*������7������t����p�������E����.PrTת�.�����6}��"�?�|� ԍ�������W_��d6勞��1�/`5]�s�i2���	]�Ԉ�9���=�ؼ1�.���k_~��/�M�������-
�ٖV܍�2d�̱<�2'��챾���[�{���
�*AX��7gO�g��}ތ�֣�kjR/7��,�A.�:���6v�)��_?`~���E�f�r�.=��e��M�E�w�	�EjG�ׇf�$��,�X�?����NĖ#��GO	��ZA�Zq�%��Ⱦ�q�U�V���ypN�������a��@[�6��5DSO=�<y�"kũz͢.e`�����ݧ��գ/qq3�.���p�ⅹ��e�+��L�c�_���{y܅^(����d�������Y���1& �ב��2�,��R5^<͍e�]Y��*x~s���V8̅����_Ff��$�q�b�P�� u�j�4S�B�Q/WP����^�l�ݍR�U)�Vz:��8Zo�/]�Ds���L,�D�,Io�T�S (�,�7��=��}��.j:�u�E�*š���glbL�wށ���W� �H������,W
�控w�}ioN�`.��L'tO��2�b�c�t /u�}Ӯ��)@�c�'%I褧2;�$��ZS�3�S�:ӉnCڢ�J�/�r���Q�X@'���^\��`���A+A��N �܀,����{+��T�'�j0�z;#`f⼨T��'Ɔa�UI~����fҳ�R���9�w޿��ϒ��u�4A��
��5ʵe˗��ٓ��u���큁Af"��M���R��+��P�����U-�ץg�E���8�T!v94P��g��O�0��"#1���z�<���g�a��ps��n��8o��l
1�챧S%D���7��4�O��ܦ��bb(5���l�`3��2�c8&�����-�����nK>��H 3��������*~AZI�0�t��}Wtk�馛@Tj\Ƽw��R��E�fB_2L1ߴ^�@3K�&#|��5$�Of��_f��9����2����������v>?8<�J�������޽�,���?�Ț�͛?�p�/��2�ۿ�ۏ>�h5�Y�-^��lڴ���p�������{׮���G�bM�%D[��kx(����*����|��a���G����_�R�sG�����?4�?�R���Lr9e�`ڶ�S�3�F8~���/��I���n�q�Y�W���p�?��ի�z����&�����O�?oǯqq+�c���o~�ŝ;�f�R*�Z��j��?�����-[A����+�رCé!���}�󟟘��.���U)'~�w~GCn݆(]��gv<{�]w֛���Y�T;\O��֭��'?	z.�s�AF��c������0�w~O_���s�z��sL��1�擇�a�T(�-���j�7�
�$���Ū�,���B���$���{y�T������+x��j���FF�W�\i��'N+WZW]�u���#�_o6�w�j�8t�@�`�W�<�w�@��L�'Ǜ��NgY:::��ݼi�k�:6<�0S�tq
/^655y��������ʼ%ˍeR�iˎ���|Js[�c��A3�#k�J>`��y`�f�Al��:3��`���G��'�F�Y��;�S��c,����]��PI�����<95U�(u�v����Jǁ���{u����K1��Z�tE�ө6֜�v<eL$n�r�����k� V2������]4j���fY��?�؎J�^KX�]Q�|��������}�����ر����l�"c���߲1
��&�B�_DZ�����A)o�r*���S�(x+��t��0����*�����Σ5i�U@�u��Y)�˭J����V����ݍf��`�vK	�Kv9�Z�bD����ۘ��hsJ������B�.�:lR��zA��2ӆK��c'�`$U�1�l�iEI
���ʪ�i�A`{�jh�J�Z�c"r�ˁC{���̂yv��h���aw��s��te@���<z4���:�m�T�6�f��*�E�X�����UX��BRv��*"��{2�ә*kVr�(�GM��	�f�����h�Bw���V1�$"R�{��S��]{�Xn3��)��Z�D-^�H'�!���h��������S���K&���Q����QCP��֎%�2��l�@k�U'��3z9i�wD�j���s�%���ߞTͨ9/E�q~�Z��Bc��Au��,�>K�'��7�	��5�O���4AO3�'I���y��J����]��O?��c�)��p�$��:��3���7]w�u��-т_���[�oEb�1w�	���Z�f�L���lH�=��F�.q��`�Ej�y����L�h���@���.oh��ڔ�THr���CV�����;�����Gi���^y��a-}��7s��7[�:뮍�dZ���E�=��`Ak|)f��[o��?��]�v1�B����_��_n߾��c�bf��� \�,�0]F���@Y�m��������?̞���g����������?l���c��Tk6�lԐ��W\q3��㏯^�����n�Tf1�rn���wr����'�����ˢ��S6l���]X�b}�n�w�R�|����6m��?�#�\�Uѿ�H��޸q#��Ê?0�A�`.�\)/?c�_e�&�1ۮ���'�vb�5���$�Vzk&y�ۏ{��=�FW2�tLb���D�!�h��;�izA���M$�bɖ��;���B��ߤ���(������ݐ�X֔��l.\�@^�kR.���+Ȓ|������&���۷�έ_�3�����f�R|�q ߘ��'��w�4���S���BV�a�0��2�9M���쟚8����μ�6�{�7��~�4U�H*��M�J���/q�(���-��ag�7a�Qf�����F)�O�%��9�+��+�;��V���T�3cj�"ss�U�Թc���g�~]$�:�z���
`>\��L8=�#+�j���������Ti�[r6~��sč(� ^�b�@6�R�j����ɱr9q�ML���˷^��B��$��*�qXK���D.DT^X8���TUp�vɁ�_�m�w
ouv45�%���5�>a!�U�y �l�����n��t73v֘�R9%�v���֞i
O�=L�I���h�w6�-q���,Hu�L��b�pc�
6�E�R6��Ra ��Sd��hLa��v'�جd��Q�+i<�r��~���,���2�֙�8�X
�+AT�kx����}Ѝ��s���'��U���`>����g^��D'�y�ņ�m&��f\S4�W�82��D���s_7*�9����h�#s3�c�97���%٘�<"9���:Q6���EI���)d	9�? ������g>c�ᮓ]~�m���c�2LLr�W0A�$}ƌN��������[��T~�W�rӦM6��b��s��m��ŏY5�.iɒF�������\oʀw�[�g�"�~��E�Ї'�	9�����׿��dZdd}�nK������w8���0���q��y�f����2����kF�@J m�0Ø4���P�obb��pY��.w�+��v>�ʾ����d��(�֬=�9z*`/�~�����B�ZM-Y������f/���� H�bexxޖ-[��>t�W.��Z�Î��nػ����O?����>��+f�;v� 6�) K�裏��5��G�J�w~�{��#@�]t_a��(1����_ͣ���o�V�%�F,h�`*{�?5��C}���R�0�(����`���K��\p߳j�fo�����e���R��\F��T���)�Rv�d�SѰ�YUNZs�C1�]VR˝�rŲ��y&����fS��K���:$��l�ժ���:u�	*�m/'S�=R�'J.���&��ћҍ�%R�ڍ���k�KuBJk�1�+����m��� m.WgF<���)Y�����*�1)�J��+V���		3#��Y��a�3#ƪg����RG)o3�'�"�R�5��5�����[j�w�ֱ9C��
��BGw���?j+9���0�X��̉j�|	���#x����MNN����捌�O�81�)涕J�c�(��e��lS܌�R�QGF�e^P1�
"㕖?�ӕ�r��[��Y#��z=dŬkS1��pa���?�J�_@�B�����`\�Pk'�6ɶ���03OA3Fۍ�Q�;O��&�m._C�?:{�����|�#�'(��E��SP���f��H�c=B�?N�m���t i������صz���hP7[�maF���+9�9.���y�eDn��3.��%���D"AF^v�����f�a�s>S�}㴲�Z�<��obY������&_T7Y�je�9����
�3p�|>?<;�����^�es��VFR�n�H����y��S��Yt9����Z]�&S�0�}�	�]+O����c)��H  ��IDAT��Bt��@��"�\���.R��p�ž
 �~��$z�R��7̅rA�.��5�5@mn)���Z�f��:&\������w���P�h�Gз�A!�w�}��UW]�i�2��b�؊w?��2���K/�����K�o*�?*u�x�Lѕh�m)}vN[�S�d&����,W��&Z�y�U�P��u�|.�Ӝ�<�q�u׽���gH��m�O�W����mrbs�ꫯfN�x�	��I�v��mUw~�;��5w&\��"����2�7^�}�w!��ꫯ�D.+dZ4������pOѯ �ܾ};Sm�_�q́d8��s�e?p����Q�{���f��`�Ͽ��#�l8�\i�R�����<�������[na���d����?�яX;o^v�eL`�{;q�;<|��ף�o��o�PM��O��'�]_�E����_��W^ݷo��/���t�1𧑑ydr�����^|�ŏ>��#	ϒ_l[g�0B�:����k�KH1;���իY�#��VԸ��s�Ź����O��#/v��WL�QIm+~U�,k*�� �y(!'����c=wڴ��Z�ٛ
	[M�����e`F0\ǜ׳|����gV���+�"��+�=z���TX��>3��8O���>�498���h�#f%ԓ�L1S3c�d$�yX��-�:Rf]����m!���;���l�Tu�(�ˑ@_�mL��D��������a�C��A8 �
�P�td]mt�V�pw������n��V�/Uj;t�p)
��O��9A�,%�"��/WI����6/8ȝ��$�J�5�����9T2������6�j��NWy������g��S)��V���Pj�� ���,d�y���L���V3���T��N��\+ntt�)� �;c�6�bXa)��rlPPK=R@o���������k��Ok9Â�@�]]ݫW��i��/r7$�zn�	���	Sg�u�kZ��y�ĝs��V������fFTG����y@)Zap�BJX�����٬M��(+��?3X�řg��/i#�}b1����=���Q�6�Tr�9�����=v,�ϖ���2�"3�[��)գ��<42~T���]D��[9�K��$��Hs�%evhf-�d�.�M�q������"St-�ˋ���&ӘYS�Eނ|9��d�gh�ڳ����i�Mɢ%�D�4=*9���wT���n�����
i�FI�f��5���l5c��7l؀�@�X��l����aT7ٺ�R����kxp�Jl�B�5��lx�����Km�)���QI��ʻ>; ��6-F�R����A~L&;͌o+�,�wS�y��s�狎ʊf �F�BD���l۶��k�e��z�)k9���kg���&���_����>�Q�cD��9�V�ڵ�ZNV���c��FiKG���}�2GǑ�zA�l�ls�z{z�-wGh��D�/>�Y��~ಚX-"��+@K���Y,V3Ō�w!
e��Z�Q�B�����d3�Sz_��˗/e#	n������٩�E/�S �g�!t�$oq�����O|�x_�;<y+)L�0n��?�s�����_�W�%�W����q��r��_6�w�i�L��?%��k'��������[��l&� �U^vc��{��g-�X�d��j���c-4���E�y����Vk�w$�۴Ap���<�3V�Sbd���U����tm���W4?1=�P�\mr*9~����^N�6<�	�Þ5�� ��v[ک��i�ͺ�iϘ��A�-!��rIK5g�I�$\��-Z9������ĉ�)�]�g��Wh�����&-�L":nS�b:Qx�Z�}r����ӌ�BdU�Fk��=ɽ*;7ö�ȸ���\�tdͲCD��*�a1K�.�J������\��b���`~_� ��e#� �����;��r�^,+�ַ�ž]�n�=����7�2�CX��'���A9�q��YG����S�2�:����z
�t�+�m��l4~��,O$3���Z�~���t/Z%3��
���D�q����	�Z�4��j�b�0��	/Z�'�q�g0�hM�<���+���[$���y����.�t�h��'��'N݀�H��O؎������U�n���s:}�F��x(>��ۄ�aP�?ODɋِ�[���=��ԥlQ��JU��ZŬ�V!<�4��[	np�� ַ�ew��L�E�~uYYe���9*QK��n��E1elDo��v
��`�sA�o|M>$^|�l+����B�j�� s?��X��m[6o�5�-��b���H�%�<a&#E�l�l�A�H��R3cN���9R�+tL�3�@�iꮉ��.��#��f5�
R&����"_6CE����=��<Okl��QŵsA�'�b5
�=J����n"ὰ�N����z�����`��{��!�A��{o����c���Z�vF[��2��4 ���]��A;��!�i���hv���ۖM	�r�ʕ���1�I�ꋰ'�&�j6B��P�I�G���[��f@<6�u�L��wߝJ���Q.�fa�ݻWӎ��S�~�[��>��s��)���/����{��ǋpp~�W~��w%.ٕ+�,Y�(�cz�u�%����xq��#�.K*���:��}�16<��.䋦xz"̀�-~��-1e*F6����+w��"�:z,�Q)h2�I�D:9�u�~�;�y衇L�*e�'�֯�[�:4�'{��aϟ��������k֜�я~�~����{�c���9��8�%�(��E�*D7���Z����W�e�;v��M+�.�d�=�����\�+�8�u�n����Z
�
���s:$�����u�9�;e
�u0\̋'���{�@��"A%/�-%�~���'_Kbgf29������5�k9yO_��2����Nܙ���#X��.�Ȥ[]�R��3-���x*U�N[�l�{���p�V+�����#K&B��{�'6m٬R  1��j�|��P�j�������(����\?��Q���� ��=EDBX���ގ��>,�v��>����t�D簣�'����a����3WLN�*�MV�ڴ����8�,��1���Q�;El�����uՌ�\`��ѧ�̇BŗSgW�J�h��n\^̸����b��y�����ڤ�����]�e9g������'��:������L)P|�U��B��eK�ƨE�ѹ����%���g�yLE� mA>�,c̜̬ԠGd�B�<v'��ty(Z|߾D	|N��`��SʦM��J��]�9~RoiW��og�A���L�� $,1&�`�����||y�.LY&������^��1��s�$!���vա�qՃ���ƶ��z%P�R�7o(�����'�az��E�Ώ�l�:>5�?4h+�:�T�@'��g��w�N9�KQl���Q�ӈ�����-l���5�*5��p������1��==�:����\FL�|��h��k�.�'�]���F^ԂV����Or%�+�~���B]�jլg���eKW �K2��#�/�g�oć��5�iH]���]ޗ*�������}������W\���O�vkQ�)Lc�����c�=v����H�6�-��w������(���9���I�%sADi�&��^�L�8����o1�F�Q��E��>9�è"{��g�g��$q'jjf�d5^+ɨ�Q��h)�|�A�������z�w_q���>8A�K/���ͷ$����[��,��7n�*��W�VP���	�BT,��M�ӟal�K姶ok��L��k@�#m��X�u3亣�r�}�qہ���p߾T�����{�6]�����n^��Q�ȓka��+�j��^�pdzf���㱂-P��r���}/�295���5��N*�Ǹ���G��sS����pA�W����mٲ����`���H&\�g9������С��n��f�)w����{��@kR��%�`��,�����ň���lZs@������H-�+/��B �4g4�t��,a+�#D�pm�!Ȕ�y���J� ���0V��ԫ����VWw7ҹfa�� b/E6;*}CbDu�t�ڃF��������5��FUe`D�$���8�PC.�&L���%���.g$筬b�yK�-e���U;��5z2�%��J=y|F<g�i�e�R��x���6�c:�������Hld$g&��+SR쯿��O�Y19l�Q��4�##Ò�4�z�*��Z�G���k�ZM��s���?1>��5�f�G"!�&�z0�=�-��������p�M��z��UjsY�m#'��xˤ���3$+�=��D�J��xN��4�号��U��"��/]��TN�����OI�����$^�2���̀N�D�}U,%�G
��'��_�E�T��h$�Yr걱S����3��B�	�O��dGF��7����M&zOd���@Oߣ���n�<!IN]3�ttk	#�P�e���q�*�ͨ��C5ͫe<�oέ0��s�Ӭ8�;��J�j�S��cZ9�_D�V;�mI��)�C`ڄ.e�=��B��+�]�i=Z$9A�bSb2�r��52�Y3Ug��=��V5zT����(����i�J�9
��p7���{.j�������2!����E���������wW�Z��d��|E/�a��OXܷn�:N��;�_Q�/��Y�ڣ��O#�C���(Y�k
�6wJ@�ein|�XSޑ�Gʰ%����C��6��1�ΰ�;��k�y N%z}�#/�� ľ}�tGq���������~\�̘��v-��S|ʸ�=ʸ�m �nL�գ2/��y.�g��ٴm&�&-D@w^���s%�Q\,.F��0�`���o�o�}T�CU�R&_v�e|q��ͼ�A��￟���n� w{Y��2�R�̪��a��ܹs'��o���,�~�~t�$L����̹"o����Y��_xĭn��v4odDG/�ӕ
�l�t���V�$�ӻt�2`�K/�B�O�]|�Ū�FT�����f�(��^��~���3�ܡ�:��,+;\�|-����z�E{��=��lo�RVľ��FN����1\z&Ӟ�_�X�Q1N�=����5��ؐ�
A�=�?�|˃��3�<c�ߚ5g9r��8{���=e�CA�ЊK�z�Y�ҳ�;�PŚL����<`�J2�#pw`�5S�����HW����ȩ���a��@*-#��^W� ����=�})�I+=#E�V֩��o����r��5���ZtI�˰�gօp+V��K/9p���QQl�����7��G �C)I���[�T4�6�b�<c`' =�$,�&���%�c��y�{<ms#�a4���Й��謘���R�*'��#����&���7���_��G>�6��d!�Zg��rf�	9������~���e`o|�`�<�P(��N��.B- ��Ible����h�9E��âϢ&�h��O�}�o+�d9�}�>�o���~��Yh%�G1U��H�N�d�u���˻:{Z�+V-�C�mߪRIfP�P�ɩ��?,��ؙ
�T�#�J�3ZC���P�5 ����2/˖��x���ݚ&5+�lM��#m��Z(�j�Z����,wv�ڤ%���O�DQT_�h!�M�tT�:*��B��!���6f������lM#��:]�����F�sɋQ��������d`=�}��Π�s��E��J�7A�֒��$�3ӳ��ɱS������
�=�ro;��ƣEO%��Y/0��ήA���YrPBi���y�5z�A4 |���O9X����̐�������D��Q~�%k0Ͽ^x!s�{���HX�@/�c�6#ĮDr";�]q��[�&���"�#w�������a����T��b(mV��u�~.��+x(3�K�����e�x��[E����Yܠ�y���L��#�X,�'�fS��לs��k1�4�����{?RI�@Ht��QDÛ��&Q�G�W�PA@?���2v�[���ѯ��u�]�w�>���m�:�(yOl��bt{�pQ��6���x�����	����Y�ˢ��U)������矿��˷m�a�5{��'��Mh�C"��d�7����/^6��Zy&Ȁ�/[�����a��������7�x#7D@3�����W(��H
�U��Z|��A�z��[��V^���g �ib���o�_Nn?6��#2x����c�J��N�� -����� ���:K���͛��ښ�d����A=|��Z�a}��-���cG�T�f����J���˖WgfK�,YD�^��d��^��G�
R�aLyf�XG��+%g�f9&X_��XP��8=D�X������측�������W�����B����B|3�L�0E���x���sA8�џN��>��S|��؍���tQ�G�����1�˖,��U^�~m��J�f�116Y)u�9k-�}�W׮[���ǉ���m3����<uj<�q�ˊ�K�����K��>q(3e�}-����dY����ZQw%���d�/_v���b�3iL���{�Q�Uw�U��s7+[�-+Lčsծ��J�|jrꌕg��ǎ�����^��͕K��VL�MTg�{^ڳ���K�, ֲ��RgGy85�l�L�2-�V��H̓N�t�2`�z*�Lu��E��IeC�Cɂ=5�B��=�V��4�#�}}�;�s&!�\�bY����W*�ݯ��hhX#��1���dK@�<��c���k�Y�$1��P-��v��?�������b٬�Zo��Ð8a����͜wv2G�bt�td�Q�R]�NK:�bKS-��]Z��Ǥ��+Q���{�Zm�3�4[͟��PZ�@ ���"��L���?ݡ/*B	3��C�F���qbMo3���$:J�`yI�-�R�"� R�l�Z4*V5/��5pf�)V:*�l���6����Yc>A��`�uD���J�I��Tɑ�E�j���Z�Jrm�[�T��3>�6�|w������FX�	��\ˈӸ>e�w$�hb-z�k_���jk	-x�����4�8c}.�1|��1�P�dS�;)C�T3��Ox��=�9�%����rʃ�p��^+�����n1?�UMf������ �.e3<��*j�y�aks�4S�@�������yĬ����Iβ�-�F2�'/
�QL?ngg��R0��E4�XkS�'�Ʊ�y_�4\��h�3�[����`R�M�"��	�Ц�.����ɯp�?��?�zVZ�a�'y���U�H�mI&��0�m��m��կ26])�䮻��q��������y/��b)U9��Zٮօ9u�*c@��s�=G��*��>�(�
�b� ���2H�����z~���,�.[��y����^{�u����w�q�e�]V	����/Y!��fC[l��/}��{�մ(G�""+j�ƍ����3�<���F�A-�BdDS�+K�B�Ƭ5��MiB� ��"��z�M*U�C(O�U�(�</����Y[�=��0����X�@�>rA�5Q͊�bH;w�Bi1�z,\�+�}�ml`]��.�L��Pi�P=t"`��[Y9h��Mi-41W�X��@V7�0���I�J[�N�v�(��w�JG���*i��G8��șm^��f�,���
_7}�3���r��U�5��������R3{�?�믾v`ժ�H�j4����P�"W��S����9IQc��id*Г'S�4C�f�����̞�*q�c$��������F�HqXZC��'_>i��<��a��#;���	y���&4���a��{� m;l�1C^YσF���"�1�ҢԬ�p̿�m����*d��BiX;$��E�H]�͜���)J�aN�-��b���}�s^xی�b;�?��m۞�iE��S�����>�)���L��
eX9cnr����_���?��c+pNWgro)�O�z�փ&�j֚�?GY������<���U�.�R���5�F�� *�g��F��z�mP�t�;�r&��Jm�i�Z��#��ƴ��M�Q���irrN�C�:6�V���-Z<==i��={��ی^���aO�En=����8KQ��J���f#�/6�i�<�J�,��H�bZ�՗�g�)�0;o^OW�d-��N(-y��{�
N�3w�&���Y�����׊��ŨmqQ�t1�e�\bU�W�c�y�0!|����`e<����Gr�ʋ�Ri�����-^�(�͛�b��Cp�<��:��4d��W�1�D�8�|�e��W�(Ȝ	�1�&�2r��2q�w�����-+q��iv�w���P�wЋ��)7�Ġ��N'�\�Y6�1cgP5{����Qz�v��Ni�9ڑ������z��Hɕ���m���i������A_��j�O�$;&@�c��>�1V
�d]ge�d?HL���m��˓�}���Fvx:�'1^F"W�Q��s�)�\?�z�!��w�wAE%�4;~�v��#G_xᅳ׮a��I$/���L.�`� b���������Tx��H$�2���h�뮽���2��1$����i��9J�Uՙ��6�����1�	�S"���;w޼a�ѣeP��c�Gw-�/���;���5�\����W�������?�O�<�p!�
LU�7^<;;}��^X����0cLu����FG+劇7�)��{�.0ߩS'w�z�� ��\C3;���m_�WMycQs�M�zI��c[~f#V���f��2�<]b�I��Ī�`��Nt��"�о�`C���X���X��D3L\K����ߌ~.�TH�Ɏգ�SF)pt�ʲk^����3K5-�L��ޘ��r��G:x���#�v_c����O����I�q���)|yo���)*0:t��z��ɱ�Jy�|����/�$7��f�+�tZ�4?���-�Ǐ�U��Q)B�-*DS�Bc��������L�h+V�NMΎ��H�g�:t�hGg�"&�'�,P�0�l�����V#]�ԉ��=F锱`u���� 1��nJ�v�L�^�z�973p�a�V�0�t8�'�kE��V��G�[�~+ƌ৊�h)�as�z��!o���J�Ń>�i��Y�=�oT׮M-�c��t�M�b���%ܸI������'�GԊY;��63B�z��T�m/q�R,:��ј�)s�i���Uaf���)�Yj�Ȓ'
md�}��j�#8��-6�s
�u��+V-+%F���w�x*&���wn�ܾ����p�x�ǅ#�"��ױ�p�6!BGt���XQ�e�[�RR7~��^:��5w*�xz)��D*b��jۃj-%�\Hg����Ɉx8Ê��5�J��Ua��V��q.Z���O�3�C� �����X���xbJv��n���5s��2�i��/oT0,�ߔ�y�]wu��|z��%��ٲF˲���_��C�*�		ܗ䟼"!�� 	��n�@��`0�<a[�eY�dM�<�<���3��]�s�F�n�K�>��޿����黨���*�BQ]��KU�@�*�9Z�Ga�@6i�n%༲,��yɪARž¹�wI��Y�)g!'0�̥ԋ����
���f�1OZ����LA�,�q�$j��L�#�	7���9�2�%8S-wʍ�xi�V�d��&ǭ���8�ǖ�̕�ҫ�)g��kHųN�M-�;v����������3�Ow:{�@�Mz� Q�뮻�y����q�h]��$�N�y����^�x֝�(p	��_�~�S�N9rD2��;�$��
�9zuuY�J'��~]@XJo������6[2)$X��^��}0Jmy��7��={���Wt��KVu�a��Ā4T-Э�_�*d��]��fx?��z�A+��-[�YX��o��o񻓑�?�?BT�`�fI�b���u}��'�)4�׊�X	&3�0f�*�w�N*c����z}&"�q�ɉeE:���D��#K�+�����n)���N$�6�g�c��PG}�>8n	���OTBf��̀d�U�w����Y%�9������	3�6�^_��r���{�t+�q�K5�Bfo2: }$v����pA#���2��{�I� C�Ơ$B ��D��e>?�L������^��zz���e5-5�T���\j)�d���+��,�|% �}��	O5@���.L�7�5��XठIz0Q�#��W���n��6���#�,����}�ц���j-Ҩ<ha��v<���q����g�Z�����J�����*�?V�	��\}S�x�
����J��Lb�J�����qO��M��/kJ������$����$�=�N��Ç���d[~�_���ϟ��Z�ޞ�@�%�JT�
�MQ��W�j�4TR�Z�����9ڋū|��N�8�8�O�����q�������y�W�DP5�u��Z=�ô�:>Z0����/Y�D�25=65=A��ŋ�i��L[���4gsvbA*�S�m뜒r�u{%@���4y�aa!�2�V4)��L�b^QT'�C��A�(�5[s���g&��ZL��s|hNHܱ�\&[�4��g�7]yk)5 ]��/A��(2e/�J�@���	g9�.�TB'������e"�D��C����<Ȯ (I�Y�V����l�(K����I�?u�t�I����^�B�9��t�0�P"NB1�T�ۑam�{�v���U �<}d�<_j���xƏ���e+��a(�����qiA|��f�W��[�}OqS��▫:]�,�~P�S���c���'ߑ���޺l�2��w��-%$q�i�&������N�,yD=D`���%���ijj�kli=w��+����SMA����K��F���/?���)��	�A�u\_ܟ�0�J��u���x�ǎ--�Ȯ���p�|Gg��3�N�Ow<A�Ȼ���;�Ԕ�V���O�B� �n%Wn	�h
b����)p�/R
cw���`�dq5z�g�}V�Uwۿ�Nu6��G%�B'�Lf:ڍ�A7Ѱ5E�.@!��KL�^�?0>h�u�nHq��㧢,�HP�
�Ryꩧ��:��������..�!mh�\�2䝤W���t4u���4���,��C��CK��K��暮�K�����=k��ζ�t:�oM:?�t� �Ν;u��z뭲u=n�3C1a�@�w�]S�M�֪���Ʀ��zM2��_�%�����/�`� �d���Gm���g�#y�N;��~]�����Z��_�����v�����$/��Bq�O�S �.��=Z�W�Щ�$"x5�S��CC#�SX/B��5]�Mg�|�����Fb>��i����kw�����k6n���	h���̞��,s����Lc3ZW���6j���9Ǯ&D������B�? %���������W�����8��7p^nv�/�6Y�!2W0{���tN-�O��tg�V�BLgS��Y�6�K%d;dJ��GI�SٙG�5D�P��%RGP�����N?NPd��àT�k�bY�F���d���?�	��?��?~��}˖-�x�{]�0���~��|pp ��p�?������^�bY�b��W�b�
����%�Q��p�3��5�QP�O����D��S��3�Z������㤑�,���L#���7[�.���¦|��9kh_�7�T��.H.Z�YT�X�_K%�[r9�$Ѹ���q�.�ć��N��seR`,3��Ps�jE	���/���d]��-2��З��H��ə$��/
#�X"��/*Rji�2"}\�9��1i#�vĪ���i��3�T�ј��c9_�7��;_k5�C�O΢��Öii�+V�����Yo����a����G74֫R������"@_��h۶m� �)��S�V�?;�[(�i���d������N�,�K��
��H�Ձ��p���a�ë�؄���i!�S�-�/�8ڧf�	D���a�5 1�O�����O����}��r%x.���	����Oig�&�����*ӻ"e��av�d��m[I�!�-�lu�.�k_�ڗ��%r`�\�G<�H=��p��K�����A�.�H�y�߻��n����{�9LL����Z�Sd!:��;%I�K;�����Z�޶����3�ui��ӝp�4��۷Oo����8�,J�<�q��%�W_}U���I�k����E�4H͛��O�>�G�G�@U��h�n�����}�7o�<�Z�ޅSmK�>�n|�d�jY5����'�x�G/����B����U��{�%T�akf�Dҟ|�I��`����Ѷ��k�:��o1��k�-����/�r�p+R �i��(�dL�N�[�i�4cٕ&�S�6�����Cӥ������
zZ�9����º<S�p�^VRN�E���^���7d����K��L$N7?uꔬD��E�CK@�c�����&A�YbC�<�s�y���	��dg��)��X	s
����G ebj���W�GK�|Cf���� LI_��D3I5�,@��t��Ȟ!EiC�q1
�R�)���n<q�ė��e��F��2(�� %�"M���Ss��bȌ��Gk9�s�ޢ�l���J����v����{�j�z�M����#Ƶ�ZꮮNx	B���W����&� �P0��eI���Vs^�j�^�jzz��]��v���,��ڵ��7C����K�����\.���*C��������
�ɐa���à�@ Xհc��jqа�I/�}��c�U�E"<��M1v�X�A�d��V�1D*�ծ2�Q�Y�?㗟�o����#�5��J����	+��~z֖-���G��Z+�<�$G��k��
Nn^r��rȀJ�.�Z	Rj��6���ٳg�h͡n�k�.��q�����
?�˱hA��eapH���p��M��NL�����l��Ͱ��]��Ue&Ӡ�i���ѭ�!~G��Җ���uBt�
�Y6k�^<��%�m�>ѫa���J@�k`:� ��*N{��h��s�xz�x�_����z	ӤQ�v:+v��N�DɊ3�wŐ�i�q�f��:_n}Ji��i	Bjf$�>�a�? �P2�/�7�G4�;e�A�ȑC�@����J��!� a[1lkA3H:���<���n��^�ߓ�Σe�� �R� �i�9�Ǝ68b�1�-m�r[3��iT��f6����<��ux��Fx�ԩ&��II���XF�T#���+�Xy��y��Gw~��4�w����i~������g�y&�c��$�Ms"����}����ڨ�8���i�~:�Ȧ��ɡ�|��7� �S�/U�������.��Uv@������w���;�t! �C��K�֜_�[��ֳ���$��_Is�ǈId�C�>�^�f���6)y�lE�doo�3Z�rS'��=ƪ��j���C��@ ��ݻu����u;�ˎz뭷@ZQ�H����GɫsP�뮻4c���2)8�'-M3���M����
];��K����m�>��O^SU>�9�|��ݛ7o�ifd�D3�~��
�Ђw�W"�+ޛ�c.UGf:M��c5��L��"3�4�h��`���i�Pj}��ԄC��WӨXa%$��I�B��+���=��������ެ����є�m�w��໦��%�;$�~jnVV�Z�o��c��믵r)ba ˒�冑F��;�j��c!��.��.p}@>6�^�ߨ�y�-���_�̀����l"�$�R�ň@�}�P��P���c��M���)� ��3�OL2���s�Eҁ#䗢Sp��9�U�m<�m�,J�(؈rW�+�����v�K�(� ��<yzݺ����'����_��MK�]�a�:�M�/����w�d���' �%"�y�jE�9B�߫a#�HU�p�;)t���>I�&z��*�UL}ǃ���F#�4j�b��T�_��╽d��1�l�:e��:f��JxJi��=�(/��#�`����-8���W��퉁�&cp���!&���wz�-.p&W�ց5g�ђ��`Kb_FB�Ig?�:����� ���i��1S�打�;�APג����m�2����
G�Gx�4T�~}"Ŭ�20��HR������+ta����8J�L�v��K"����	��I����DC�Q��ИIe�Ԫ$����D�d�#&ܓ���݈�t,N ��Z�Y�A�PN��B`%}ƍ�%���p� �v��lH��!���R�=���kM����*��a��F�n�]rv����
c?���B�a$]�y�'&Ɛ�xRɣ2"��|&��z#��6[���Y���� /��{LJ�_�������Ą`�e�X�R�H�n߾]��믿���֨�Mi_����j�Νt�Е��{���!��H�l�m۶}���&�6��̢ŋME�j[�l������೪����D�7I��.���)�ĩ	�f��[���H�&��O~�~��$�mnf��k!��Hs�����w�8q��W_��~�u4󚱿�����j'x���Vm͚�7�|3�#��z�tlB�(��n����H`����z"���&�--;v��{yߋzJg��]�;wέ����_o�N��!����!i���h�_����۶�[t�����dR�t�5Q��򊹵g���x���BLK3�#��O�X�V�������ڱZm9j_���Lq�����ƶ�/�LWj3�_\��H���S�B}1>T('�
�={nz��UO׊S�Bj�Dd0����J���	\RQ!\��&�pL�V��E��|	�q|�hI8��3�F��ק�:{�~��tb|
�l���֮i�^X -�����H�@�EZ�9=� �jm�&v�n�x K��׀�-���ЫIt#��[���,���>'��|r�66B�LS����ut�!!(����Y�Kz6��h,Yb��T�C�a��'h2�x�ͦ=��'f*A����۽��P�8q�&�7;G3�߿xhhtpph��E��w���&9&��r劽{��x֭_C�D������ӕ�[>�����U��\		2p�D�~g���}^	��0����F�H��S�XY�bѤ dTq�0@o��0�����I�ُ	�0��ZP�M$�jfY����t��O4�҉r-��ef'':[[�Z�ϝ9�����,�/�\Z�rE"45477����Dgƣa�ZP3
�DP,�[ۚQ���Ah��C�.��Թ��w�����cv�:�X�j�-�ZT�X����hbm�F�՘��g`nf
���u���[������3S����Z���9�x��;���
��z�\X���a���ѣG.됟?����]�gf�+7�l�r^�/���tӻd���JT�{Nm	S	�g�~�:�M��E�.��܂�lk�&(:%����؄�?$G�ם���s��J��j����LN��a-S).>�T�B{{�Nfٴɱ���]LF��x��ΧJJ,v<{��ZDx�]8�Q�2a�^����Pި?I����F\ DN��i4�&�&�^$ҭ-�S�SX]�{������Ih��i�3��Q�f��O0:~g�kq�1+0���\a!o��1�A"O4e�6�rͦC��>�\��M,������_|�׾��/�����e(	�_(.Y�l`�ʁ����k`��c�g$ʉ��E40�� �KI$^F�4VݪU�46�v�޸��~Z�o�r���M7�dܤK�R��ܕ�����+Hd�2��3�/��]�:s���l���+7W����[;�˗���,[��߾}�s�������}�╇��������4����&�D:7��okk��Y���ci��X��ɓg���K_���r��͚��/X�����G��x>�?��r���ߒ�����]��R977/�&yW����ֶ�����n�+�9����}�^�tE2J�K"΅��O~�W���k�l��c�ӂ,#MM͚�'Nn�z��n��~zrr"��U���/���[:uk�ׯߨQ=��ǅ�N�8Ӑn����y�ʆ��������W��X]�6���LKS����w{���;��u��ۅ�RY�\mjh*�s��d�lOWw�T�l�e��:���c�u�͕fL��/�}�{u��Dr����a7�:�s�\�dR��aK-�m59x��V�7 i*:zqaGt!.m��By�W�\��21PP��Fr�m��� ��w�}$�r��3�:U�F��l�"�aλ��_c��z�K��r�"�#��YڴwIk��n.]�=�mڪ?I�^4:����x�)��ռ�T�K�.�w��R�o� ]8:OV
��s3����������5>6�ꊀ��wv���-�����*�2�d�X��#iO?5���8uw�]�-%_z���ZLsv�������m�=�BC�)��^���h�@���p��T��JcSft�p��Y�W�hEwk�D�ƾv�7�yO%4Hpz��75R��9o��eÙ��P�d�L�
Ӫ��HyB����C�s�d����ruQw�Ղ\r����U˭B67s���ɐ�Hr��<��)̢���1j'�%M֜����{
9���K���l��R-�bt�/���;3��ԐL��mV)��f��X"㥁���B�8/J�L�Q`QK&P��ӗʤ'�dfk�z�@�jM���_�d�\�%kzN>���	�Ea�(M�&�u�	J�T[�m�A���.���h�	�'����M
���3�@3@T�$v�oRO9�/Ľ��<D��@�Vx�.9Q��D�'��Q2�������I�m���Q,M��0Ҙ"�M��P�ܼB2lkH�ҭ�2	�[���	���?.���mm��B7�.TWP��>s	X���Ro��q�AN���G��"��ڦM���V݊ނ�-p�k�2Ð�S���D'��l7��N�c�h�4`9�%t�<�EbW�@=S�HtI[��'\ǘe�.��)���H�X�6��
ڱ DH^R6�@��x�&��P���n|.Tb�ޖ�]P����!�8ig�#��bI`(գ�R��P��{j��N�E�H���?�a�<Θ��I�cE��_1ju�!�k.	o��t$��N���:1�F��kn��y����r1
t�r���K��O�d&b=4������3�#������x(ɛ$ϚRvK��[u���챓'O�4� ��&�I�JRsp��7kA59/���SO=s�w}�ע�%��|P �*wZĨ*��5<��f�iz�i�����ug65.�?� ��~���l��<��)�"}JkmeSS�$�z	L��W�Ӥ�0JK �lnn^K/	���9k�Tأ�����߹����D����{)zCCV&�v�$3A�W_}U�!Qs��H.i ��լ
�I��z�O��߭�?~\3O�!R���j��G.��"XCI���m	]�=��)J��8=�^�=�*��J��lc��IJ(ڄ,}�F����B��CmQ���
}AfP9?��0��,_�lѢ�F|�(;�}�&��:C����o���$=kn-���r-��t����'$g��2h���ErZ0;�\ͧ�u��_��_�1���q��iz���l޼YO�Va���K���(Н;w�]���^����˗@��]�7@Mo��%�)Y�P eB{R��i���������MH���e�u	���|
��N�C��/)y!~;6*�U
�CT��΂Yr�)bhQ�	Q��X�Ĉ��4�1N(I#���ԝ5ǯel~��V���th�a�RX�OBYFk`�M�3�I^�|�S]m�S=ٍ\����T:I6tGW{CSc�SG����G܃unFɤx�A9�!*�%Zo7\�����GƑ�H� !Kv~c� J���P������+/�g��K����H>���s��\<l���E��Ņ�غ��N&Y��PXp[��ײ�Ke˂ҍ��e�󅨑�A^�hR�y�a+��u�$uO���41<u�f&L)�1+XO;�}�W�<E�:YT��dHM�?	^y�#�~�
��J���i!�Q�i!W���8��RBDW�2-�F%�
��
�P�#�UE�C���].%�TM�	�Ơy�T"��&�ɂA
�m˵���}�d��U--M����%1���m�#Āu~�}��=�'ZV)~�ha�����2xd�'VG�iaF��]�#�hw��$��a�ͭ��欂��Ŋ~._2�2>Q�R(�:dr4����c�
G�<$좳b&����+gfmᤁ�u�5zܶm�|c~~N7#i�X,x�R+e���zŻ��z�����L��2�pdt(�x��;�C/�{����a	�ի��]t�W6l^"8n�Ls��C=d���\�3>P����ڽ��D�����[X�֚i�b�tCA"�5����IJ��g���9=,�%P��%쩐-�2��������RǄlH
4!����,p���1>>�wnp����ޡ�.���}H#�lp�֭Ҧ�^"!X���P�}H�B������B���qu7p�B�2, �x1�&�A�#�Z�v1�tUM��$ʡE/;u��h��0�y �&MK��ŗ�WQ�R�����<�U�~G��V��򊃰>�4d�m�ssQtE�X֑�ΰ�1)��#!U�&َW��%Q`�>	�z�)��e�$�)�O�>:>FH�쯁N���Q��	
:��}Qw>t���m��FF���'����_Ϣ��n�Y%�-��ӧ���%@>�{���c�I��/��S�4����^��-��P����[3G�Hݫ��LM�"���r�a���Ĕm���`����B�딌&�DBtJP�; ���n�[�~�wV�v*a/&R�q���;NԻy)�Bs�:xO��;�R�UO �R����G�H�LmĜ�Gm5Z!p�n5S��-��o`�uo��\���]����g�?�]�7�M-j'���q�m�ZJ�l�rm�;��bQ��j��W �B�q�#\�� k"."�-� ,�C�A���� �T$��<5�����R���	(D�&��,���3B`hGP���z�br�@��T�1ME:U�X��Qh������k8��$`�� p���� /|U=�#p�v�^�fNh<A�����)^���Y}�;A�a�����#[�[�:GLC�7	��D�8iN�6�!`�g�$7�J!-	�$� �B�2B��.�]������� #�P(��WG��J���6��	�K� ��^�<�%pGl�Pf6$�SΨ�*D-�������DLG,�R*�39Ѥ���"�$ѹj�*�?Mf�j7��o�C�lx�N�8Q�^�*�,�?^�R��t��Ё/�_��Pi�G�i��]����u#�����f�&����#G���@�r�-�=�R��V}�ђ��9�f��b^���ڡ���Y�cn���ϼ}J�g�&˚ji��Nl����:�,cR��-ۻ)���!����
rQ���gvvF�5V�O;	R�_��G�
R�.��ׇdk��?���64�R��gϞիW?�KO��ƣ}�ӫݭP����߿s���{�����~ )��!�G��*I��g��v����nh�j�4�	u�>͘��O<�O��O�A�a�|!/U�e˖�}�{�m[4�7�xc�S���ױ�Ǆ�~�a@.r���Do+�g��ړ�E��Iw�{��o��/�*a�5%�p�p��s�)�==���Ji3J��zqm��۷�}���F�]#�6#�S��܃�9ӽV0�����#hkC��%, �	�i� ���΂��p��E�y����:C�5�vI(<Д�g�9� 4 Kq+D}�̨�zÝ����*�[�^q�2�q��y��u�5�\#,+!��J��h��W��_wze�R���9v���_�k7�%�R���#ځt��M6lX'�~��ۚ.=�TiS�lK-�b�u�@&���Ma�'���Gx�[�[s���dў8k��j�/���i�GqR2d`��l�T ļ��
	 ;��R��y@���~(t�t=+�GސX��{ң����3�� I�
i.�ba82r����)�����zշ�m�W�I�Lf���ٸi����a�Ë��A��)$x��#���C����֗\�m�$ H�2g��3I���,����o�C�P6���yK%`~r�76Պ���&Б�Wt�-����t����ӢƁ�؈��w'�C:Iw{���'S��q���'f�m�L���Gl�ZX����}�"�k9��R�s��1�wİ�,*X{��Ƣ��./|QxGܳ��F�P�;Lcİx|Z�j�|l�dU]hCBaI�h��ۧ;\��j�M	sSO@� "?��L�6�J��F2�P2��@N�%4:�ت1�@_��S�ȐӖЊP�Ixw2���`NBj�5�%.s6Z������]a���?u��O>I	3q��uw�}��՚���=z��-��uىUu�l�UK2�����|߻߻u�v�EK�kn��%pgu$���ᗪ��Bp�lV��"ǜ�f�>���7�Aӑ����ɭX�J���ze�>
�f�-Fn��g|b��g�����]\���SO=����<��#�|h]tP�;v󭷼�;'�g���q3 ���@��uF+m�@O{{������o�/iP�3F.�$i<4$�������m۶E�F��ݱg�FRuRHx�5`r�,'����_��_��_i�\�-{�9� ��bQ��[o�a�"	�:3ޤN��y$��\IΔQ�j��Mن��\�Hwj�.]�Ԍ�K.����:22��z={���pll��w��a���ң��۷o5����誅�[�[���>�ч.]$�]� �hiպl��/~����݋��.h������^p{�DR�V-gnIZզ�W�dsJ�I���U;�>e�p�W(�vr��t�W_}Ub�f���\�֫��v[U��q8!C
�311i}P��d�h��V�]��ӭi�T���43^�3ʩ�B��L��AgJC"�˺�x�Kc ���
eLS��x�Q祋��B�k��H�8����� ���?��pik	p��$W�̮]�t-�fC[��k�%/��WY皖�Y�na}��О��
��9��`��#[��#�����A�׌�E+���_w_�Y�@�'�bLy��1c�K�3'�'i�-��6���)j�p���B���>�M��H��ؙ������1w�H�Zh�\���>�p۲If��O�89>1<<(�:*��ɆT�"P<�c^LPhA
�`E�Ŷ�)���1ݪ�Zȟ�-�2C����t�T��m!�ȎdӃ`$t���@Q]	3Y�I�q�!A��oIE��G.J�g;R_�C��M,� d��&W�mX%$!#l��֜\���F�|��+b��>�7C;k�!��,wv/H�@�ѡ"`
�yR��%CPw�[YWRD�ϱ\�^QB�U�t�@��/9E~�"8��'��RC�j���.��]�5:��T���r�q&��k��Z-�\��D�z
���}��T~q���g���=WBˤ�%O�l���~�+fI��4ۆtB��<��ɂDؚ�: z�c`��,�6������O�&��W�W���:" ��8gΞ"{2�-���8p� Q����%Լ�*>|8_�'�N�i��U�%�X
j��^�1������%��4��r�w>����~��S�55�E��ɮ.k�1�֎F%B�������u�]�bKӘK�ٸ0N�<�o�X�ʙ9S�n�{�)F���@����e��C7���6�u����{�'?�	�1��|��a���^�I��	��d�T?yN��}C�p��h�����Y�d���:$RO|�B�z�D�+���_�l߾]����R궚U͉�D&c]�_�ы���SC��[n��3Ɇb�y�t`�E�EM���?����W L�AzM���������|��;r��p�����P�Ni����]��S�N�������.&]I`���D����e5uF��]��n�O�z����ΰ��)�ɇ5�1@N�߅�H��%�u��GuZ4s�O� �tm�� �)�JSϞ��ZY��Lc���!Zs�B��հ;/.�4
8`�#���� �DVvK��̀^�v����:"�z�5kV�зz��t�!�4z����)���/���KlB蜢7�N�A�Jݷ���Gq�2i�\�k�>��#O�eb	�V�ְN�q��F�!ǂS6�Ӊ?��#^��SQ(3r�pgt:J�?�m3��h�LA^�ϩ��̱�'���z[*CZ��5f�vHs�~Ca�:��:}<�,*H��c��7�X��,ԛb�����g���k�.5�j!��5��?���J�\�U��&�0���k�>O���薄�
�����l�7g#�.���O�N�н~G�FWʎP�b��F҉�bf�����e@�D��#ɉ���DWR�eS��xt>o	��.��^�d�aj��p�R��g��M����Y�������TJ�M�
}�ɻy@~���B�ˮ"�!vgl!�M�қ5���l)�?#�'��G�r��57 �p�a<Žw8� ��*�V�8�3�'�$��0��r�ģ���՜������ $I�i��΅}�0���`�f,�H#ŐlM5T��Z��A�4eԁ���x���d��CvKҫVϞ=�w�^�a�;I'zz-�.���+�a���϶��!���������[Ȕ�}�Y_���n��,⯂׊�>������S�.Xb] 4��	?�i� ��kh=���7�l��h򞞮7��H�?S0���K�D��h���c���/����ظ�9�,I�R-�E$p
E-k=Q(䅺v������ӳi��g��o�3#�r�r'�M�[�����;��۷aÆ�zH(SpMK�����ٳ�[m��ڵ������hB��Z�;w��JJ5�D�C�¦ȃSy���oݺU�WXD�Dkq��!P�ƍ�35''O��	)P`�^Ҙq�\w�֑�	�]�a�ƅ����o�߿_�N_��N��M\s͆7���־c�͹������f��vә3�����a[xv�M����?��#z�7�|S�L;�;	7�0���7��wfQ�㙳g��q�_��_cW n�.�A�g�\9y2���;ke5�Q��-�z�D8��Ƞ*1��\a�`Mi�T��4�ǅL/��U̡��|�5ɤ��=�Io��ׂJ2���܃��<2�8Z ���]�V��"5���1�	gϞ��dN�G`���:����'ՠ���Df���R�w�?,g�5j��DR��89�$증Z��|�_ڴ��Q4Û�|���`nΊ�Fծ�Y �N�9X[�������P2�_�54fpp���E�5���ݼ�Zp�D'�(Q��1v;;]���y=S<$�#2ƳHRB�P*a` $g��W�;D*m�NAS�DF��\�kP������%Ja� �\�m�u%^�w2�Y)��x�������Ɔ�r��2��k����!3�9��!�ʉ����$��O6z�/��pa�XH���{�>�l�[��{wXO��4GH}������X풚w'��=E��I-N�N4u��v�`6ȃ�R����аH���P��ؼ��������0|�ϖvu�19�Jv��a��G�]G[��|����8���:E��q��$�U/H���D�S���]L{�k�!R����6���oB����`GX*t1�U�X{Q�VV�XC2,F��o����k��P�'�诘t��@�IjD�.1���W��
��֭ˇ\Ǭ`�U�T��0g�Æ���AɄÖ_��B�R!��k�݋ۉE<򋇘l<�[��R����U&�M�H}啗�N�gۯ\ ���f����_���b��<����;2�ug@��)o�.T�7�Z��L���hOv�dy�Yo����=��o��6ضm�R�f��r:85̆� ���%XO���S��3㭷�J�hy�|�����ϝ�|������h���.��)���/���H��&)���U����~���aG�1.�K�F6�����f��~�#d�"���R�P��覆&�$��D-�{b"%$���2#B��Ⱦ��ܽ{7�9�n�+h<�M�6���KG�4cӼ	fif�~��^��_GG�P������_�켃V��L��_������H�8u.FF���;�;"7I�寽����������]��]�;.^��ҥ�¸�+�s�9�D�LgG�?�a����>��J��օ�ӝ�W�j�0Q�-Gks�����͆
�S����0�CX�����W�;�V|�Ν�oZhd�n��9!�"jv���2���dT�^����f�x�B�zG�@qAgފ��睧�#M�Ǒ�g�B�PGRs�bc$�	�#��(��7jO'�|�ưE]L`���M/K&�0��?��T���I�lp�s�F�41	��9�3@�B�R8����y�Ř��l�P�]�~��������C��C�
���B����J{s'�1?�'�&�@A  �vc$o#�Ǧ������ja ���������Al�mw�Πz����+��c��C�6i'c/�3��ѣP�[0��Pl:aOjU�
&果��:��ށ>��YY��ca�u� $��c�Rœ�=-�,����	"�D�lύ�M��N��J;�9s���76��u�	Epf��ZKx��d���ڐ8�rq�]��P�sϦ�`A��^k8A�2�'�)%.�۴ɨ�c�Fy
� J��u&��{tn�7�Nґ�srQ<���Hj������*??�ТJ��h���W�k5���uI'�@�e�/_a0<��0�?zS��M-q2��ࡡB.�RHi�/��:e�L��5�$���a�Տ�p�Zl_����҇��"�����\��%lAd�cI	'�Q��g�g�I8cĩ�똊`�O���2�,4D|�Y��-��E��FN�^Y��"���^�3J���S������.������,I-Q�ދ/|����_�������NX������������H�	� n�;�s׮]lэ7J�0x��wh`��DH���<%�S���$ �3�)E�\$�eѩ��/����Œ�(���w܆GY�PR���G���Gj�y��=�裏j>���������g�y��ge.5;fez;���~��~���C�L���A�A8���������?�s��ъ�ٲe�~y��S��{z��l���E T�J�mܸ^{��0�nF�rU	�ƬO4`��|�A��� W#t>�K�J5��a#]��xʿ��oQ����Bz�_I!3�EJ���RB56��=���Mw�q�ΎfIo�s�u>�W�:|��3��bQϙ�|z�/~�B�7�|3����	Q(@��.]�zr �H��ZS���1*��V᧞��7�<��МxAC�p�p���ŝCr�俤�'\��."� Љ>�z{yͪ����p͒I�$F�tIWgTڴ�|���x����ʕ�B޲(��buZ��+SS"�"ܢ+�s`�>O&�^�܆;��#�z�իW^�l��ޔb5���(�'����ר闌[5��E�P��}����۷�`piA{.���нJ[�Z{M簽����Ys�Q�j�u�X��0>-`�ĬQi̚s-�&A�Ś�L��m�͉c��C��/�.Q#�e5?�a��D�p-F���s�������y~nN�B*$�SgrIV�7!��`�yqA<2���L=��=8�p�G�?
Alc<�?E+b�T+A!_o���'O�k���2<eE��3SV�f�3����XKk�����\�T�B�I�wĠ���Jر<Pw�v�������]���'Y�@$U�!O����� �H� �h�"�3�qn� �;Q�{�۔��1bb���+��FI��T� ����{ 3���pt6�ݩyϓ^�����4�\A�Q'�!�`�`�L��K"�8$�&�GJ&~l�HBE���,N -�E��<[��c¿����h�A����$��&qr��JZ�����6�d�SVxV��`�ƻ�@q�!���Tnp����~
�j��*=��gMu�׮]�q�/. ;O�MJ_����v�<��)%�}O�	�X{���(������)� �Ap&����A��-�m6l*��c��7Aa~8�ށ�J^���L�,%w��_�������w� *.	";v����T�������|�^ R	����2�x1��'ĸi��oQu/X�˄��z�vm{�z�	S���MR�/�q-|
�	&�S�%�����!����+I0ЕB-6�J�����w�>�쳚�O~�a�g��:t��a'Դo���mÞ�*�(�g��5�}��56�d�-�jV[���?�����J�!g��sxi� ����ʼ[Gx�1���MN�������������ֿ��i`Z�ӧOl!|u�{�"�UpΗ,�-F�8>�-�WM��ͤ&������׾�e:w�p��@WJ�jҴ�����}��8|�M��f�&Ұ@'��s�iZ�� �ts�	�4=���;v���護ު��m��hM��y����/��
y�AA�ǎ��;.Om�Y��f#�,(���6�B�M���#���"0x\(OF�㟫�.�A�Ѣb�y�W��L9��Eﰌ=�ֺ�K�-�rSx�%�$�GDB���	������l�����_�Ս[�CG���XQ�K/�D�)���� $���5?x(��&s�iN�	 �����Q����\�n7�t��`��nif$��G��I ׅ�v��X��%:������>��BAt�x^P����
C@�8G0�H�Ł��J�Jưc�Ss�.!&����?�T����a�p^��Jx7K�>�4<Ϟ�iWL۔z�g*i~�X<���k��Q�r���EƢ�c�}����~ڇ���m��+�\ LNOЊ[���a	�vg�I��"�i;���@�ā0�Q����y`����G/��(Y� �q�pN�k`�|�r�c\�Fp# �����y�fb	e��뮻N��я~DV 
���&���ĉ�&�%��1n�Z�65�-�Ʋ�_�3?9a�Gvp�K�S���T��Ε��#5.����5�Tvzjօ]&�J����	���ҽ���B�K"v���}b�`����F� �=���5
(_�!Z��s<DJ���x�-�"�#ո`t�s�6R*��ƛ^n�
��D�:����G�&��|f�G(@� P2��>���;�1$�XY,~�5R~��N���a��ss��>��С�/������?�x�B��4�K��K�VQ���?��PF�V^:U|�;ޡ�<y2��%�,}�Ձ+�J�ot&lPMY��;+K����|)���j�x�rnv^��ϥQH�i]k	�%�}��u=99�.���=28X,q�������?���k�W*agtN�,i��[�^{�m7OMN� %�7~�r���^�rx�:ɦ���!(�zKy��x���ޫ�I|ͪ�{(��c�� ڻt��S�k���Y-����_}�U�r��;w���+����XM�D�hHWWwssl;� V��u� ��9��fsW�Ă� �]w�ktt\�C�f��t:�ʫ%_�nusKc[{�/>�����^N����F
\��$��0$ 
��˫?�O���ۚ7]��#ޚtH<��ɥK�8�Z��[�� Uq`��di���V��]pC��70���z:9�T;�zΔ��������P�/�V͍��0����1��fh2ͫ^R
٪y�`Ii��z)�U��n�_��`49�}*%�3N֪	tG�u���Z�n��ȕ��u"���(��� ��.���=B�$.ONN9��L�&�I�hGuj��{!�5��v�y�G�B�i�b6YM B�T�-���Z�;2��#�\Ě�m�W&��0�0��K���H�;q���+EL�䬷u�t3�/��JXs��TH��)[Q��7BQr���IK��ۙ�.�(P-��'b��!Q�ŵ�1)h}'T+���4�a�׍�NsA�X���c����-�Ӡ���v��-�=,RSY-��<��6�<MB�@�����gc�\f�!q�)qP�bQ8��-���`�x�m޿X�s",_C��K���h�.��XB�MI'Phrzq6����/�Zc�1V���4.&>^���P6��)�A�����/8�.����%�4JiG>�#��¾$!��?�0o��erL (�1�ފ���(z�2O+a+!��x4��}Z"�]4�j�h�g>�?����Z`k5d�!��P�ɐk�FgrH�(���P;G����.Г7��u���)֨*jl�ѧ�" ��I �{��ٳ`G�Y��+�gǎ�<��ѣG��F;�2��,�$C5�HRik��s�%:���{�{��ޕ+W�K��W���${R�ǂp���������k��i' AJ(8U��'R�uͱc�֭[�z�:A����>��ۣ_�#��$�Y�=6l ���h8���ޘ��K�8�)�Ӵ�b��WM�R��~������y��)�HR3���庅��9-NDn�#�aЛ�Kh<��iH$��7�����!g��mظ��CU
	�4B-z�s�=�{�nA��_]`%�=�X53�4	5�xXZP�$ /0�4Q}}�aC�|�rsC�l-�3��L<���~p��o߾�ر�D������u��_���W�����q�3�c�>S�������[>���n޼9������=��Eչ��o����@����Ӹh55QB�ps�J�S���E�R4�4Τ	��'�(� l����n������l�,��4!�6771r3���2��N>s������_����6N�+�Z��z����$���D+>�d�;͡@�^��sk��]���&�q�>���"�HJ�RB�$�CE0	RHҰ [�ɾ���r�!��N�58nz�!�Xq�E�@9���&t��n	~"4c���&;*��D�|�hU��IM��'�;���n��s޿�b�i �E�*�-T�R0t+����<Q��,FFƢ������÷��"�մr�p"' E$��W��V�~�*k�'Qi!�V�$=�+���N���d�ό�4�k���Ii6|f�2Pm(��u��M_(�<��sͺ���m�Holq-��.\�v����>���&���������9���r4u�V�S�B����%rUC�@@ ��9Q!�"I��IC�c���A���+%�e�G�5,0�C��ȏ� ���׀ղ�N�Q���ҪnՐ��r� �W,��������V^$��'B�_�J�޲���SS��%>hNw�7h�5'{>2�l�(4�@!-�J����iH����"�������lkz�� ��G�S}�X�Rc�|(^A?U��Y�� �d�E�!����+1�@F����8�o=��;���L��%�ԯ�٪o������l�!W�۶m�Z"<*�C�Nv��Fr@�.I�(��]�z���&'&�)��d�\)��j	��}v6��k�����}�cd��G��ڻw��I��,i"�E=+�ϵ��1�h~d��H�%}����˭�bBpm�h���;k|im[��<yx�]��Y=��ߡ������/�KZa,�=����!O���r�&���IX�w�wkN�������'�������<�E���ɜ�{��- t�'>��/��$v#�ZP�� 
�h��������u�&����>��O
^��?�v����[5/�ѹ8�|2��!��������L�������qO=F��RW�N(�����M���������_�*:��'����W�\ibbLb@#ٳg��e@'�ɐ4�t3Ȩ�(�P{-��t�M���v���k��v�u�Ar��[�	��PQB��mIr��TP��W ��S��D�Xտ:���؝zS���u��s���$4 Uz�������6ģ)�N{{�XA���j��	���jJ''�pG�=oAWw�������?��D8�z#�[�"��<�\ˤu��&�D\�|yddtӦ��BI�.�
I�Ǌ�$�5x,�F������I�$�?���?i64�T�PuA�"�a�:��E-H�˄4X�B���b!P�Q�~�^��$���HJ���/X���*��bm���#1��J!E�s
��z�[�ڵ�YS�D�'�P����#�I|
����t��X,o@����.�/0#J^��QwR��vb��EQ����._�������R	!Z�#-h���+�Z�^�`)c��F��(�\�?��?��N4����ό�<.[��7�H-o�I��˖v�+{�܀�%S�>��ca5��媳X��A0��|�}�o�8��=|�]�I2.��O^ŤOB�10�HA��Ǐv�M)om���7����p6� 2�h�"�@L��G�u���
WI�
܏���0K�F޴�{Xo<�xhi��h[	��7"�	�Nc�C
��n.;��0��<]��A��Q��$!	�r+=�]IF(�`/ܫL�	��&B�k�C��(]�:��&	�+�z�"����9�1u�	3`��.��j0G/�H��&��`<������^���hzq�,]EQҜ��u��o�ypp��[̱��%�e�n��R��I�p�Zť]��7n�x��B��i�3�4iaҲz�W^yE�D�����t�M7�$-BF�^u�C3]��	�H�h{$��Ls�6��/��j$���"��9��kB�-����ѣF����~��������Μ>���'�P�Ş.�ɘ�A����v�������СCV�������/�O$��^���Eh��ms��$tQ�Rп\�ܲM� t�WR���$�̱w�� {��@����2$M�G4���~��~A� :�l�����V��Lp?���#V(\�p!�Br^J%;,C�� 2iN%+ͦ���s���۩��}��8n��^%�{���mZA��Z,Ͷ���ů��B�C��+��tuvg�Ơ�)��Z�-�*0z뭷�>}Z�	����cc�HjL�ޓ>����ݷx����g͓�tL]�� ��ƍ�ҧ}���0ѡo�����B�EgdD�O�	�;�c�R�B�$D�A��/^&���#�$����J����KA'�%�G;�8dښ紓e��)�H�\ժ��0#�� �4��$fa�χl��;�����B�A\kx�Pv��}H��q>�@�@�])���bi���AFɸz)l���Ř`=Tc�՜2��VRЂ���a��rYP^;k]�)K��������5W�Er}�x=�X5Lkn�}�#��wG�W�M)�Z��h��y'�g��C5�!gΣ�e���w�kat�B�{gn����U�,�C锃�c���t�Z�2.*���2L�A��g�<�?�g²�vke�#�<3�����h~�I&ՠ	��N�(`B.PT8�g
V#�ͺ#��');�Q�d�7�#�y�
ᅁD���4�U�P�Y��U�'��hk���<JQ׿��%A!�{��Uݝ�0�(;>�Yo�˞���j&�x��Q�@d�ɨUOeܲIr��53����?������aci't��	I�1c!�^@*�W58��C&�#o�����fm@sJ��D�<:5���Z��'%���Q�@c�4:�;�Q<���#�g59�~�@=+�G�))�*NSaG��������m���u�i�V���İ0tC��'ƒ[�du��l6����\��`A�8m!Lb&�B؃KKq��;�Wqh�+='�d�R&~��Ih�[ZM�JzJ� >���M�ť_o��������R��5X&ը{J��[1�S�}:�:��ۺu��Ա�GW�Y#9�;��>r�*	��IA#���a���_���裏?~|̩^�C��^N5;���~��W�����w�ޭY����¦w�u� z��QD�N����d�*`���[��[	�#�;k�t6c�7y�r�l����K5T]���=K-	�@�z�7hg
�i`\2�R!��֢����w�}��}��'i��N�5� D��hǑ�u��[zYm!��V���v���=��c�=���>��3�F�H3)=������<��������O�'�	���m���r�-=���	�	MYtԄ��#�l�0^r�((��B��;q��т}:�۷o�Z�;w.鬳���t���kk��K%������ռ�kժ�ӳt?�x��b������ØC�h�WgsU�����?��>!�h�\?V
�%؞>1A����s���[-��ӪeO��e_-Րmli�p�2�I���	\�X���NN�(u���E
Pso|"8�24;�w�D.i$�Pϕ�Jy�$��Y'*�Tc�P��c�;P賰����,����߸�[����!�k��BV>M3�h�I�h�c1(�y�����BB�۔����lCkO7R�p��r���jaw)�Y�7�LS.V�D����A�(���Ia���d�XK�+��#��5Ŭ�2H{,�ʤZ9p����y�*h��U��R�޹|U��E�)���g��!}̓��Ջ5Ɉ�n���!�ìd��%��8�(�c	���(26������x�p2,�c�s��"��W��3�Z��� �e�I�a���%���3Sǡ��,
Y��e���Fli/Tv��IΞ�ӕ�6h�� 6�giS��i���N��Z@W$�һ̤�HKn�j���P<n��
6Ɋ�VtK��. �K��_,Ă3Y��t��-r�����%�4�Rlq�q���n��T��]���M��k�PTQ�V0�7�~\��I"ݼ�k0�#�#[���=�1����|~:�P��v��2�=�a�?�q�x@�Qr1���*��H��&ܫA�����?�n��ΑA2�����4���m��v�w��}~��~Lg�0�`���xȀ��H����L"M�uX�����߰~��vV�C��/�H`���҄\�9�R��4J���^��N�����5��H������m2?q��AS���;XC�%hB���?��=�!@�Θ[�j��Ç�聍����g�yF7��JN�|y`@��'�]�M���M���L���Lo��B�#�>fv�h��K/��y;r��"�cǎI�x*[�����F<v㍻5�O=��VDZ#����t���1�EM#�_Ƙ0;G��5�\�q�Va�ΝC4*�����33SdXd$x�m���z<~7�gϞ֖v('�{�9��`��}�D��}�#@ R����W�B�;J�+{@�
G#��6*�L�!$|4�4*
5M��� ��8��c�͛��G�M�&A�o��gki0�H����`�����;�i �I6oںf��3g���6* ҂�];y�J�6��q�V)�T���F�h�� !Ӿŵ��.Zԫ'����I�`N�*T�i��X�Py�Y�r���PLU/�a2a��kq���r���^?�f޲D���^��>P>/+1E�0�ăBr�d��@�j�;"h�t0���7Q+�������eSgD�b��b�����g$��`�zS��	���6 �s"��Tr�Q:��H��II�jn�����A�H��!p@T�Z=�j\	�,��׆'��=��s��h�8�1���D�7�iq�����?KU�YI�^��]��d�	ڥ�م��T�L���j�GF�T��@W��_[C:����ӽda��А	��L����B��y���X�D�����i,�	B2��^)��������_1v�3��;+�74l��W,3Kb��f�*scV%�s�S9v<Q�'�J���M͙��n)͙Y�`���Q�\�ăX�R�[0WJ�X\�+���n�h˕�!��nmn�"���9I��M񗊳�)[%d�s��T������������>�������g*��d�d|xh�ah���<�]���T�Z)A���d���S�
�KT��g�!
�ń���u�����􋾖�]�v�3)�ӹ�lG{�y��c��(j��{-p)�_��/��2�3&n������cx�p1�ܔd�5����><do���X�阥ai���)�Ni>m�WGjo& �AZ
w4���B�p�D-�v���%����kn��vAl6gx]+�GX�H�0�`��d�Eqy"��f�m׼���`��]�l�v������R7��M�檵�t$�����bian~��+6ñx�Z+Λ����_+B[ԕ�8'��f��߿D����$x=z���n&[�����R�g�_�۽{7�Ρѱ��a)��Vc�2k�6��I"�ܞI���3#"�)v����I��CI�D��B�OG��c.�[d�h�n��V���#2b0�ْ�����e}�zV�X�oɬ:/�R��Cod��Zwg��ɪ�x���Mޛ\b]R��{�y�Wt�[n���`���~z�=���>��o�1��Z�f��\\ЮK�͍142Q,K���K	þ��kgN��mK�Tȗ^zq�ԭv���LOG�ʥ����R�<51662D��|n���P.k^��,�]�bhd�̹���[���������-[��O��K�yG�3g_��^P�;t��eп��ѣ��h2u^$�6lؠW��p^��������o������7ޘ��lmm.�K��L{������|���;p��̒�ə���Xl�g�2�(Ztn�'��n޶x�R͆6�M7������_|Q���#�H |��nn��)�ݱǵ{�ZJkS[*�߸Ѣ�CC�_�>т�^�z�Y3�N�W���떳��ܵk܄��ʕ���k�wj��9s�>װ��}nA��҅�7����Mp������lڴI_����;w\'�;jt���R�I_�p��і���	D��?qX�jI�UR��N.[�D��!%�q�J��H���X:��U�%���5c����$f��H�����%��d��>���jG�]�_�=4�?�2쉉[�9�йj���MMw���t�&'p�eK��V�.Ц��!��;�h���'O��=����띜p
��r�D�RlZh����!M����u��['O�H�R�W.����6���%KڼeV�]M�39<p�S3/	����;!���'>HfK����X�9����*�z���)c���"}l��B%��ܜ��7�7 �F�8��A�����M�F����,	1W��L��Q�U&�llk��#0>�:7j=�։����%�[-���J�R��}�W�X�y�R�.[�ߚ�M���dK�UH,�M;�F��R*ꡲ%����l:���L�7��E�HA�j5���E�`s�U��4����E���x7bA����<m<�A��d$%A_��E���5wT<F0�����ѐ6ע.��Yt���j�0|�m�5�=U��2�����<DsY�0�J�W���bhl���Vok�d�:h �IO�?ӥ+a���ˤS�V��8TL����<�[�C��i�zn��-����wtvv��Á\��|��qe��<wnn!E��"�
7U}+���9ಏs3�Q�Y_��H��<�s�a�@��ơ�:1ӊ��S6���K�Jw���Y��  X��v_�aH��I�d6�9 o&�|�&^l"�ɤsc�"J0�<�V��n�ǐ	�3KU`��� ��95�T��d��F��"�rň�7 M95E��	�4Vb���"+H��һ.��뮻t�fiQ���iBt���?���y�-d�k���P"U�q�E�K=.x=B0�P��{�H��8��X�~=�u�(-2�SanJ��R՘Ț�u�֡<���(�7��{��($~J*���O�f@O��y�!��~X�G�JC���T�@��Ԁ�+��$|P�<:r���Y�B`�s��^Ѐ��r*��P6XN������m5ZV&G�߿��W�V{I�C�@��uj�h�)ӃDC�GㄪT�\�+k���mu4�������u4�:y�ǔĝV���_נ�\% �D��G��Y����6O"��C-Yb�ǫa_��_�Zz�_������TfI��ܹ��p6�\�[ˡ�<e���ܜF�>��4<�O�>��>XӮ�5�8��v��B����a�&�*P8N��GOhɂ�'�#�u(��`B�H婦��<}���I�щ�ME)�F�k
����&��sMyr�[�Q�E�-Y�8����R ��Q��W�Zf|���� �Q�:w�N���!��1x�Y�V%˙p�&P���m�H���J��k���)`P���v-�źç>����{����&\��[iW�ȋϩ��D�tOb����VD]�}i�Ȣ���&,x��q����ω(��%s��!�A	'� ���e�  AP�=� ]��lV���,�+�&���4b��1�_(����j�2����=�$��4M!Sg�� A�h�=�{g�f;����·��V�&�$H��B�ԡ\�{����Gd�7V���p���sޣ}��P�	ŉD��l�jk���=֭����}�a�	�W�	��M�%o��ם�`SDU�_;���u�Yt��-dyeIi/%޶�r����Ui���H�������xUVM4��ۗ2!��V�����֫?4[�b*����#�,
Ĳ<����=��1`��Z2 ��Bp������&:�,��>��I$�4uz��m���h�����*M7���������G�y�Y��fS�͍�&��h�)ܽX7菙�?��R.~�����[��@ɭ�$���@�� l������P�����A�-5iꤹ�a���=s��@��PA�0�*���e &7�'�bRs<�F�Yqa�89k��O�e~�1G������Ϣ�߬�ir>�h������v�lbQ����A�,���E�{�� 8�4��N� m@CU����G�B��֦�H���ݝ�hN��5 ���,A���/��CJ�!>x�G;�97�?��1�CÔ/���;�5/W;�.D��T��_��NP�=�~�y�6%���v�B�5���޸s��o�[Q�x���Ջ�]�ј�ğ�xL����� ����g^r]sI�4�W��6���*�c�8#�=AT �Ľ�X��J�@���8��􄽽'Ϟ�������k7n�nK�L�>>��_�q����w��O�<ӡ�������V;�s�6K�]�7��4E�֬e��C8������?��Vw�[�^Z�ba�v�5������?�񳘆��l�F�����̻�����ۇ?����HC�'�
�X1ޢ��[�`�Mٹ��p�4 ]#ɇ��[�:�l���јFR�t�\��O<�ZL�ox�1�t:���k7�omo�}�k�4��E1����w��܋G|���զ|�/MA�CO�G�7�!
�2+/^���{�o����p���T{�曇o���Dg��{�����|>{�@�����y�޽��Ϟ=��"���s�Nʯ~���Z�^���J=Ц��֛ڠ���d6���F1/��Բ���(�+��u/*<�dkg��46Eg�
�蟨�߰@g��^����ˏ���~�X':V�����ݽ]��E m^��c��$��|�>�'�<�:48��ѩ�����H���T�Ľ@7�7�� gD��	5x-J��ۧ�馿�]�a�Eh<C����N������ٳd�R���
�D������g `M���W4c���Ar���^��M '�yI��Y�C	+I�qVIG��s�ֿ�˯�h�#����7C�t���`pt�M�)�Eh�I8�fn_�F��eARO/*�L}�Q�D��OYjaQU�~�@'�3<�x�����$��v>��*	�md6��C���`�f��W)���G��b���$l֍����.·&4��ٗe�Օg�Y��ؘH�����Ko�Y�`|��]T�d�Ef����uH(VNy�%^݊��`�R����������nM4e*�C�z���A�<�_h��eu`��0S\�/K؄.�~���8 V�TH��b�x�B%�g�X��h�}3�VTB;XB�P_ 5�R�U�΄�I�Vc�M�)���IT�%� 0��ǘ���v�e!���tAb����'���)���O�I�Q��G	�b�)f�x�{D�(�� ���ݓt��S��T(B�S�?Y%�O�?�`C5G�$Q�X����'t2` ur�E@= - �(��Ҏ����'I��񳘳B�5[�jK�$F"sc�j�<2K�n��g������h'~�(�j�lh�XixX��X�f�g��.`�R��W�I+b9�
�V�r�L,�>��DT�],12i"��ǺF�Q���ӟ�T�C�g��P�������w4<�jL	�{���/�����UԎ8��/�������Ǻ��얒m�#�;*����;ꇢ؏>��K�X�P�VDX�V̲\���~MS+CCL��Wi����f�X~��_��'?����O�^њ��T�p��#�Is�lӲ|��τᨕZxӧ�߼q�o��o�����'��O�N����3�����/j��~�EF�j�D���5���/MD�������N���D�jO5;�?y��JC1g�hbV��k/��.:����4������kK�˥�����_��_��|�	U�1�L�gVU����d�qQ��V��bu�*@�V � /�Va6̄SI]*�M�o�\4�@T�8z�F����?�޽���C}B�Y�2߮fA .a�F�T`~#<�)�ZU��L��#:Q"w[(��$������Xi\���#��۠(Mcs}f�����-NrsV.�1�L�U��U�꣒ [����Q�x0�sC��-M���Ճ��3F�2��Z(r
�U�@3ņ
��g�w�V<sӓ����wBl	�F�pN)���&逡�<�n�OC]  Fnn���J�$���M?��Wf�P?�H6!%��w[����&ª4ԇ3 �Y畆�K|�4�AOx�\u�����J���Z$�����������ѿ����W� ��������1��n���\We�I��a��nQ��iwggs���g�� �D�8��x�?菨���tr>�~��|f���|��i��!F����Y}KH����;�q�@G��O��@]�`���h�ѻ�v#�D�#���N5�a=ZF��7�-���g)oƣ~�{ ���\�C�Z߹dss둨���^Hv�$j�zYָN������!n>�#k�X�N�V�eo� bխ,�fj>ӫW�R�_#�t��Ltg�41�����x�	�3n�q|�M���Z�k����`�o��D���3KŪ�bϪYjw��/>���xNG��M�%9n���v��N���Rw�~o(5;f�Z�͍eJ���#-K�2�s�����>�\W��Ue�����o��o��X����������[9�BF���+�%����Y���j�}�ݲrzb��Z�؏6��D$q��rr|Fa�ɼ��g�����bL�yj��*
qnX����G5=��hkۺ�^�z�lbf�w��.����z�}��W_}}~bp\��h���*��OL�k�b�7��Ҕ���M�>f l�m���&�����?%�����h��걖H��?u�H����Z�������|Úi�/_zQ�I��{�,�Ώ�E�y��P�����+�+�Z}[U�Lf���t�Z�ß��/~�O��{A�+׮��wew����GO��eU}��ߓ�������������ÿ�ɇ�������ß�P�n��Ck`����H�2a�����/��@wj�j�}���y��l͢�葄���h��]g�hY�.��;qj/,���\t���bjhvg��Ç���{��-�����+{e� ��*��x~��m�W?���&�_>���{�Y���j[����f���������#/D���o4ȝ���ӳ�/�/��v�:v&�!/bw:YAW	���TN�/'G!Z"�l ����%�o�\��T�2d�����ww�ܸ����W��>?�����o���Aa�/���Xŧ�~��to��[7E��ǧ'泾{�H69'r?wO�nb�g'xB�	y�ԝ{��wO2-��7�Te��� 2�q�ZC0����0a��F��X�}@/͚�4(x�[7%Vtg�9(��	��`/�jQ��E��x꾷�ͼ`��{?4����w�7�� ��>����3#aC�pԴu1�Z�x�E�PySv+����A���;�{��	f�+D��f��b�?:r����s�IlD�i;�<��P0+£(���[�X�V1sd��L��� ,#��%.0\�-|����Fӗ�)��K�>:��b�|��m�<�2lU}ݳ�3"��cLc�K\���.�$7�|&s�VFK�u�g���!�����z�&��W �0�������<��|�z�����=���Y��<6f+�gm)g���2U@Q|�l�(%��Ю�AsBbj4�PkG��b'�wN����^w�͈%�{�A���U��X��a�"lo$�0�"��'��H/lf/�x�8^<�S����r�l�ZV�2-�mb?硖:�v�уtt%Pb	_f1��ow%��`Y{ES�3�a�d�нp��=��N���7Q�zѯ��Ѩ|H�1\E������������pVR{�mB��މv�x	.�8r�b��}�Y(��,8�#�"6Bg_:�37���;ư�Z��S
^?L��=~��/���4DB�44��M�k��?{��0��p��3�&^�-û޻�B-�p����'���2$�24��B����ϓ�WzOsKr����������=�x�]*�X��>�K��8�(��VJ��.���w{3K̍ۖA�I��o���n"}۪n�i��(0�G�Gil�Xh䚩n�����?�����7�`��	����������S-�w�������3]��{�Y�ƍ�Z��/��R0�>ym�t��1Vc�X��Q#��l�_���ʾ�vS���-	����4#���{��M�G*���c�e��[;^�ƘO�6m����/)u���%��6�=}��0��[�?����h��mo�%�j@G^5�L)izY
_%DZO�{��!�L@��\��O�Ii0���X���{���W�N����Q��W�ܵ"l�o͔DZ��~KqA�F��UHa���I�OQz���tF����{KvP}c�m/Dq��ɚ��6�`hD�ȆM%hqH5e���h����'x�T?����?/�9DrR�R���=� `:KR
$�6O�x��{�:ȡĺ��_"�����m'��M5�x�TC}x�n+0�?���0��T77�$uv��?b��^�s���[MC�<�{nh�{rr�n��i� @01��0y,�܁S�,+C7?��[`?��B@J���P�W����_II�<�x��Ft��K��\�i�,D�v���Q�ᷦ
v5���;���k�i��i�&���kU��̢@Ҽ2xh�\u�9A��%T�����	�mo�l�.t̄��a9k�	֨������EU�1bhІ)� �`3Cx��I
\3xl���*�"��=Eʱ)U.�� [iܯZb�%�G#Qm��c�F4����M���7��*���!��7�-=@
�pc<���WWn���ԛ�Dۭ���ձ1D�Z����*��������)p֟O&gε��M�?k�%��� ������O��1e{����L�1h8��o�[��Vl�����%��[Vu��'"usg;&%?:��{��s�X�b��#fzs�Zo8����`K����W�3k�C}�kpdJ�~���H{�������gz�V�@^VV�z�*��,T�!���x�	+l�x�A�U��}�rGH��'������j �C���4T�����ׯ_�\�����!$ɱ��+�AmZVֳ���C^�P��`�sa����O�tzdV+b�ž�3�50�Q,���(P�Cr���}%�)��A��7�y���
`}-2Ω�S��\�{�2}d���������ܿbu��ŀ�zieP�fs{�;�wxx"y&�&�!�=h�`1�)5�ټxaX���yW���/~!�HՀ[�nU�L��|��߾z���9�rc��..�����q7 |A�Ѓ���oP�/�M���k��Z��"i �(��;X���,4�r-���������7���b����Ma�S�B޾}K���o�saM��o��wŬ���@SiE���-'g���x�[o��ǝ�{����+7���d���H��<�Ų�ҍs?4�V��K K��a�a����C��+l�2��V[���!_
lEh����o?���8��C	s{G���7w���Zg�x䰿o�#g���_|a`�A������
��}��ܡ;=���G������!1ͨ�ʎ�X�ċ��r���k����t}HaG���E�AOg��I�zbӉ�'ӳ��p89=y�Y�>'J!n"��bz�U���c�_4��,��?�1�Ѽ��5n(3�������Zs\�x?+�vB =��[���o]�ӭ��Oo޺�����z�R�76r�/�M�t6�~����ƹ�Fh�d���Lw��5��7�k�s�|�U�����i����x�	�����;�  p�藢�'Sm�
��.X�eh�����.i��-f}����|����a?m�y�'�?�7+8�5�5ȭuK!$�����1m�":�I��no2���%�p�6���ҏ�%���=?`iU�.	�\�ln�4��(����c�~r`;���S���ptzCb�.�!G������q�,e�z���OW��=�"j�w>!����z��������θ����|l,��{���-Ma1G�����	
7(�vшg̮�G�ǉ7���XRч�-C̖S-FG�c����H�h*�aF"LM/	*O>�(#�K�C�#�:Я�:jX�k������~9&����I"^��%��p@��\i.x�cE�æ�3E�C#��a,Ċ�6�ы��X�������b�O�X!�F�P�}�`��$j
�A'���[$̀(B̽���#��?���|=�s�-���)͊M�����a)�O'~��D�>�裏�2d�l�d�{��b�@#y�╄�S������q���<�>+C����dOq� F��b�(�OϠs
X�������X#�����H?Į,A����R�T�^�C�qx����ۿͽ]w�+bbD� �P��]f$ΎME��oy�����y��jI�Z{:!d����9캛FA
c��G����5�a4@횰�_��_F`54�wh�G����qAQ�m���zC��so���������Z
v
�i4*�#�O9����Coԫ`_d%!j��Ć��_��ԝ��/�R��ѓ��c�SlBVa�s��K{���C=w�_��XP��$nn�O�_��W4f�c�ѣu��(��Pi�,z��q�FȲ���"{͈�h�J��d�(��Q�	�'�
��쿾�c��_z5P��t}�7�I0/:#鞨7z��2y<�\ot+8@��Lh4&�N,h������sL�z��]H���C���F��]!�a���B��_Q����>��O������6K�#�ԢE{�Ĕ:m���P�I[#�zz�G�7�2�FT��&q�b�So����%N�ӟ�������+m��#���J,�$�������im�R{O���9��5���
(6��S(�_S���}A5J%���-7p `jE�"L^*���9�u5��O��v��.���� ��iB����9�Ja
!�.��0�V��k�g]�Y�ux����"��MJ�
E9��yvz�ԥ��V��Y�]��������g�'�f`!o�u_�vEK|x|�%��ܴ� �`�X}�^��aJC���LtcԮc?�D�v�5��3��p�|&u}��5j�&k�^��nm.@�a����ў�)dm5�<�O��f��{7���o�3����m[}�r�@�����ګI��>"�"���6�-�O�����VS�� ���*�Y����^yO��L�����t���{��cָ�cb�mx�K9���NN�8r�H������ϧ���A�0P������XE����Lu�?(�Y'+�-#�06�
��x3��7���D!T�B`F��ʗ/�AnrZ�\�V��J
�G]D�B�!�L�|�]�!B�D�2a8�!p\��V3T`��E��q]T���z�{���k`�M�����d]|���+@T�q`�{��ޢ}��$^�����3�M,�F�M}���_@L0A�ޱ&��d��Uw��m���(C��Euj������j����o��ᢈ����S\̅�`.y苧A���d�,J��ee>f��cK>��s������o�_�qݗ�\�C\A�F��3�"����_c�Q�7gs���-����(��'VY���������/��'Ѫ��O�3�0yϠj�ztLI3��Bᡋ�_��	�:|�����}�{"3�h��zZ�������/��g��?o�.���|���9;;���Ȓd���@�_�e�!�-�19=��mg��x��	��z����z��g�]Ho����ŋ}���S���l�Burv��8�m)�þh�c������ǟjCaf����s�L�aѤ ee��^��5!V�ѵJ:ATo������`������m�=~x�����ypx��`o���B1�v�77uZO7ǣ?}��E��:I7=�H��1��/~�����z��������7�v�j�=��hx�/¾o��Ϟ�@�"��"�tYЎ���;���P/5�/dF�Gb�p�pҽ�w�ܱhW��|~�a�ׯ����ϰJp|Ro]CD��B
_
��Ą���4Z���3�����
2���� �w������{i�S7vJ���-9����?y�ؒ�g3$�tʋ��޲�t�Ŝ"�t4�$��[�JA��]n�{&������e׾|y�����D��"��hi�mV ���)����+�>i���%O�΂�4i*�wtxD����b����o?��8URG�U=	��x��:Lh�=O(��Ed�U�ո^*�"�<��bg�F�͍�h��,ƥ9�B}�?��-:D���+�N�"n\�	i����������~��ߟ��~d�_!9��h�
?}�Gh EbJ]`�#^�B�����"@+�u%eN�aj(����
!����1��~�[��D�j��A��ۨ�|�ᚠ
\�,��Gu��$H���7�����t\�8=��%Kp�M0�[&=�p%���R#�	#��V1ܔDY�)x�'�II����v����װ`��É��6�y1��!ņc������O�ҽЕ�H}���I��
_�L�s0�z9�����$��� bn�#s����=��T��Q�ƅ:�Z�.<��#������%��@�bn<Fk�%rQ���:X@�a6�b'�'H2����" Kz���y":��X�Zt��~�������T�E�H�uH��}��Є��*Ŷք�a����0�"4ƍa����dbauck�)t�#��@lb�E�b��TO' H��&����aX)6��y4x�g�F�������w��/�l�����c��v��7^C������7����;M�>��w?𪳖���s1m�Eym韄Oݼi����-4�Û>$��׿�5u������G}����_��~��?~����!t�-���{ｧY��_ռ��,�q�4�a�ާ��%C�"^���5M�PV��'�$������,qKT8B1�{�1mJ�b��&jMd��L�Ц�x�<1�d��j�6�zId��"�1�)}2��j�8�v�0�L<\��5�ύG����]#؜hXu7쎸��Ŋ�&-�h<�������W��D S"��4�k�(w!p��:d��$���h��qfa.�K�-|�"�*48Bq�A�X��$����'>�b��GJ�"��4H�|����"DN�٥+Q�Q��� �p"A�ƺ7�+�̫����63JBm3�y���0"dV�@�@L7nDӇ��p�j����ӟ>����?2��޾��b�.���=%��BU��,���~�<�M�C �DУ)f�V4�%I�M{�K�!Ioޟ�ck�y��A�5��b��M���Avr��W����������v6��W���O���^>n��͞�r���DSHN9�9P6��re�p�&$���&��M���ŋ�.s�@��֑ݝ-@+n�M�D �/�5'?`kk�>?&Ϭٹ+�y�Dֺ���[`|�6@��%�:	2������Y���Ȋr^O������a�){�Q���l�~���\13~Z�a����`(Ĝ���jU*Ϭ6A��@�KBn>/���C�E\��ά�C?Mj�.�eM�a���uss��p^;�>5�r����ZzC�cYb�+���V�r��2MrGQ�?�FYS�3��xh�@��{�KcjJbF���-fY�%���)�T����6U߆�)����xc���?ȯ]�2����g\�43�DWh��768'�K�n��uU���X�����^>�T�s�ܞ�S�+]���.��O��}'������)�&��t+̐"��Va�*w�]=���bw��M'V�cg{S���)X@�x"0w׬��yۺfo�44�
�ja����\������H����qr|��D�z����j^f�nf�Mp4�7[&u4}Qn\�2�b̧�{&�����8��}�h�8�3cj�n�`M�^�YSV�Xq	�99<ӛ�t�.�	r��.�CћNW�(s�?99}��k����n�}�*�g'G�X�i'G���	��YT�x8�~�@XW�xoǊˌï>��(�`���pt�ꕤ*O��"_{p�g	t9����H�쳨Q�5������}�
��xf�����\��?��iz����ɱV�`�����Ջ[7��N��Zj�E}��y�j���O�}�����+q��;�؊Y�o�=}���o��'�˿������{�ῳ�9��G?��亄��mD�m�@����7D�h�ض��5�HK{����P�c��k׬O�;�^�x��c�}JlZ��E�ոw��'VK7N�5z�鴓�EPN���:���X�J`I9��ʘa���7�w����u�>=�zpe{{��ٚ�s�&v8���M�g��d>Kww�yf>�gOͧ���$J������s2�6F��Ϲ ���Ç�
����bp�4��]K*�j%�/�+�/�|�cWЊ����E�Q_m��m�e���R�tNN${Ͻ(z���y�`��5T����4�Y��s���2�'a21#��v���J��'�i���k䇇6M�W�?�����^�b1��𑇯iR����+z��5��vp���sD��Y�<��!��Xh^�/��L&I����K��\}ba�z��Hhk���}N�ϯ9�?9mۤ���}J���E�p4FL�W��j��Hш�?�n�m�	�8y0�'�c�5y#���b�@��T�Q�����S�����Ϗ�%k�w6���DS/$�*(K��r���Y�YHX��#e��+0�u�,s\i�h���t�v�X\�,C����F8�(�K�闕�5]���v��{u��� /�7����(2�?~�JŔ*g�i��)ʄ8�{���rvz��mLXՓ�o�������ps��$4�n#�F�z����s�y�"&,j6f��Y�e�Ʈ:4�q��
����$4��j&�"=7��{ �I;w嵅�'��}�!��i���!������`c��[�^3#H0Y�`D�Q��p
��x�>�0_N�����2�������nH �ɚ6�z
1�$�. /)�{l�s�����ъ(��[3������M'X�P��:�-J�����'L,Bi:�R�)u�)�ɉ�y�9|j1$��G��L��\�T�c�q�{�,��a)��'�����&�L��v:9î�"��zl�$����K����+墌%�5k���3q�>�P�v��K�^�(v�DAl��NO�[�?�sU�1P�6s��V}�n�2ڍ�^��]-f�b.V�(�;���ܣ\�лLR�Ϡ���A����5��6��]ξ������	ʽ���  S���� L#@�'j��H=U�\L�*�t��zUj��<@�n~td�Obk`,�g�������?>��C����w�{@�>�Gw89>&���6-��l�%AI%�t Lx���(d1#b�a4T�9�q�L/�_�@J<��xs�2�S��]wm[R�W_}u��}�|څ6�t�&^�d���E�?P!n{��6�������5�e�`-�Z�����~+�4t�H�w�XCI��c��fz��z���@�*�&��K�����|��������;w\�v��1�7��x��(J��v��N�P�i���B�qxJ�qS@.㰪B�e��4r��+���$`��v_' 4vJX"l�Έ�<�J����]$�XĽ�%�U�}�tJq�q�E���k7�Y��J�͠Q�Nߜ��ȕ�j1L�������P�|�uFO�{���	�e�1�|�^Q6K�:[Y[���;�U&���f�KC�5��j���32�14��ߴZ�B�����,�:6X�F�t1�?z����?��ps|�����7�鿭�'ǹ��3��ol�M7�(&)�����4ۛ�(u@�"�n�}������;�oa�A�d�}�Is�bF��mp��C&p%��IP�Ds{;��~4����&� tݽh�P;{���%Mk�K5��I�k����r}7\k����$z�+�ZiQ�"q�F뵫�8\�N��~������H;fy[-��C��}I~��i�i�C-�j2�R 垣y�#���lL �W�e���36??��W���n�)�F"T��r���R���=X`m�q�V�_�!�8�"��� S�PR��67p�v'ȨR/�����[�Te�Ý�p+ി��Q*�h8 n���KEG�ǰ툺�?8�w��b�e
IZW<&4�1]w�v�y#5{�{�S������y�4�J�l��!X*�{�<���p���� @���o���n޼��ߧ&01�� �n߾�e�E`�^�}�lG�v�u��Lʪп�[3�\�n9zs��_�a);��_~�����|���փn{� ��
�;�I�t��w}L�hw�^�����r0��g��3+�"�}c<~�[o�Jӷ��b:�y+-֨���ڲ�w:�fT�6ƣ{w��)�.�v߼���kW�)�����Y����S[����m�n�[��޹m6M�,�r���J[�w�S�qZ:�7�5P����t�o��ƃ�>�
�{�i��9�*�$��y�ٓ��V�Kt�s��1^+����2$�%uj���ܫ,���0n\��J�g����r���v�?;��㡮,�E����R H�p�J�w�w�ȸG�ր1
��h����Y-̳'�k������e����+b�+bZk�螑��iF��u;�R(y_�ŉ���|��A!y���f����b{1��o\s��B�R���S+t2��ݽ}�����I�N�g'�3�YV��c��Χ3]�12;�f��7�2(��*��7��lK|��:4�Z�Fc��f��ejZLiǴ���� �o\&��&�o�VM�h��yj�D�����nn���(�Wtט���U�! ��'��B�����Vz�6t��4A��r}����!Mf��k�16��� �y���!����~9��Ȳ�Ԣ{jz�)�����n{U���XWna	gz�V�{ξ��G�qa� =��q<����uvÑY
���zMzZ�W ��0���WM��p �T�A�(�${���3�fx���V��b�Ef[#ӥ�:q	�>Ǻr�\��l`Mf]lF�&�(�@�^�I�-��S���Y��LxE���\ΌL��9�EipYp��kZ�Y���P���)��`7w�VpP0���V����o�˕�k"�{�����#]�z���tcs<�����|2u�M��y����t���s���J�M�4�{['��Ը#�|z�Q�Y����w�Q<@[�W�Wv�����5Ll4Q�c�q�Ua2?��N����q>% ��V��a� ���b30���Ŋ�2a��}W���������+;	ey��m��Im�`�����H�����"Y�8��Ԭ�^����"Vf}g+�	
�!्�o�������uLq�d}��!��z���\TU7�2�N����O�T�����\bN��:{���"����|ǌ�;rlm������`�x�󗾫_�@4@���B�5�+��LhL��e�8cGICO�۷o����Ãi4��-^����qr�ZJ��Fh+�d�s6-����RО���u�)�"�ӓ	�:}�U��M^G�"L�9�d[��R��(�M�X#�tvnj�ѝ;�5��d������Cp`���x>/h� ��	޸qU!��,�͋���76�Q����Y��z6�m<��\��3A��/~>2�Z���}'�+Zcw����z�eC�<��6 Zmq�ݳ����&S!����k^X�ƕ+�~p�z���[o�%R�e?h�l�����N�ب���bQ8'1�+Ӡ>��lOS;��t.`WXUH?k=��J��1�w�J�V?�^b���)]�z^�A�@	~�8t>�,��kO|."�,Otü�:II�7Z�&R�O�������-����K3&�ݻ��3�7o^�=	�ӱ�rq�d!W�RT,;Ȃ=E���v�ѐ@���iZ������I�]�w`�òX�r�n}ԩ���۴z�F-�jk�y=�o�{r|��@)T���~�32#9	�� Yl%�ܹ�_�@�!n��Ϟ�仌��>n��C�����>�-L���r����L'��#��X�����c�;�}�6ڦ0��ގ%��s)�X��3�AdPicoow�t��0��؆&פ(q]��Z�"��X�)���1��f$ �<�*1�|��N��3%M�̭"U�sm��FK�˛����W����P@}o�v��������S�/��e��\1*��5K���g�"��*�+�� �D(�{�� �͂���ê4ߋv�6?cu��	�-�^ѓ�.�q�f�?�Z58���Ϟ=!���P��h{<"D̖:7��f\"p��^ �N���IB 7�U�į�آu�YXg��yE�ګ��JkOJhE��S�COWĹ�k�V���狉������ɋ8|����F�����z�kt����f�H2+�G|�Z!��!M�l�YS�m �}ߞ����^7���1vK,"���t�e� mЯ�f4/��,�2���:��跶k�-|�@񚝞��E��g�ܜ·�C��l�JY�@1�Joө�`^�u�[�j�n�'��B�E(������K,����f�ͱ��VE%a��|���K�n�m|�,�k}-]!��K��Ƣ?�ZV�D�
D��esD�!*Z���)�� �h#�<7F�r �i����ީ	C17' ?f$a�K3Ҭ\�_����p�x�P�:�q(`�Í>�i:tU�)�Y��o��`7�`q1����^!Q��ɱ��� ja1����]?�Ł�y�.:�;,�Y�ˆ��a�3��&���S�������� q=Yl�8$���3�cw����8/Z;�T�H�>�flL�P]b�uOH)п�|��}���Ɲ�DjSS�ң��f^	]8�e[���3���J�������z��j��f��V�ە�_��M��-pI	��zCa���~���>�x0,轛4(�L��'X�>r����1ƕ��e�/v�z����+ws���s���WG�����>�ۊ1 q���8���@��ٖO���x}�G�����Ӟx�J�Q�mon`5ߊ �Pn0�q�X�|Q�Yڵ����bG=j����}����\o��NOҐ�3�{e-���$�Em�$f�+�ƆP��z�$�7���l�<b��>�-��n�38n~Ծ	�\\fsl�=U1���l��T�X�Y��b�����7oV�l�b{���X�b�cu;�LM�󡔢�1i(��ko�Țd(���G1-�tlv���ֳ��6Q,q�5����4����(���\��Ң���M�p����ٳGn�����3�t�ؓh�1���.Z�c�%�Nψ7|�f���,/�|�k�����ա�k[Pn���cl1��+t�s�H�Z4Ѣ$��k׽ �j�.���b�(Xbt ��R��9�c�):�=���3�"�@B�<u�� �7F�֍ZV�b"�Ύ_���dzS��߸F��U��xh�|�at�iֵҍ��27��,��;�d>sŻ�C®Yv�l
��C�U�L�4��Ζ�ͦ���"hBZ
����ZTGc��N&3����r6���ߋݸz����x1��ˬg�G؁�}�׀I�����>~Ҫ��u��Q��C;&�E*ih����UtQ1%�A(���.��}��wB�yH�I�$'���py�v�w97�H�]��q��S	�	�m���1Am'/��ʶo��#�^9��*n��D���e�3ۮ���	������5��M�ђ��n�qw�!q�=+��`���k0�X4��XNH(�`����C<y����!�]�I<�'�"�崳��\w+���;�46���>!N����Db�z+GI3L�,�4腔�Cs�^^�2r�Pۆ�D�䎛{���`ʯ��p�X��&A���:;?���Ǐ��z����b���2rb���mߒ(W[~E�2E�� ��R��?�~��� j��2R�_�V�h'�������<���tO�ס� )`�Z겯���޽{�	�HU�Ӹnܸ�
Ǣ'BQ$�֡z"���<���������Y�k|x�[�bh����[�ȡ��m�kפݡ=s� i�G#�Uu�L$��k��*���u�-�4��p%F�9�z)��R��.��i%�k�R+Z��g��}go��I���
�[��^o�ç&~T����t��S8��.��b����H��5+~�H�0�<�!�HA�)�΀B�:g
ˍ�t���Z?��n�EaH���L<���w���7S�C:��v�����g��`֩��U�
ɵkHMT *c
�1� ���@��җ ����atÈ	��z��J��y���6 ����皩�̈́�a�N��1�v���C��@�0j�(�ّ*�q�B�z-�F��E=��tN�Q�Z]۬BK�ƫ��C}�rH��0�5�&%7�^�JAw���o�&b��>�`#K��~�
��	o���L��چm�RM����Q���h������D�`Jz��nC 13�'���CSч#�A3����w��T���}Qr��*UF���ۏ�,�d��j�,K�x��������O����c���beƣύw����W/�4��2����]?���'Evc\-N�a���e^3��6��Ά�Zo����,SK9���=.�g�).,B?M2M���	[���s�������]Y6�z�6�¬C�o���&ˠ.����N:�:A{;�,-I��u�-"�9�� �e]E�"J-&;�#��x��ܚ��,���i*DY�������K��"ć��4��Q;�~dlƌ�)�}���h�{VN���7�ck֗6L꜅�6F����G���Ӟ����/�iA'Й[�3̷MH�O�plT:g�-�g�x���P�����{�C����e��.��u5����	�qXH��c��@k7�@<�00���N{�۷���t�}ϖ@5I��_�ݴ�9��
G0z웥gfNq#�;ēYp��H³��J���mBf�������ۼuw�wPj��"���Z
+�2�$�Ũ�N�����YvEw���: 
ֿ5[L߸{DM &P5%�ʲ&��@ݲ��X��c�ŝ[���I�'r��
����ܺ��o~��a��ߑH�\���?��N��C+P��o�i�6�f��#�`���-����Iz#�lđ�YJ�$w}z���V��B��o��AY
�4�n����]�����(��t!ھ}�*�n�u���!�����/^<7@3���NҬ���2�������,��h�W�ZPs��<n�4��+�uhf�I9OYɗ�N9_�bd��ӓW'�s���S�{��+^CD�L�/��g�?�B��r��x|��O篦'U{G�"���ē5h{�ԯ �M60�K�Za��'V �S�լ~��3>i3΂G�O�7y�4�����O^�%��7愚ϬY0����,�������~�����{�ӟ=n e�]�	i���M�gֆ���A��j�g���?���R��6a0:�j,�"��3�\0���A�$��N�ce�?
1��H_�̂J)����_BoЏ�<�PK�q��0=�>��4�~r+���k��P���dմ���t��W_
W|��9�f��Ϟ|��{6;�.���ԫ٠�=~�����F�|��K�0����1�g�ۢ'F����R�M������8�y\c����D��^'i[�b1?�N,�'�a��?;�GiR��4/ΧE�c�΋��'�`�ubyE=Ӱ�i�Wm�(�E���� �-"Tj�V�D7WU��ly�:Ƨ'B�C�Q�f�")�e����L�i9�-�837���.��rӽ�%��M��ai7t�cE#hR�	��:-?����Y�J��V�o<�p9ݧ�|JN$Y���e���@�	��D����?�I�;xR��q�����ԕ�y�4�"�Mґ�X�-l+���i��:����p�
9qHb<��S��������c��E4�hE�Ӕf��K�vj���8��M��Uh9:Zj���� ��OO��Sb#�2K❹g�h��	?�����m�f����^�V��[�B�i}�݈3S�`r����b����Ė㇡��e����	B*��KdS0;D9==�u��)⒤7rI�C�@�:��e�t@���Gw�M���eMZ��٬=�����'�G�8�fm
�����Y"ޙa��1x�'��'u,~�d³ܺ��6�Bw��׶��3�/�2.K$P��%�n�%v�g<���m�,L�ɝ�X�Y�=��y
�њNU3�L�q={�Io����eU+x�V1g���v*]�&g��7�9��������n��	"{qQ����a��4I&��N�6%Â�Ere5�Ҹ}ҳ��ڈ�9����DS퇢�Z�xF���'���6X
F�.����L��q+,�=Lot��#X�����G)�&c�
�	�C?|��G��sw0硊�<-G�)���ū��]�A�)��4�b�&1��j����<��k/�(g�G���`Y�U-܉��W^2���Xa��+���2{g��`��.���k�(�����hV��^��dn�w�r��������eZ!�>��s�Aݿ.�hУ���M{qjM(�����(�8�o�$C�1ac$�*�:J���8�db��L�<�N��-�Ua.l:��0�Ɋ��Aq&�!:.k/��C~8��%!N��J����	15TPl��ñӰ�Q��BM�K_�j��^DNk�E#��v`͡��o���'Ӷ�l��!��f��ph��V�g���qd�۲��$��UFv:jF$z4;w^F}ښ�lG�����Xz��M�rm��=��n6�V�L��Ċ��m��6=�����ĵ��
��%�|�n�2-bH�ͭQ/ی�,⤸tU�҄ C���]Z-�I�<�,�x���`�L`�tG��z��[LbA���7�_�Ԅq�i�)*|�,��0�-l�#n�C/s�9�>������Q��1��xh��b�Ͳ2�XL �_���jhB�� 郸���&6p?'nd�|k����uܐ$K�Ϫ�#YO\�|��|���Wi��4�lL�%�'ͅ�;�lơC܍�%��pj,w=���xĚr��*�*��M��dl���["��I�q'�fw�#sɼ_�v-���SL`�U�ʓʓ����\y.=l9FU��Q��N�#'A��������*k�I��"�R�d����N�;#N��?d_\P�{-�i�/��֎^t���-bܖk���K��Ȳ��'oˆ�Y<4^V���,Q]VQ`Œ h��&ţg�8���	XlҶ((�wc�e�,9�RIl<�K;�F�����Rq���kW��>�E�\�� �W�K������a��.��I�F��V����C��Ø��^���H����`SE�h%W�� d��ڼ����L�IE��.��&*����6�pl�f|�}�qco���+Fh��6�Vu6繍c��^�w�ᕮu<y���ןgiy����C+ABo���B�E�]1$x&D�\�Yc�M�D��~/�h$'�����#gc;��Z-H�͝��,��s��HF%1����u�!�?]U~l���[)��3�w���W�#ZΖ���	��6�.�0�:iUqz���/­�#��,�Y���̹�Ί6LǪX���p�4m��U�i#p�!�P�8�k������C�q2B�8h���y��_R7���C��YD�)��fP��k��B�p�G1S��yiP�	��d	z���W]���x4��"��d�D�&�ZKw?�Ԝ�*wɷ�;Y�1V�<�bG.
?ٮ�-��:�'iuQ0��g�i7A�S�J��1g��yF�G,8NQ�50���sg�צ�C���*���	�d��JͭL
�3>���B=�h0Z�ZU�X,� ����&�1+$�)�e�"��"�O[�K�y�,�P;	�$q.�����7ƃ�5[Vy����,�T��`�oB�]pb]h�
��,t���}�{�Q�cm�q}z��X��Q{��I�7��4m�U��>xe��}����fjg�Xc�Z�9,(�3�*bw�]�!r�:��|��w��rܐF���u����\;�-&�~�����li�J�����8f~�6-���N�6�\<��G�c�-�ru�$���*�H�f9�<qj�4U��y�>(҉'k��)�eA]�Ƙ��8�J`4�`��CAg?�7�k�Q�SB?ô��1��~�t�q0�)�*���xB��'c�*G�F��'A����7�#���	ޏH��	�����ml&A��^���w|8v�*�����[t��ݽz����xb`&0�$�㹎'�WluǷ��ə�΃��᭾T�U�j��\!��k��N�Q���γ���Gc��q���Un��tB6qu������������8>s&����#E�ݚ��2�@��������+W\?��ԐS��Kx۪ah�l���zv?�������$�<��4�X#>[{v�)�y��Rn�����5�8��6�ŗ�\������鱥C�Ӫ�������1G�'��,�I4Q$x��t6]�1,�r��\�Ϗ��Q��4�}hK?r7JVLn�OV��=:�f^�!��t�d�6��o�m�5D�&�`�v���G�C->[��yf\�gڹ�oiɪi�a���FnvH�).��Y�Li��|>MV��{�/sݬ*�y�N'K���%��D\<WhϑT�ƎS�rJ��<Z�Ŕ}���u_9c���o6��W�l�~����,E~�*	(<����M�Bi�b	hEs�h�p)2�W���yK�y\dU�G�'�U���<�<�X�⨢�	�!��u���J���c6ArG���>�RT{s�e�2��YC�B]��^��EKL�*��4�R73�s�j�����Z��ƞ�:��J�tw�I�~�(wZ���,�чXk)���֖jHB�9��)>S_�%��9(=F6����zE�ER/�e���n�a����\IB���~:����=��[Z� ���'�4=�Zhj��3�g�	�k:�<H�%��Ժ=��2�{��{iYMSg5�mY� �2X�ޥ��:���ob�_Y%.|�6s�q�>��âYդr1f���+�&(J=�I�i�CńV�I�^�*��X�h�_�}�h"z+��QY�%��M��P�٨��I�K�"@��u� kj�[P)k�%�ֶV=h`�F�;�tv�-��*jd�d���s4�:8I�
�o�}w�#֎�kk���e�:g�ϣ�f�YG�mL�PI�AdbY'.%�Z����$X��	�r�ŝ�%ͳ��B�A2tfU�M'S�	�B����9�(�&Cg�s������y�Q�[n���Zi����,���++̟-�Qi�i�e���4�M�~�y�l	��@�O�,8I�[Z3ޢNť�v�[��x��Q.���P%�T�&$���,����:{y�Up]��>�u�Wc�!�+Ի�
���-�>u��W�eHk�r&MZ�x5���^�-�N�U�.���KkM��`f�cxܡ�v�k\M�.�0N!j�U�Z;�`Qk�~���l�
v��'�� ��WG�Y��٥��wzGTY��󠳖-�L���?��^��XΘG�Kw"ͪZS���uYu���-�!�0�D�L:ZK��I��:��:'8/g����L�zH��g^��A� [�-KV��$Ihz+y7M0�p��$k7:O��6����"�ٚX:^����DWQ�5�y���A0�k���W�wG��#�(�$�.�uz�u7�˺Ȭ�3ͺ+P{E�4D�%Y���J'<�{P&q��ڌ��~����*i��Ђu�1�Y/_Z�]F���;M��N���>�fW�s$2��.s��%���8���wm�эs�,���u�&�J�C�[���  ל�~u/�N�P��h^UQD��n��W�`��*Z�� �;���L��\rBwDn_�ݙ�:m-U�ny�[���t�"g?	�v?�X��>�w��I�w�X(q�����)d�d����mh5�(n�d����$�e��:$t�����,s����%����(bxV�~\��S�;v�Ƶ)�E֚!#q��a�~�8�8)��|�y�{���R��*.`|1f�_�mQ��2���t=�k�i�hHZw���nY`)�9�~�^���?��k� ��5!�ԃcE�n��B��żn�h;5o��~?-�F�^�*wT^���oYL�X��P�
��]���$_Bȸ|�C�|�&T���,��D
n��TX1*�~�X̚�������iQ!�+�֦,�k���>���v����?!A���>6Me�Q�+�=H�p}<��í��Sǔ�U}}�O�⯚�)���W���5�4XS��ڶ��=�y0I�/|�nk_UD�e]�]��-I�������t?_�?:���^ē�t̉���
�El���دm.��ĵM�K�w�e+�k��ܝi�ꨍ������#�c�k�֗0�����	�Z����̭�0)�i<(�>j�>�*��Ғ	�X�O���12�R���U�Q�U�x�(�V%Q(�騘K|櫱���jn��<<-	��&'�l�����p��x���1kT!}#����	Ʌ�`E�\�ܹKɑ5q2��l���(��	*�>�Qu0	�z9� |�`E��U���^$M/͢������;{w���	!����ZP���4FC���,�����۾�_Ʊ����(��}�,c���7�;�}y�/p]%nQIBLU{�|l:��˰(,\W�����9�N0N�Q5�l�;kË�W~��X*�Y�Ҥl��a���FāE/�B��|�	�͊��6V���E�iB��b1E�tU���K��t�i�E��pTz8av��,¦(���.ycW�E(��������i��R�1U�f??��W�h�o���ޖ��o*�Y{]����E�����M8�ĺY*ޒhm:me�~\.o���u�&]u�$V�㱆��a߮��ƹ#{,Y5���g���eD��`�F�r�o�*y�i8O����%�r!E�eyɒ&Ais\�9G��'.0�`r��M0�Qs�g!WV+`]�M����;!2M������Wl�f:�F�����Z�?>��8�:f��]K�_��^ee���O�ӕņ���8�Ǌ�ob�Ow��ӛ�V��o�%#�I��ׄzm��Mw��m޵-/�c��L�)��vyb�b�M�B�@0��aeڍ�B�,�vY�����C��!٪�&�����׮��Qf$
��1�JW�q$*W���cEf�'4ա��;z-�|��O�kV똬��;���z��ekr�{��r-��n7�>��P�x���O���w��qV2�.�F���ru��
�%�G��R�,��l��/Kڶ�q��y��e;>�ubt�Z���.��dw���l�W�TL�4C�R�}֌FG� ��]����j�L�v���.Q!o����WI���^W�{�f��Ӎ��#��×����	�����ʢ� �k��>�$��%�aoB�g����U)����K�6��9�֔��_��b-�ֶn+kڋ��I��LGz�ئ��;��ںź�3�T�а2�˯�t�إj2����i��kb���dL�y�t��'kc�+�BH��z<ĕ�?���8�Hϑl����2KM0�7����E�-�Y��,`���P~�r"5��x�$d�,%H瀯���W�L��#�}��7�J�K4�^^9W��^�X\<��%3�^��*��Q�u괙/0@/�ז��3U	�dK��M,��U-�,�o�����,zڄܫZ'��%mӥ"h��?�n��ăG�tWd�"]�X�f�V�-�]�l�{tt$��[�n�liR�=a�IZ��c]��@�)l��qY|t�骒�D��c�S��Gx�d��r�vW�Le��sp�i��r��˟;3_�.M���:P*?��n�i�}��ٮ�WS^�
�;���1�x�����Q��'�RlP� ��u���kI���|�J�$���\:]ʣ�$i����nR8�`x-���ߒt��c�Y���,� ��ߋ����y�{�cef�Ī3ԙ�r^�&k�Q��M�������Z\�b��!�x�n�Y�X��~p�̞_.�4�b'���x@㼍�������a�g��0Hn��h��+]w�h����a�d2��|��Kw�@V����5�䟵�X��[�Xو0��[�ֆ_u���_"ۦ�[#��Zc�e��{i��s������P�Q���q�Bٸ{'�e��%�ɖp���K�;���*�I��n�,�6�ʥ�
�]�C��L�V �f��\���X!�!�'�����k�H8v�:��^窮�2���R�U7���i �%t��V�q��٤.R�+����P��A޵�(���i��7e�"I`�A�Y֍�ˢ�
$����!���d�I����!
u�ga/Ț��
��SaEz{~ҍ���.�t�̤�sho�g�����;�煇��U��
�i�r��W�k����c���c�l����t�����&^<��o/̺\��KY��d;Pf�:g�r5�vPkQ̻ı�JW���cR�t���?i.���^μ�/I�|�
��=;�ؿU�Z��}��XR�J@�\܂��{6���è..�E���de�q��僿�ǧƶ�fi��r�K)2�1]�\B�IqvDi�m�;����.��NA�X���|+�rv�(ݳ�fUj.�g����� �<�tE��_jy} �򹯣�6���]��埗E%�
�����m)B�Xgza;z��xA�]J�M����ZcVM't��ǭ}����^1�CfC��D�kgڬ�$���qvH���_.K.~����߿�}�fz!��?�r1����O�1�4�JT�M���&��-��k�++�v�ڇ��s]U����������;��JkC_ۣ�Y�ג9ğt��~����^���寋$��E�z�o/w�	x7Y��U��Ig�S��5�u����_]�����5kf�?Ck�d\�k��+����;??����h�ACu�橗O��։ϳ ��m��v��$lq��c�-��|�N�+���m'�;���&-'�8 ��wi�^���M$�\<�{B"����խ��s�Pg���==G2m��p�֟�Y����= �:q�|i6J"W_]���Ō�O�,���v��UI��74�>���6箳>���P��z+̷	�,,W�/��� AFv�l|��w� �ֽ�=W���}+�7�#�t�ڮC{:�fV9��'��%��V�i���,��8�,S��6�(���H���_9�+ߦa��K��z���\r٫�;uw3��h,A-n���<�C�;E;��WXsG�̇s�[��G�u�uD��ǵJ���8�/|�����I�vV��*X���岸���[bL�I�w[������+�.�����\�X]��}�ݹ�+��.H���l��k�>u��oB���Y1�p�$�������4H�5��,wg�C��ug=/[���MՉZ�gi�� �{,��`H���'�n��╁�JX�����|z9���-5�������r���b3�[�liV����tqĒ�m$�В,�<�s�^���_���g����H��
�\\��_kg�R��R�ՋqHT���ӸV)vU�]��뾅�����"�f����g�&k��\�0�c袄��k{u�z~�w�%z�S���HW������1��Ss�t�_����KlWͥsL/,�ڨ��	IV� �&�̷i�~���{�ڷe��tv]�})?]�U݉�~��\��-��٥�z[1��'��\|�b�W�9�+��x����x��7�7+����%;�]�8�(#/Ny9�l�Qv�������0.���_����������n�⩹�����4�%�$ɥԸ����4���\��p��/e#ݣ}ɬ;t�^0�/�Z��d����^|z��9s��Å}Y�3<Ѿ�BzمU�d�˵�t����/�.�g�i�������zͿ�C���u�n)*�d;�J��e$����o��Y��׭F�W�/�s� �y&S7+���!�m_�j�Q/�ꠝ5V�t����ƣ�bQ�m?oQлt��Z��18�M����H��y��JW��d�ww��CQ��Rd��Z]��1c����+�������4M�6�8�4���#~�����u��^m�y�:�I/9~k��h�^��?�ڐ\�d��|�V��@�Ju�4l_���u�Ԗ�0�6���G���
G������Aᒵ��V��
�� 6k&jwչ�:7�����;��<��f�i��d�e�l�U�����[M����Vlr�����9+ *7�����5��gˑ�������/C!� ������ג�b�O�5�:����ZF5��E�h����$�91y�+��,��朵��xȫj���Z3S��o�۲�pƚp�>%��^��*^r����
�fտ�r��Ь��C�q2���^L3���c'�[DD�$ĉvn�M�<9I�?K�Bӱ��I�K_\��9]�Nڹ(�$Ĭ�5��Ʃ�a	�>Y�t�N�.�3�.���:����?���μ��°B����.��V�ux�i�74I�x�؛�`���g~�^g�i��H�U���ժLY�$����~��u�}^��4�\/�#�<��-7du��ß^������`�`��	1�r��2�5�N�r$�t��Z�h�kA���gi������ޛ=�uw�Ug�K�ht��F�@IQ���-ɒ5r؞�˄��ᙉG���0�����<;�+����'����F&%Q"E� A;��z߻�~��~�yN�:˽}�R��ty��:UY[�/����d�jKw��6ne�Ko�+�-�ڑ��2��Z��)R�F��4G	*�p�b��}!CL����y�7��u�G2FQ�������£r�#?٢Ȧ9�/�:3��'����{�_C�z�U���U}
�ʼ��>v`�wwU�
�����J���!D���֕����E: �*�m��q�E��袂	�g�����3K�ns�hA�܂�1��bVZ�'Lf���#�Bٟ*=s2Ug��N�kK���k.�#^�L����{�7���25�w�� ����g�a�)�Em��D2����JE]�{R>-���/�+]�"IITq:�B�)G���(�F�`�_Ǒs��@�e�GE�1�튻V�0v,�s��|K>��(Lޢ:�_��=�������V<�t��f�.��T�����Yws��X�����W<��@]��̍����9o��E�m��:eGU����8Lϻ^z1=�C| �(�Y��f���<���5�u�1�%�cƚo�!
��_E��ŷ��Y�ki]V$�x�$j��<������2�9Wef��S�8�CeT��+FB�\	�X|IYmm�c�>R��W�w{�t�n��e�i��ꅋ���J?[�%�3LuE������,ǚ#{�J%�����zr|�՛H�n֋��T�$�6�䏢.�����̙T�E���3/�zb�tWD�OJA<:]"tbz�KH�R��{�3�⇘aY4+�X�5��Բ�����[&5:�[Q.�yo�U�蜈) m��=�Tb��2sbY��٦�S  ��IDAT+�� ǮC�����%��l)��%N���4hkv��E�2C�=��dv�Ȇ��;�ɥ����a��(���~w�UZ+A�J�m٧U�G���k�h6�9ّ�6�<?�i)ܜ��ePu��n�
�2c?3ߏ��\Ɩ���V��k�ך����ꓸ����NOP�U{P���n�!5�Y2��U~��0dG���B��NjCpf\��)�jOG�jZ�H5�|�����La?d�Z��=�Uz=��Н�Q���;�}���3��W�4�~�+���T���C��6
{�O��7��T���KR�!��g�o�i�k-v��^H^F��+��<��}�E�@�����*\S�Yg��O�L�Wb��,��o`!=�C�qM�z�N.�N�����>��?;��W�e���L�Ry����qL0Hu���وi�D�3����m�gW&O^��!c�d��>��_�~�5�Y�-22������������w�h����?K��3�kήɣat/�ă�`Y����[���� V�&���}�H�Ȓ!@�P��'�-z�D�a�!����g���t��F���̎��N����E�J{�ϯ��b��D,���$(����W`���+��u���Q�Z��-F!�=�"c�J
g�����PR�l� &�,=���8rF�^r�����c���.�N����ʺ�;�ZG)ӆ�q{w�D֊3���͋��f�I<[�bD���MBo�Zŧ5�c�H�X�X`բF�N����|���E��~BL�>�'D'��5}�[�=ɝ���ʒ�&N�j��r)�nv1$�I��eF�Z�<�R���u�\1G��lY-�8�ꈝ/I��nzx`�{(��7�F��:	��\���b�L���Q�of7�NQ�/��yFaaս�!����4e�)���t�X�e˷g�h�񬲮T	R�/�^e�{t�W]7?fm��T���:	�h[�#y����M����6�щ�6��L��MA�N.�!�����@6@%�e(�pQ$���I�*Ao6˶��jY��V���L�Gf{�c�	��s�06K�����Ce]&��Zv�Ĵ(癤
��m.�0�n /Q
���1�C��Y�=�툯�H��Uq���Ӽz!����3���^��/5?�����I0�_N��s�J��]_I�.�Ѷ�f|v�����B��9�#�pO�|��H�3�ϔdJ+g��!'/������Q]�{^��kz�+�O2��b)��I��Q��m���ϙ����n�b�d�U��O��A���w��0�=ܫ�<��Ê�2H��3<�n�O�ݫν�zC�hNM���ln�=ʹ>����𗔓���^����Sf�aa���ɰ�����_���d��y�4��)�s��Y�Ͻ����<|�m���Y��>�}��ya�{>OLLWTD�mL���v��ZT8uO<�G�� ��)����+^t\�<�AL!=}(��lLi�Y>����bVٷ��+l����#Yh�Q�7���-U�
��ӧ�������S�ͯԾR��>J�E��kl�K���Fd�P{�tC�Q{�<ɜk��ݕ�kJ��w�2�9��R�P)�,-m���Ë�^�ͦ���M����t��oQ��hm�t��g���2��w�Ja��G���=*�֋��� 8��N���j�h2﩮=�/��B�>�<��R!Ύ�X�����ނ]S^���K}���Ά���</�+;�?Cޮ3mH��[52�40?e�Wd�܏�ɦ0S�����A)li����m����~�<�kny>���iwc�ɮk�����s�>��� ���qW����w$���s|ҳ�*�[���gd[~�:H�}�x>�!,�A��֎v�"�����<�+H-ģ���+a��_
���D>$��'�S//
���5��If���i�ȓ��٫�܇f�r�������nXOy��U�VA���C��fp��#�&��P9nP�V��
���F��|5��JO�^(�$��d�3�Zm$��<�ە���4E��dA�嵔�����rꮵ�e�d�e)v��|&I�ەG���p敖�?�
�8q��+|^8*��7��M�嗙=5{��k)l���Ԗ^j����i�]x��B��L�����ɯ��Ta�y$��)e4�^y2O�hZ��/��I6��`Z�WH䋛����f,�0�u�g8j��.�"y��E�#����^ܠW	*ݺx��%T&CNB%���������ygS�k�m?��G<e�`}�g�13����sdd��$��nR.]���8���0�^-W=�K}R������A��5�q�+{���ɤL���e����׀�,_�]�.А��x%-�i_��U�{_p�>$�_eڷ��5��G�C�r���'��2�zWp�y���5����{�̟�U��f>��\��?Pw5ݒ���Xv]���u���^��pi��ܸ�>��LV���ԍ.��(2 53+z��+y�?��1,�̔�������}�v��ZH>Z3���s���d�H/��d(\�n�y���Q4�(�(R/y��D�ϓp��6Hd�O.��!NpG��8���GN^}��CCg/�f{A��!WA���h}�R㞚�-���<d�0�|����(�c�.Sx~~�iԞ~z�X�F0?C2 �O{{��g@U���S�I��j�4�A�����x��n�r�8�G�)ED\[$�Β��nJ���I���^-�d�L}��Y|��ٽ����_�S�R��	]���R�(�fL$��1� ��r?u:�u��;��[�����q�|�|ٴB�Dޯ9��^���Ot~�d^��[THF���)�z��u�}
���1w�N|�.��V�Gi�T(ߏ�����5y
��.@F��Б�mu��(��Q��5��,� �ͣ�67m��b2)�$
�(s��az����l�_ϥ�)ӠR��.�@���χL���U5�Ĥ]�'�[��]9�)�f²/��^�]�袶��^le�oK������a����g���cL�	J���1�=C�J��4$/�3�K��"��)7�8�� ��$�%x�h4�}?�t��y����f�a�$�(�B9��T�VI\��}(,������p�t���L!���<�V�re�]N�[��7$W{��*l�xh2����$��oS��^���f�>J%I6�T=V���)^h����z/����x�2(A�e��S�K颥(+&z5�ȩ��c�����~n(lE/)�y�g��yɢ��T�!�
�)*��.[�و�nB���ϵe��ѭ]D�?����Wh�%��#�h������4D?�3�
���.j������W�@�P!�赖zѶ��*�= Z�h�Yk1y�SH�fd�\,���h�ڍ��ӹ�ڑd��*����(}8p������?��п��|�?��A���S�W����}���g�$�>4`�3���m�9h�=�����~�*�~l2��<����0b@|f��b��^y&��)��5�[��k*7"ʢ3�lY`�n
ه�lrMn4�[��W�/1ư(q2��83���;�Jn�H50��\J�|�3�����2��/w��p��x�Μ��Z�_Z}|�ׄ~H�o*kt����x�B�/�èY6+)\�}H��g�^Q�bUњIS>(ͽ~�� T*a�0<��t�m�^��]�UEKWY3̈��b�Ӂ���'[���[�^)�E�g����G�?Jj_Əm�øtZ��Uw!�]]Nǿ�$�˪��X�ݮ�oQa�g���e�^
y��AdYdi��|��H�*z���[��'��S��f:*3y���^t&h�6�Xk���Z�+�o�$�+��j0�� 7�����^���N����~����G�(y�Үv 2�'\�������B���B����j��<1��B���pB�~`O|��Y�\��c�1�*��6H{be�R�92��e�&�u���R��So!��S�Sq�Q������$�c.��V]�S��X�'[�tM�x^`�b� K��]�6l!I{��+䟅�WW�3��S�쒹���f���S!P�W�r���L(�B����TE��0�i��t�cP�W*Ҍ�t�����B8����XL(40&C�y�[�2r_Y�0S]h�9kǝ6y8�U�
�1�K�Ƕ.�`�\��Rn���h�S�_�?g,�[��G�����o��M�{L!w�o��a����f3��\�j�v���ul��*$�&f@��?Ks�Ƣ0�S�d
�g������(�#r�>�P��Q��Է������)Ϧtb?� V��B�,��T�z��b�{mr��^�:OL1�Qy������2v�$���C��PI�%���Ӻ�������9>3�zp�T.��b��j�X�Qo�Cl�H���%o�gv��ia�n	�����0͋Z�8�J/y?�
y��y��ofI�oD�no]�?�w�o�ei#�=����L�����
Z4���Im�����si�=���C*��J&���S��	�ž3�O[�������b@������{�,�B�lʏr����i�]Ԯ� �;&�õ{�!����������p��M�xE!#�WN���ޓ�$�Œh���%�(���S�]�y2/�)\Y���<��u}:!��d����BV���+�`K�i��1fX�y�zt� ����$�����!�u�ͦT�ìt����(�d���B��e�g*Rv�͖�Az�~hw�y���u"/T�_�$��Ϧ�
����pu���3�U�����~�-�_QQ8�fo��=�
eC��=��B��v_�&C��QQ���ⶏ���t�ըLW[�wGjOX��!L�Ϸ�����J�T���̴��*��b����9C���C���V!X���3�L67��F�w�2���<�Y�)pO��iy��K���O�E�	��lY�C�A�H�/|7�VKE��d>�����'>�O� 0[��bnO��ٲ2?����A�]�V�ߜ︴�b�S~v	|2H��{Ϧ���v��&���{�Hԑ�a���}(�RIF�T*b��|��|6��+�7P���N�S����T*b2��d�xe�]������d��0
�؁�5T��E�(�U>����V�i�c����D�ϒ00,����#Ms��'��^�J�M�[�⩛D��T��j7%����bh�ڪ��z�A�P��phlxcc������Ÿ����V|X��.t��&�24�U~�:�J��l�}��.�A�_�!'�E�W+6MSH'�\��&Xr��-�a҉�7��I����#O;@3���p@#r�s\��R�>Ow�[A0:��z�٬����0���~�w��
�� \m�+o�δ��G-��=7���`���[�"w��X�b.�JH��]�����h��i��,Y�|��(����I������|�}��}���q���	U�B1{�J�e�ԕjlc0�j�7'w�G:r�;A��n33��<�# �.;Ģ9�#� ����������,������ []�������* ��� O�����(~��d���fC"N�e���J���=�>���2�U�i������ ?<<uH���Z��hC��F�=ѐ��N�VÂ	I��=osssjr��?��n�e�����V�<��K�D������[ܨ7�����x��h�`>�	�$j\ZZ@G�-�P*U��ǉ�rM����D�ש�I�Dkgh��H^P����V�MCS
�e�iۄ���=G�E6��o�Z`��^�D���p��ߠ�fQ��$�cI��ށW.��,//�mm�6�s1:(�r�;�P�đ;��
O<���	�'����N�(ڈ��P�<zkbb���P%]SF�J�Y�������!�N�?�?QhAJlQQ���&����@4@;):j�!K:ު�b�����x�eP��C[��1�##3f	c�,Z����U�B�@����o�`�بb)+�F�/E�F�x.m�|�}�#��Pi���lӉ�q>hYef�k�b�"� Rl�>�D�����ev�fǤD�A����ښ9R�J�AI�h<_^_�z��A�)�����,��Q�>�~��/�����*$Y#Z�;;up
�G�1ọ�L���HK.\+09� �����H`;V�e��-�FӢ���2A[J���F	��5;�1�u�n7~�>���&x��x����H��B?��0���'+����ٺ_��g�y���8 n����D��:#Mc/��4��R)�U�v�M���."?�N�(��(A��LC�j��K� g������.a#�J�La�x9��@r�r0^Ѓ��� I��:)�\]Y���ܼ)G$B���程�zn&8^�mB?X�m�����`��bA���t�����y���%T]*���M�{.�� K~	��C��_rd���	��P����WB	�o��H?o�eͲfE�V��A�1��[9I|�\�=�y���pJR�,���{�VVV�_.ah< �k� lI�����RQ� "�nRl0�#�C-�p'�܍Ut;5�TV�M���ͯ�V�[:��6���t!��s����bkSq�fvq;�Q�	N{%�M�7��J��H��e`�j��Vie]�<���`qO�J�>���v苝'b4�
%�+�+\&�0&r6�T8f������?�-L���A]��yEav�{�[�\�C�r��d\8G.�=A$f���U��2��'�gz���
�!�ԡ�1��- �@;n���q\ rtW�#�*=���0��<p�:pW���CD�#�I��&{�ed�N+G�h�>:6�T�7�G�IT�ц>�$
��L)F|,d�%s���G
�E�#���V��^�!�W``�3�([XiC%Z�� (k�U��`&TI�&�h�)��2����
�ؠ��9�X2H�����7�?��l��$��J(��jq����n�$�'�.��m}m�|��[� �^vDGGI�f�1.*���g�6Ɩ�i����JYb	�nI��z>8� x��F�f+	����u@�"����������$@ܑ1�}̪��6kZyx2���`�,����X�����i�}P"����^XXpKį*`��Of�ZR
��<Sq6�H�T���cP���Ӡm~n�$@���S	:(v:* $����%����@"m��*eY#�G�-r���AVv@���I�j|y . ׀��c�->���@x壝�Fstt�P�vc�D�aua�q#ա���d	�٪�;!qN��nwZ��\1v�nw�5���#�Y$�B�g��h��?93G`�����6Z:�����)�(�{�F�F��C��r����⍀p���(�<Bxl��]-�����*L0���&�h�戛��V�Q��jf����0�<��uQ�U|Q��2����y�S�Ӊ�d�:w�hQ]���b��'4ٳ[1D4�E��x����Z��AЎ�*��7d�ب�&���p��_#	s����z�t��sB,r�
���2ʌ��ND�����c�/Q�b�B�9�W�ݿ�z��b���� i'��:R�V2#: U>��n��[X�XЊ�P̉��_�O�W���%E�� #"ǌ���jh���xD����;���v��Y��M?����t�h��h�l�a.��`X�W4͓}�껞X\�B���h���� f%l�*�[F| �Q��G�c��R�~&C/�:�K���������Ӻ��*S�|���;�`���bka��Í*������J��Th�[���f�������YV �h��Do5��_+���v���D^p!TK�2~���0X�OJ�uMh8|�������X
�����`DR/r�qݕ��%���t��D9���	��n�E�G0I�Xp���'�@%�H�k���U�>�066F{,�*��8��֎8�����9���w��~��۷�"�j�Uj�#v&�](�	~�SCgoloo�x;�++k��Ę/�5�? #.zJ��h�������i?��}b��)+����w� ��G���P55:>���<FcT>�P��~��4DƁ���	mBI+j�hs�.����>x���5j�O��"�iǾ��]�m�R{d�Y�W��q(���f>����6kGr&���Ob�o'��Í�-Ln>sۉ�HT� �l�&-(���1�g�f���S40%	���F���`m�^t��Q1t�D� �����1�<�^��[+��]��>�fo�k7ގ�>i·�����?�9�i��Ω�b7�l����'N�������=��� �`:�=v�ӧ0����K�������ښ~@��� r��U�h���.V~zp�.�<��Ǐ��i����w߻~��*|%ֽn+hͬn��}j����+�c��d�9hB�Y�(L���
��N�m��l�t���4�N@�N������̙3O]8w��Q1�A��k�ɬ��[51붿��1Di*�tE%�"IȘU�=��>x22�;��%��>qlQ
r�S��P���	��g��Ж��/��o��/�����m�[tE��=^|6�SoD��+%�� :X�ã��Yk�_2��[S�s�{$�i���8�{f�j���,;u�$xΛo���ǎ��>�NBN0FV��y��UԎ/�S�a099)u�]�~Q�;��}�'@�ի�	;���bP^�X]�Juܕ��ًo�O����92¦���54�\�zuz�0(y��4�O�7n�i��0��UGfR'��{u2RJ��Fsrjrr%l߼�<�F���?���F�	R�F��Mnn�ގe�����U;t��Ș��M��b��W?���&ɀ�l�L��f��{���Nc��Ё��
v��k[xH�sx����(Q�!5�z��"�QZ�[.BB՚tr,`��OR�[JBf.��7̒�j�z������Ĵ����"GK�6���M���?3f�FX�˴�V��_c�1N�s�	�$�Z��u�]��;m9 ��!il�
c��L��R�i3>pI*`dۼ�n��� �}�m9�2�{��*n�'4ļ�KCXE�&�jc{��:2V�>�h��TGvm���u?�i�=4�f/��}�[�܁]K��;���'��+X�_03u�����O����?���/�������� ���,^i��E!Hk~X1��Vt�{U�Q�0���|��_��W���c�aP���o��_�%
a�[h�0Ŀ�MH�{D���TjF��;�LeQmU��e��a
,#OD�aR�{K�(�h�F4��,1��u��ǟx�������}BH?Z��aK���n1ʀ����q�M�X�9׎y��|�U>BR��G�Nw�f�sօ�eU�.my�`�<x%������������-\W�<�s�2�l�A�%<��s�\haa�^k���N��V+e�p�}ޘk�a��s��Id����7� ^¯W�\�8w�~:�<
y������?��Ϟ={�^�|�0~Eix?�|�p�o~���_�x:����P9󅩩��Օ���w������m���������߻$7u��k���� o��������_m����^{l��ɟ�	����
�?�#~{�n�����z�g@0@��O� Ͽ}�.�������4���O��p��s�=Nx�����;������'���RS�~&f�|��th�,�\wx�U�z�C�{�*�|q�|F�y�a���7>eg8/ٙ%�p4P��@^`V@"���v��yP�3Y�|�@<��ut �wpr}kܜ�@ �I��Ff�@-*��a�[�
Wh&�m�����'�oFS$�j����cb|�7s�=��%/����P|>(�+U�r���hG��ق" ��JS;�Z�m|gy�o�4m�sm�,��2��T��b.Y�ֽ�n��1Jӄ̪%�>6�GGIÃ� p渥�Z����ֽsl�!O�&o�����N&I櫯b>H2�������A�-���*V��b���Q�]cw�ت���@m��s㇎t��޵��޹�W�K#w�.�/�i�����{�dE۲����
�Xlu:]#�d���?����?�%!��c���,�m�Z�D�tS�����up�Q�V�<�eƇO���[*qZ�-��5��l�ܖb�f��e��uɱ�|��jx��G�<�v�ld��R� ��_��J�
��L��U%��Q�o��a�u�!�<��Fbt���K����ɒ��Av�	���Gn݋�4�P�(������~�"�E�Ϧ%�2�u|���5
{7(�J���V��R���kAH�6XX��"��L;��r9�������?��˗/ߞ���a�J�	]J<�>8��c>�:��[���3�+��C�_]�\��l����ƽ{w�ju�'� A��O?�(}��M�@���7�����+��ɣ�FG��0�\Y�;0s�H��v����OO}��g7V׿�͗67w�>~��͛P)����NLN�P�����x����ܞ884t�(\�ܸ𱧁>'&H�9B�7p-�!`�����ޙ3g���/��꫿�˿|��������:�4�
�;ypqiqyu������>����щ
�����of!d#�|���#�$�,z��Q����~��|B��v5�I�N$�����T��(Q�e�:�Q,�@���N�f�kY�ly��،��m1��l�#��v��2jDOnn�>2�G͔8��Ab%Lï}/�^kWƞQV�7��6�x�Z�R�T�#��Z�E���Ա�Tb\�>ٺ����PE��i��%��=;�3�l
n��t�ġ*�|ɮb|HX���+B'�K�&''��Y��0�7779zE|�Q�b,"f�x_YJ sT�5��5LN#U�� �H �Ph�Rm��	Ê=��K�|?��?�E+Ve<4����o������&�Hl�$�I'�����C�ՐVf�.&D�]�öCm]%*ꯘH�.ב�P��`gA�� 6Ekؗ���)��4���Ӣ3�@��,^qKL0-{�T`V�ӡ���ur�L;�h2��:D~�Ƒ�N?�,���^%'���b�I�8���Թ]��`�l}@yP���6�܇���jʾ��Wl�\����q'��Ǫ���̌�5Y�Ш�ϗ��w���n��ʧ�"��8�~hF����J���!-�w��N[?��g�}%�(`����R�q�
`���(_��@P ���_��'N�~����ݻ'ۋ_��/^|�w��x%�C�v�֭[��;w�P���Ν���W^y��1��566<���:���yd�^_^�z�*�� ����}>�x r�+�;2�iw���=u��9������+"?T��a<@_���ΝØ�����ʫ��o��o��_��7���&���t~~2Ea@ ��R:��@�<Lb�.�3��O��/�Y�d�!�)ѦH�șZt5���Ս3�8���[��[�-Fa
�4��/,B��s��C����4{'��05���d�s��K��On��ƭ�[��i��7��X%O���0��#�@�p�yS|أ��z�O*�������6��h��`W�ͼ��^�V�1��f��4Gj!�$� �G��;m��j@`Zp�6;��!����:��(,��������D���,�K[��ӇCٮcITFF1�v�P�vj����f�����yⷡ9Z�o%FTL���neh\=\���%�Y�[1��GF~ס l�=���$��v��PR9a4�&��-�� �~�V��o�������޺5�_�K�����V'*U�:.��4&��+~��;Ak}{������ߢI2ux���;�:��ŋ����w�Neh�T��:�v�ϱ�XP�Z�:�l���&1\���&���<�j� |�_�H�����@��?Lt�'����n5;��N�;���J����Z��61T�ᒃ`j�ٳ�p~����<�Ba��>g�
�L?�d�>D��u��7�����:쭁�J��u��6Rc�$َ�ns�L9��U��M��6��͑��F�f��*�ƙ6Ɣ���n�T%DJ�[�6� ��!�e'�M��2{��V �g���X֤]��a��O���R�Ò[
����9�WJZ�G��8~��ܸu��b�:��l߸uwlx��?u�ʕRyh�����������7��� �v�on���\�tih���r�����8���9�:�n���S�hы���:�����Ͽ�K��{��{'���s���o~�駟~0?�:62z����#�W�];z�����'?�)0/��ӧO���/�;���1�Z���������~���Η�^ဤ������:��z���/����<�- 5H3p�'N _�	(���?���+v<����4�WMNN.,�כ���t�t�2����Ry��/��o�����ck��_�~�����{ua�.^�x���p��W7��wv�C��F� �E��C��h�b���m�ux��������Q�)�����������-�1N7[�)2�H�)b��=��4�P�a k��*(N��ڶS��*�GJ@a�r���.A����VPx��`�V��e�/���d̑A��%�|"e�c� �uW�a0J�n:BK�,�iGŖ1�e�.��c�%2&�6<�H��wǴ/gC�S�J�h��$�K1f��162�D6����)\!o�Cɀ�Q�5��d���SƟ���zqsüTb��76
��F�bM�à[����wp
�S �(�8���1���/y�E]j5�͉�P�$t|=z�����ך�Tb�1�t8+[90&vf�J���8�S9VP�P�sWZG	o�찏�v��O�o�d�\*�������d֬�l�n�g�8��b3Ȭ�a^#-g��[�?�E���A{U=`2X��b#��6��?e͚E-[W~���.w�UL���"pY<�|?��ښ<txuu���e@	���0����"�d�b�QɅ��,E�LΏ�ଢ଼�ց z M�}����a{��<DQwnς��H���z��������ӡ��Ü�B�pL�͋�j�A���}�_�u�B����]���Ν;��t�a��n޼)�e��w�w��j����@%�p�?��?Cf���o}�=r����,D��ݯ��.\@'��?���/��3_�Y����h/�����ҭT��W`�i�*�`l�GG��2��/�"�,Z�������x�@�w�y�Q#����:ZP�6�����g���x��������AW���ס���zHqC��✷�� Ů���mَ�iq�^�r�d{�fN4FFF&���=�������n�iK���1Dm��!�x|]z�[
4Tm�o"㎣�#]��(;���S@�D;,F�*������: r�'�A�� �P�x@3Yh���PF�vD��9��."���R,���Q�vK��ju܀N2w�ȷd��467�6�w�k�F;$�t��*���oM
���,�u��caܗ:az��F��8~#��9y��!�Y���%�\rtH�����_��?��O�@)��˳�w��w�Yk��0��m�Ȏ��8��ɦY9!m}R�2�s�������g΀
�=	��O/��q�&G�v}��*>5K���M�YhV�&�]�;arۚ�>ޠV{Qr�ZO�U�k��	�_"��NI�މק1TR��
�i 
h[miw<s�[v��nt��udN��� ����xi2h��˰�R�?i�`yh����R��̯œ0ᮃ4b𜽒D2��D�I����h��+tTrr��)o�� �i5��:�U�����X�q��	��ҥ0���^��P��k����#�<?4<r��k�뛣�C�6�-��X������v+����C�)�R���I|x�Ӧ�#ã��&��on�+�ǁ�y�V�� e(����;�z��t}���?~ir�ރm���<4%'�޻�`n�+_������\H huk�Vu���O~��ݻ�w���@�Q�����7�|�K�${t�N�~�w��˫�zsB9����=���V�7 z���.�S��>
l��饻��~����u�V�-�N�j�L�Nޝ�w��M�G�0��Tb��hPt�_�A�%^Cny��O|��|�g �7���hg����	�}�' Ԯ\��|W��
������C��t���oG���j�dg�����m6w�$�<��g��B�5�ĸ�)Y�&� $_��Db����G�K)N[�q�ߢH�M#�T��f�3M��N���$<�)�}��m���US�bP"��$x��tQ�8���;�!m��f@n�sMEe�Y�@A���"���ec��Ų;.=+zC�߻��&s�/��a4T���d�Ų��2)����Yˋ�#'8O`&~8y�$���ӧϞ=��WVV��`͈g�J�)1cW�]�9�}3}�2r��-�=��P%�:܄��S$ђ�.k��*:�k{#E�=L�w
�۔�kahWw�$
nIV��QV0��(}E�ċ����p"�lm��<�n���2���d�����K�{r�]+�9S\�er8�d�6m��x�z��Y�v-�k���Β%I��Y={���k5k�q�*�׭�L(���бcǦ��ů��ˁ)�g@#��555%�jr[@�Q��|�_����0(�����ę� ��9r�r��'�	�R�(-<����߿��K׮\A����!	���g��r�
*�6+~u��K���_z	����3h^kkK�_�z�ͨ����ǿ��o����U��܉&�- �@ �N4�">:�ꫯ��'NHH�.��Ν�7n;"X9)��b�(��B)5t�
�sџ�e&J���6��J�� �~��~d` �]������|Dtģ?o1�4���Z��BW'�iM|���$13��Ah����DV�����$�UD����q��e�ԇ	��,��,�Zh6R)BI��@%Ɲ,3���jZ���^�th���ia[�A�룶��0�k����6t�X�)r �A��$�_?G��B2&�$~�*�V����NfO`D�~��?:<"@�du�ԈZ�o�p��%ћ�#(A.g��:9�cA^�W=�|��)�OW��.��
�3̵&�
dJ��{�g?�ٱ�1й���h���)v���;�fǥ�t��q	_ƇEc
�����p7޷�<015q�|����o|���l�M>}X�ʓp�l*����Mk�J�tW7����"����T��p��n��־QJ0LЍ�4^�a|݇�����w67ס]Z��Sr��	��#\{-���Pڏ��,���p�.���}�-:*�Hz=,�<��g�_m��UGd�)�Мɟ!Ff�͛2���&�9�X�46.\��`�Y�V��2������&g�p �=T0���N��9��K�T=�49u\��ŷ�+��G�d�i�bk���K?�C	���������N=�8r^�qD�x���#���X��СCtj����̱���޼yk|b��s�j�_[_�3X��w�"�99I!�&�&66����?���:<24159??7}�h�ZҞ�v��~�Z���-,-ݸu�̹s��fff޽|�ڍ� �:<226���x��._�6::^k4�R9l4�A87�0s�Xuh���������N�������ux���s���L��������!o�x�?H7"�W�.Ŗpk����8�w�TVet���E��5zp�������nݺ�?�����_�յ�W���0�:����B�4����m$���ZI|]�p�Q�&������7�HT�*O��&�{�Y�( ��&d��=�̔��U~�N'.=qneT�z�D�)��	�Ȝ�Ҽ���M���UM�k��2j�\���W��$���敡9OI�K/nXH���OL2	�B���@�� �;$|�#��8X�l
m�K#-�URcª8�@�=������)��l�`[J�"Ju����9��/�'~�' A�{�%
Z �T�S!J,g�T���2�S�M��YV�$�4Z���+Z܎�L%Ѣͦ�QLߚ��Iod$�t�ъXs�t���=���Xͷ;(�]<re�_��,j��I�؎c�t+�{�I8xJO��,d����ݵ�{��L�]�O��d����W��.kOy̪���yEuf7����z�Y��U����%��h����aﱔv��6���xezz�avv�NMZ[[��9�m��%o�'�2��)vb������ծ�?LLL<���go�y�GD�s���������J�G�/<����ݺm�U{��1`�V 5^�p�����DԎ�?�S?%g�>�O ���pT���W��5P�w�8I4����w)��x�ѣGG�ǟ@oxO�?y�С�������� @�ƍ�p4mlb�����
WWW��oM�I�osݎ�6�H���N���F4��!�*��+�c'N�	����g����/��[������������r���A1��Ѧ��S8⦙jF�ҙ5hs�0�#7!���s[���A�s��R5�t1y����yƔu���.9��	������F��]QҔ^���'��){q��鄤)�5��L}���ך#b�=arP"bb�V�H�#�vǃi�G5��2}��c1W+�D�������pHH���V�	\��.��t=ۜ�H٦�2�+q��OGؾ E��/�%����${z
����=��YXp����Σ�������믾6L��O�[*xAPx?��+&���kECf�����@������H����;wnc�I�r�@Y�mqF�� Ư�L�jyED<���Bd�TFN��@[�����e������)^�Z'#��$3	3�x�gz�ݨ|u����NAl���eS�r&4{��f��ud�i����w�R�������?2˼�oѮ3-#`�76�Mc����E�P���Is�<�,�43�,��I�I��u���1��l��O�=u��c�v�����+�+e �m�\ ~��B�r�sO�8.�T�aa�o# ������;;tY	�@~aV�E���Y�&'A��ݻC##Gff^��Pԗ����/�S=~��nmnoݼ}krr�I��peu�%��?�Q�������믿������,N#�: tnnn�eG��t)_{�s���S�O����mnm��V�ܻ�*h��_�ã�P;�'��8�	�����ҥKx-�s��%���	�E����v�
�WX�� �����j�����VMr�vU�Ѧ0p�2˨7!:�&�rUXoԫVn�?����~�����}��v�Q���Q�>�CZ���!O
/�W`[�$�+���1��$���5�����x�g�V*���%��b�$�L���5�_z/�����_�k9�M����-�Yԍ�PcW��+e�f�$1bÏ�+��]���B�7ve�6����V��T�������κ��(&5��.Ya`X�R�a�,�f�͟��� �8b�@��"���
>�s�����G
ĸ����H?A ��޽{ЮN�8!>�l?K��KM�t�������#t����EI]XX � o#����n�e�L3�y5He�Q��O���l]x� o�o'n%R��}q��#Wr� �R��H�����O��i���cLf'Q6K�1Һ�tgB����O4�.�dm��+$���̗]Ӯ��|;���SH��o�y�Q�
�)JQ�	��I:l�l6y�z�b�z�����e�	������ѣG�����w(��8�r(Z��
�<q괰Mp?20(��!��R;������<|��+�����x�	�	X�wϟ?/T}�ӟ;������?������O|��W_EC���WW��_��8;;��3�H�6����8�9H�é�)��#��KK�	P�z~~����_��׿V��I���<ym|���F�$+A�ݻwgff@r��)�P2���>��7n���; Rd޽r�ʩS�����/`��m_2n5�#L����q��Q ة�˲L����.S�ޖ�t]�J�f��N�����σ6��ym�}�]�sD�tmcÒ�)q`救���6�җd.	
��N|oM|ہc]���f�C,{	�ݖjF_JxW�=�X�,m�O�h���N>D���a�{�����ś�u��k[�-�Ōl�R�؝&ߒ.���:����j��x}^�m��V�Ӭ��!�w�\�z�=w��.�e�˛�t��C�u��%ކ���[���V��y� ���J���+�B�:-�h�-��><�)O��l�ǀ1vs4�4�E&�x+?D:�ݣq����(��Х%���+�_�-2�����R�|�رv'�q����̋3Ӈ����{��{���.\�v���6�W�^ů�����t��-E%������D�ܜ�v�s���]@�o�����%��k;�Y�4�m.h�:���Ke�I�(.7��[X�G|*�;Aֈ��N��m���	ϩ�k���f
��@��-�s��h��V._"�:�D��M`=��k$Vk,���S^�ǫ#�**��,�k�o-�c�f�
ٮv�$��Nv̝��ńH�߽Q��ybS�ބ�C+��'�H<���a� �ֿcLkq�-�����Ϙ�&n�̅8�2{G�j��*�P�#y�l7�&��Qr�^�r)�E�U[&&��Y��5�!rٯ��7��CC]�I�Y\��a���4P�F����;+Ӭ6�b�05�-���9#eX���w���M`�!Ve�jGNP�ʤ��R�&��N��1��9~B���Aˡ�Z�hUv\5>>���y�������6�DD��I_��(<�y�& �_�n^_[;~�h����y	彲�����'!��W�s����D���G�W���N�|bz�䥷/�~Z������863��s��wv��C������O���ӏ=�����R�>~���'�N¥U����ҙ��v"����9����ȱ�ǿ�����%
F�m(�!�T~��7n߹32�ll�|����]mw�+����j����嫗	A�I�\Y��zk�ޜ��@� b�굥����ͱ��}���r�̙S�)Fڵ���������(������E/���j�]���k���Vc�2u���}�����gά��9|���ѵ-%���k���P���N�f�協��<�{hj����3s/��&P#�0�w�F��1dt����"W�6Q��Rq��0���)�\3��N(]�x�dRu���>�K��ì�Ӭe�����7�v��kUUQE9�W*7���0�՞�*����a÷��X�+G��y���	9��eA3����U�Þ�B�2ӤD���Ͻ<Y:�O�X�i�}��^�
�ܖ�>��u�B�Y�3[�g9EJ�v#C�D�
�5�]�.y�w��5��<)�0�:���z����.u�0�Bֽ��Z�qtG	�/v5��/����������mnlq���5�L+++ ��#ƑILC���D��J ф7{��7�4"S_Y�@�-ux�6H�|�\"�QĎ�+*2�j��!�5UX��N�B���C�O�	���:5��!K�ZU�Q����lR�KF��������*i�h�W	g_��G�lg#�af�R'�/9�d9���6�i�Y��[��s�a2���Ɉ����dY'F�HǸ�|q�qe'F��n���s��0C�>�E��0��ƅy쇎����^�qA'�N��!z�\SSWWW�"E�ucoTq�B�V��?)G�Q����~�+K��_C��Oh�X�sssPh��)���EΙ���������Q �\6�Q�Ց9Ɏ�ggg��䋨�k_���?�q��^�~�X�:<ܪ��޽+n!U>y��}� ��vj��;m�� �2�ť�I��`l������i�����Q0����?����ԧ@��W�w�)~`5����ðh ���~tT�B���A9X����I�b��r��j�uxT�  5�,p��%�?��O�����?���K�f���SS$�4�����Z'�,b�h5[��£��ak��"v2��Y�AϮ�����c�i�#�����ˢpz-�� ���P��Q2h,J��F�������0[a��?I�͹��L�厄?asF���я,ڍm�*����R������:*é����/ƷYċ5.�l
��S���7U���_���$
�D(W�� ��	�+��BB9۝�G��9*�:T�y뺜H�ŋ��l�ɖ��E�m�#�7�P"Z�]��í��w߻�\��E���1IǍo^Sf����Kbӎ'�eud�u��t".���y�w�>oA�ݪ�V��ɬ�@���Qfz�Ѽ����mF�6�Ht&M*�G(�#K��b�SGz��)8XC:����gONs]��s	EDFH���o6Yj���@8�U~גgUXL��}I�Ȅ����6EL���#���h���x9F�z�bT��e:����<�z���Qb��V��n6�cw�}�^����>(ͦ�'ϳ���X�s�+��&�aD�(�!����?���Ç�x�۷o��  �H(��X�"ْ��K�X<�|	7����J�`����b�u�J��J��� ��*C�v �A18B�h��hӴ�6�-�7�p�����흫7om���ͭN;�9u�����ꖖW_xa�Z.���[vd�X������6t���Y��(�~�����F5[�1V�[��|��x4A������g�yf���𛳷��� ����~`|lf�p�����@EC##�&-�F�>1q�^��|���X� �>]��nm�tZ�?�Ŀ�no�Ie�T�KޘD�u�2�)/�!��4�����/��/����gήnpD�F��\+��#b��Bݡ����gKDlF����I(J�(�1\�^2]&�x1"짲Z\+��@�`.s�N|dJ����])$Q�e���/�[�!���z`n۟,`&k�uk�W(�֦9�Π�1��0ٺ;�*�u�@d��tz/�a~�j)P�d=�a긇�gBy��hD�O`������K���&�j~�b�u�a1��.�eʎ����@{��&A��m���{ ���|�ܹs��gddT�ۂ��m��js����=@&l�<�+�g䊹�b�"J����V����#���=X=�ξ}!�Hl¢�z���E!^&*�7��@�$�$h��E1���� ����|��$W�sr�{&��Xh�y�>�%��L��d���l�'>A�ݬ�Е����F�F�)��S(��pXsP����>�q�ӓ���<��{��?��lV�Wta9�9��!�LH*�	ۅ�%&�xb�n�/�y뭷������(�V�-��bb�8�Ζ�9`�?x��N����S��(��O����`r���iO�8��L N	��'���7�ԕ+W� ~���H677��A��ʢ�b<�<?���F��{� Sĺ&\YX�����,X��hO��P#���h�5Ks����t|�;�y�����o�����;���I��~�^�ç��?����fK�a�v�))6\I�L�y	�F'�����i��%A0�Z���w�ʢ��9B�69O���ʕ
� )~�K_�v����?~o�)��d9�Z9��vμ��bĮ���Hvk�Ė�����n��xA����(�|ѩ�{���9վ�g��maz�A��� �2R3�z3P�<���7+�#n�Ч�J�@�pf��<��C��n7�y�1������b �Z�(�g�:MH��^�&���1�2��챴��NWb�7� �L��Nn ����!D�7�6������`�_��	q<�����p �NZ�N�-��Y}��f���2dfA!�ɋ�~���l��О��b��-P�q�b'Ȭ��?=0��,�oZ�#-gx�щ�0p���{C�R���.�O�L2l�`��l�EH�~E�0���^b�)��Vnw&������� R$k�f[��n'��8�x�݋�ĥ$v�Ua����69a@���IꙎ���N��HN@�Ac%� �J
7Yʴ�u��݆0�rTZ���}�$�~n�ؖ��X���!9?�ⓕ	��R��C���43ԙ�L�ő�81mT����:����܏���������ʒv[dW7�\9~�䥷���w^~m6邦�O����W�h��R��JU��!`��lxt�hd��;qO�x�snn��h?�'���ӧ��6�k'O�<=~��ŋ�i�//��s���������Y����hgg���]XZ�y�ΩS����v�}�2J~�0�4��]Et�aM�E���Z�v Xr@ѕ�-�^Ĵk4�ZQ�ו�UP5V)�̵������T���u�|������Ņ�g�D�O<q�? ,�e*�8�𖵭mLT<o��f///�,/>��S�_��f����������nl����}�ݷ�~�����/`��./cd<��Bu䛤��G}��?���J�3G����,K���O�8�����(�d0�+&Os͗J�
�ٝuN�8f,�]������	5/Faj�N`�9q��S�[N�|i�[�[\ ļ����6{��2��F�F��1Maʀ3�n�-�mѢr��)�nDӒ���JF"�pmJ˰0����CosPE�v{$~Q�D��,?�> ��h��8�r�����F��6QEm��%799)��0���������jЧ>�<ʄ
��+� ��Ep.�uM����D��v~�lh�(�^d�8d����o�	u�Z-������RU����O #�x�Ur�5!ƞ6ŐZ��Uv�;|�Az�'�^_���j!��q<^̲�SVO5J����g9��>k�y�R�<�3��5���v��
�e%}_�º�2���\U&4!>�z	���nL��̌q^�)E�����)��d�n��c���B��gI�y�C��)�d��<r����r�&p�-fȴW�W_&�ʱe[��T6�W��\�44�c�?~|i�d��#�j�i��
'('����Bk�����~E"���O�T��N|O� D�++@நq�8, �y�ǐ�Ν;kk3���� ���Ƙ<<��3� Z�ʊ���ҥKx]Γ^�v�����6�`vv�����dr�\����/��G�ye����`�x��Rڴk$&1���N��iAs�זּ�\%�Ѡ6;v��-�ӪQ�,��AKѐ��z��w~�w�������zݯ���R:I:2�z�߿����㼷���W�Pw�8��,�rma�f����mG�G�#��_�_��ׯ~���N��}M\�u9f�&b��
�>qrs�Q0��d���݅�s&�lf&�O�R��8�O��'[^�ȋ�@|ֵ�F��ǯҫuO<�K^���km�G�n�U�k�(�)����}3"s�L�G+Ui����Y���
 ��YǺ7I� q�䃹��6���	)dg㩛*�%�ڦ�Ud��G���Ƕ��\فU4??����K��@���'�� i�j6�~�\�<{�������K�*�[���qd���0�J��( rC0�!x͟��B���	�����+%����+فe��1@�v:�p�gԝ����SZ�'${h��{�O���	�:t�Sw��n�\�m&\m$gW��>g}�N���z�w��f�ѩZ�v�{$0��d<du:>`mF$��9�{�<��Ob��ӥ����s�x��(��'1�&��u����M���b������K��y�4jtW:w(x1"''>���]4�Q�k��o�l����Z�)\��`�I��R��cW�,˜��
՞�Χ�?�a���]��$���_���VWH��א��*F� "�|�[\�5[5_5��!R_ɴ����8F<��E�E-CC��_%�/��U�5:j&;w��{��c�/O?��ٳg�4�olol�LV�˛;�����������#hC�Z�m��bkxx ��<E ��ʎ�3�W�\�C��\z������?��+W�,,,����}��ɓ�q���o�:u�Oc-����76>>�@paaN��O<xp��l��Z]�i5�5���@l7n�^^��XSg�R����ӵ���%����������0�E�AG٢��jmA���C���ب���	�KJo�q� �K������?6��]}����n��8����!���b053�����h�[7N�8�y%c�P��M�H�n��vl6cy��?W�ګDbs�S��Wy[b�3��N�b@g��J�~l�׉y+J�Ww�9�X�,4�Ǌ�e���o�-m Y�"���F"v��Z�0�N��
��L��7�Ε��i��6��Jƙ]�W�z$���󸻓�oA�:-h��E�3Z�ӛ-	�R�1�3	W���+M'��YA���~1��ᙙ��_}l�Nt���{��JQ��{_�Je�]��g����2:2��q*��^{�^��`E��a˶�@��U�-�'�K�|r�
�l�����Yj�ݙ*D����Y@��R3Ey�#`IQݜ�e�Π�]gu>��K\Z�?���2�_dL�O�a�H�P���=4I��=cFk�,g-��mK�ұ�	��|�m�i�4P���U��Q�1�zM�H�=?v&��:&f�A9arP&��31-�ԣA`���Y�jK�7�?ڽ��w�*�^��9�^G����$Q�`���N�I�O�* ,�x9���Hv��sy(��
Kͻ�X��@yH�c���x���c�C�s`s�bq�ns��Ol�1���[D���������;＃�t�_7)��hgii	P��w�Y�K׮]���~�	�/<�4�$^?w�ܯ�ʯ���������j��_�����'�ʮ�/U@��m@E��I ��7n�;?�lz������T�d�i��O�����/���s�=���R*U8 E�Ӗ�*�ܶ���;8�>Ǩ�����l���_����͛7o=�	��u�D��:v+�ӟ��������R�onG�.��d{OI%��ql�{t��鲿!��D<S�X!��W�WϞ�qmV��:2;?{�O{b�P�iӉ������rәu3�J���c��PJ)6+)kq�,1�"�<��^����y�!��Y\o7hE�8�Sķ�Dg�βDp�}y`[���T؂�߬�x���B+��U��"��$��>�Ȏ�j�)3L8���� 3,*p��G�b�#'�V�ݻw[�"��9�"�9�"W\�p���ӧ���!�[o]*��tgh�&�1����cE����O���������޻|yiq��@A�ppfL{���f��'O\�v��Qk�u>�@$�v�'-=N7%8N+��X��6{��A/PY�؍l��>�.����ԭ��,�?�.�o��-��-tZ;��1�^"Swۛzm���֙���?e�Vis�J/{���ѫ�.:3�KUb��%ƃ��C,�y�q�9ǐ+�K�F�FQy�q���g��v�	:���i6:�.]��E�����B+ڂ������BN��xp��db�ŭ����?���d���i�|X8U��a^��I̛��%�%9B�ۄ�H������
廬�)�0�㓙%/�.L�)#K�L_���U{Y�I�^���lr(��kB�U�5��QZE��[>�d��gf�!LY N|�=b�;�Dl9�3�$J�N;l��� �2n O�8�?I%�b�?~��^\XZ~���olI�!
�
ͰR�;�ds^6� �j�Ʃ������|�u6�J�X]��%���q�2�R����=~l}sciy%Ҏ_�=~�+uBg��X�U���2sr�2<DK�/�mλ977'm�V�W�7���|�I	����`����_�����{�w����Ǘ�_������� ������~�s�9`Τ�)��d%�V��,yf呭�4�g��V+������X�Mɦ�d�i�b	�  �Ј�@���/�����Su�}� (�l}��ի�u�s��Ϲ'�v&�:�Iq,j�u������.F�񆌈�K�H���`�&������0���N�w�m�����{��ŋFGƳ��t�P*�UF	�K�!G�x�a�Ν>9 �-���/�Nuu�,Y���sgO��wl����ӧ��P$li�_u��v� ����bQ��R*i�CN�ilm^�|)�H�=)�d� z;����\B����ZeP�x3�����mϟ�C����BEK&u���L��R͡�����xb���Y��V�oT���hqtuR=��|�&q�5}�3�%ڴ��T���~��\�[/���S�8�.�ĲqK�	�R"�(�D�un�US��]�Q���n�lx��p��I	���jл�Ǩ��5"pA��$�}(z� �4�3H(Ω*I7
�z;$>�d�nn��CPt�-[&�k���V�<�phՈ3�O� �;x� Db�3�	dL��c?����VJϝ�J��|�p�l�JyS<��.C�`�����.w@_�J�h�|�	��9g�n���8˳{J�����/	��?���CQo�+$�/"�e����B�b��=55���M�6gRpGe���
V�T�GUn���x{f{��r*)vva(���$�
Z^�INs�E��je��*�Oy���(e�X��q���*}�bP�3Cc�jp�7h�ժ���c��G]?d�s7҄�U@LɖEP�E�_�"+�JKE(Q�	�R����_e�g��&���c�u�P�Ξ=��Y
0$��U� D�a.�D��1Cː��rrr4,)�'N�FW%�~����%	P
�,��?D���sow>�O��)Wo����p���߿k�.���]{���<����Й3�>�f�Z4E���3��
b��A[��,Zv�-<��q���U$;���p�u7n�L ݆¦Q��Ĳ� �P���(��Ǳ�Qх|�-iI��)�b���7���'�2����k2��5'N�8p��o��o`�N�:e,t����x.��/b�d�G�W��,����g��T'?呦lou����*qd�S]h\VEߌ9���.�:�G���窽�N_�ܩ`x����X*d�fLjQ�-+)9�m��3��,e��@͟#O�����0���?H[���86o̪��%x�K��n�Y����B�2:ɣ�.������
�.'$(RL�zg���N�F�|�
��l�Z��:z�(4�x<&�n�Y;V{��UP��j�:�`/Ik���vzjBb}�q���U<)泹i��k�����h�]���q������U�V��ѱs�/�$&�!�*�QߙI��]�����d?5�#��2�;A������%�������\Σ(��%��ꡃ���e>�<.�nD`�Q-�ʌ\�x��5�����v�0dy;���7@Y\��v/S�39���ϕ�7��cYjkA7���l�Űi�'�c������6<V�,R�F�m�:���z2"g�D��� ��zr/�*_�dKPy�8����:��Y�͙,r�����2M�R#�~��S�<m�Z|����ߋ����eVj�
 �s>��B�y���'GK1*������_Bfq�F�Y0�v��Q��C�e�/��;��
�HN�d��CM�F���cΟ?�uw�B0�8�hѢ���DbLj�ht9�Jer�Bѵ��'@唔�.546��OB����j^2��BA����@�x:��ї��as��U� �2����W_}�;n����NGG�C�{_fvP`Pfǎ��/?�4oh�4�&X�R�Dr6�c�B͑��/^��=|�Ț5��v�ܙ����L�d��@	��ȃ>�d�RpR:��E�s���q�J�	H�+0"\����~��m===��}�5{{%Mnck��e+0�',�Eb��_�����w���Բ���w�qq��}{�J�*�<x'� ���K7YI)�_,�29����k@���W\&,�	x�]	ΔYA��:��_kAU]�\�yzHm&3�&Q�PW����e�5�gu{��Te�2��1�J�ְ�W�U���NsK���B��Lee̪�W�GuRA���cF��*QW�,u�o���q )%5�d�'!n���ڛ���-$owI�CM?{�b�g����'�r5��j���Q�y�k�կ��rՔ�KQ��xLr*���FVh�˶4����n$D�Ԇ!�O�V�7lX�|����qe�װl�|8$O)�-T9�i�6sQ�Y��L���c=�65Pvot���涣��w8��o3�b��k-ٿ}p��tT�0���C������hi�C6�A���Jf��d��N��ҩѨ�4�o�e��T�t)�R�H�ġ1QL_DJ+3�5z��$�CFXP���U���EJ���qYo^1�%��ڎ���B}Q1��d%0�@��щY�Dծv�T�����2Y!!��Pv���?;hF�­���E-�!#2���%S�2��b���KD�E�����ٙJ�J�'܅h��xE�\|M$��)R�E�@�~"����-݀�����l�g<���E�!�~˭@6�3���?~ظq�?���{�1`���%���?�a<���^ڷo_{{��!�C���_��ee),R�*x ��9����������kS��w�>p`�a��H�����ܶm�G>�}�cmmmXcr��O��*g9�fsk�8��l6MU��"i�-X�������ǽ�DB���z���č �T/�v1� ĘF�H~ H���i����QV��b�j�����ee�|&�U����*�zz]6�x��K�
r>�U������{)���~j�C���J������˩�T��((jz��:6�ڱ���D-?̕����,�#�����ۭt?,�װ��G�E�X���oÆR�ܹs�i,7A�(��O?���;$I�Q��e�%Y� ` 蚔�'���c^���cj����^jT��lE�l>�G �f,wllTHTRoc���l@=b�;^��Ĵ�9rϟ�x���Mk֬�2�ީ�E�=3�҉3(|E6c����N3��"��c�X�~�(�U	��c�P0$�%�5ͭ-�x�;���o9a3�R?�vȜ����R;3Px�"�J���0�-ɓJsR���������'�yz�S��� ]eQB"��l�t�<y7/l첝 �Z4@?6���)-K�Y�f3Qٻ�`�@l�*{P�)��F�3�%�CR�iX��FJ(W�4yhF�;]�c�d�2�L��7-�q�r$d,`J4_��v�5D�V̿������Ġ�^W1}��B��j/������1�1�ҥ�pU�u�V����I�g�35�e�f$��X�Hi����!������g����?[��M�m�/>~���� )C*�D�Y�q{"A�L�=FF΃JK󪫮B�###��ɴl��c�' #�X�������n�:7�F@����x#��L������\w�ʕSmS�	Y�dr@E��r��ի�����\�ԩA�3<��^��׿��/~RbC^�d�]w�q��)�d�D?ņ�\��d�����T��L8ܻw/� ���Ћ�=���|����ff&0Ɨ_~���>G��ld�[���<�P�Zr���|L��N�}nlr���j*��!���^���d��e�X|Ϟ=��M�Æ����޶��ek�=���'N�����_�a6�<>x���=��x���Wnڴ��s��b�������LΜo��n�4^a!3���5��1�z��G���A9&��*i
���^�:���
������M�GSf���=E3�U�M�wR��Z}�����zU��1��R�C}u��X��)]tK���C���pUs]�He�V8�i1��LFE����˭�^n*w}�~�/� X�I�f�S���ԩS�h�j9��z��)�N�S�Q'9W���A$I)��/�K�&!6��L��iՂ�ϕ���G!)�&�S���rh'�]nM�	J%S3�S��Fzzpzy�д��B�@hb�Y��5�Xbt[����^�pxo�&`��D~�RrFO
�$OZ���Y]�tߺ	M'o}ݪj_Goo������*XEt>(�%���)g:�*r��eȜ�R\)�[Y\��Gr�ST�q��ׇP��jP�1��#|�Gt^�m�����f�����)�(���гE�L�gF=Ix�G��\��x���m�k�i�I�vV��ܱ
������H��|Tj���W��	�ܺˋ��:u��l�$�t�W`G�,���?�U�"�ܙSO1�b�W�Tb�`�Z���Z��ah��V�Ӡv�:�*�UD�B��D���#dZK��޽ۡ��! !t��jٲe@9O>�$���֭[�`���x

�L !�RQI{��(b��8����?��](�'IW�����< (����܇m۶}׮���f��o�wt�s�P4Z�f!6=�8qS���h{��;W.@�9Y��Ս�>{O��LbNV�XQH�!�),�koo�T`�O����;��_�u��+%�`g�R���S�4+�"*m���� &3v�[�L.E��]F�T!YR=}���:<�g��F��n��:�il��O�g���L���� ]�	��t�Q���R���)վQ�J�WN����ew1���l/�_�c����CIi_B���TS�tb`		#��#2��D{؜�5)��ū�Ma)��ҌL��71>:<t��7��58&���-���XFu��]�ϦW��c������L1�1��q�[�˦�Y��䦚��$��̥3�hw��k�抹cǎ�;wft�B*���Bh>g�O���i�M5/�"F����M�0󹌤���k������-)�U_k���l����k��D�⪞U��*�8	m �СC(!���Ta�!"ީ��g�H��� 6R �a���d|�-8ݏ<�#7�K�e��jT��^ì�ɋ/.��,RD�^�?i��?X���;�ĪK��t�}}��c!,��lG�>]ӯ>���66a�U���Hk.+�C���E_"��Y�tp�2ky_���^�Q\
�Tט~]���\�RB �j�&)Ʀ��0�K�V}N���zB��ɉ�f��KK$r��"c��<]LK�n���� �K�@-X^$S+�kh�[����S4����OD�nJ?$6tK.pgWe���b�.��&Ǜ��$ia��. ��Ǐ�
���e��2w�}�/����oڴ��ѣ��hC ���F��4�ӳ�P��~���L�..���u���w�umg``������ö��=��C���?������G}�C>�����?G�;6����K�������3x�$0Y�P:v�xkK�7�����F�W�\��Ԓ��n�
�u�W�|���w�vdu�p gq1%��Ezz�<,SQ�UTQ�v���dϲ@Z��ofՒ�:$��reu��,/��݋T������J��4��^E�9���Tar�?�>��٪��}0�Yj^#~zqSW}��L�z{U�Q5������D���Ν��c���'K�?��.Ԇ�����&�-t/vDKC:��!�QLr6Z�(=��v�rr8���?	�&K���^]rG���2�seG�������H��Kt>�X�"Qa'�&3��
�KJ�>sP��~� 1���V,\�p��6l8v��]w����6o���A�R����,���&SM�J��VZ �7(�˒�.�W�ϐ\mmmn�KȌQ8��R�pX���.���K9�^'EU�S�&��9�D��܇�r!�=`���; ʆ�(�>m�dK�٠�KX~��*�?X���0�=hC# �{oс�s�5�R/W�5�+����:`H�j!�^�ስPe���d�dj.2��_nJ�ݿ~�~�G��7jH�� ��ѵz�j_$�H�l6-���3�Hr�G��E2�,�Pխ �):��X��,Vp�H��̬DSBh�+� d1�_Y99&7(�R���#�E�kW&���)�1��l&���-�[p;.��Z�l.8~�hoo�M7���ĉ�/������S��,^&�m�r���=Z ��p�2۷o��Cj� J'��0R�B�*��-�%BR�)�%"|$��0Tf*��`�r<�� ���8a��O~�i���?���<��«V�¸$桹��˴�$	��	,1�����$��#&y������-G��5D��˖-����Ȯ]�*�ܹ���kp/���Jq�L��HE�{}�g~u^�@�\��g���#4^�^��a�m�ꦿ�d���lD�[��zG�	�E�b��6�c��e���%��z�谪�Wﰴ�S�9UCS{�Ϩ�_u�Y�Yg��W��L��^n	S�l[�,cF(q�)ÆN�b~�KI�#��O��OBF�N1h�%��He��ӅIC�Vq�jY�|�P�\�/R�M֧�6S�H��ؽ��A�@8VHqT�(g�\�Ȍ�@`E��-e����qd9�"qYA|������9�TrJ\' �r)�D"%�����GGzz�F�Ɗ���ǚ��TF��%��v� �����Lf �o�=�a����8�X8T���˓s@C�!jhnm�@��v�<��6��l�����g
���������ѝd��%K�[���;�ܶm����{���Shnn���j����U��Ԯ�7e�kQ���1��,��gLq9B�U��2��X�E'���ԓ%�����R�OinE������d�����l�7}�,i<8������K�xk����gubt�o����s8��!���H8k�*R��u��ab!����~����L���
�ki��6�F#�t�1�X��TH��uE�T(�(6�Ñ�k�&6��c��\SQMN�e�e��	M�??U2�;l߄�*�E��vtK@����Y�u[W���	�,ռ9N<��d�{�ҥ���Xqgg�J���uLr4�baa(�����y�ť$LbYw=�!��?ǭ5-�V�\�j�>^�Io��5ƕ}[~��٤���	m�W�O8���p���[ߙX,ןDi'�%L�R���.��8`0br�hec&��B��R�881>e�Ʀem2u�S�Q���k|�B!��K�0/бp���9��JG���'''��P��h4��n���B�(� ��u���9{�,ջ+����8H[k��.I�L&(�D(��b(�@����ƞ���JZ6;�y��鞮Ϋ��424<~a���`ldx$�MM�O��z�Y����ѝӧO��-�<o��NM'�'�`��w�^)�gq��-�3ѐl�3��ZV�� 年���UA�`8J��R4�C��Z��u��z�>�����v�9u��7с~��w�q�W��կ|����ַ��ZU�d"�����n*�Xt9!��?�)����M&0�gΜ�2-
# 6M����	m�]����ebfrf��hů��s���wv����v�������Qm�:%���͠�Ub�Ju��z��X,bAM�@��iu%�1[ׅG@ 6�V�6�i(���[*���2��A�T*��#� ҼT����Q�$��I]��%Q��2�����#J���}k�뗥Q{�6oby�F�V*�0���Rm���g.[E{���?^}5*��LQ,����Ю��
ꊉ.����Rѳ
u����U����r�Ԗ�|����z���7�%~�x�d|���qpVI�����q�g���\nӦho?9�&񡎟�J���:��1�ڊ���P�n�}N>S.o�sJ���-3(�����>*�n�~�*���B�]�Fʌr8��d��8�ix�����6/�:�P��1�o�"� �$�j��%���s����*�zt�Q�`*l?u;y��e^Jn�k�j��>p�����X ��={��<�J3eH2-�U���W�őӌCI2�az�2(%��9QLgT�]��
�s���y�)d��.zx[��B���eǎ�Ν[�b��� (�R�q)h־��I�#&��`�w�V��E��%X����>��i������p��49,@�7$�x�%蘍�P^kQ %'�]�J�p��)Bj�?'L��d;E\���%qQ��R�RR+�[�����ҭ�
d�*;�T�eH��"Dî� ?���%�Ν;{{{Ń%�L�Ϝ8�H�ϕR�h-�*�EHH>sW5�*������e$�^��6=3��X���om*J(�_{{[h�������Boo��LB�O�����1- Q	Y@�V�X�������p,V�g�zz�:�����Kߤ|�C��ߑ#G�����A<�����կ~u�8��ʦ3�}��篹�Z�r�����<v����h�o���e]p�N$"	jE��U'��C�4c(/R�Y��QL�:-Ԋ��.�^�)�g�φ�dsd_�x
[ׂ��b[�r������9_lI��Q.�m�ߓ��T;��(��L��R��.@��D���]��E����?���i?7���̂�%�L���pd4Θk��J�ɟ�R6��F��V-_�j�0�hdd�����������s�=G���;����E?-gA�Ʃ,	��c���d	���K	SV׼J�Bi�?��}����
764��)�k���)�CH�}��a�ׯ_��_�d��lvl�b�0. Eq��^�X;��N�D�EJv�ʑn��ˡ������'ڋ��w�k=�����D������,CoF?�N�����PL�)TbY�.�KzCGG|6�=9xvbrj����#��_ ���S�p ȥ��q�� �F0���J!��:{(�ĪU��Hq��'�K@j.$g�u���zp��"�k;u&�K����O�<}axdp����%���.$�m��݉4#)+D3V�Z6:fEL�[Շy{Xsk��y�_�b�����j��n�ǹ_MoZ^�m��R1�sI,��5��x�.���D�dO���JĺK9OH& ʈS���@`h���R�&��Ȳ���L�sI&g�ٴ왊[*;rQ]#��,�-
�ݗ_:�������fe��UNO'��ݥ:HE◂����@������&���X�5��lf�ۥR�
x�d�D�%���0�h6������'&f�"gϷ��Y�Jř����L._�5�������y�� �x��l6��M�R��&�o�y˖W�n�p�v���G_۵g��խ͆mshBJ4.Z���(^��C,7RK���ӳ8�:{�,x����\�l��{�%�鞾��-�O��I�I��U-�;;R	ھU"V�2o��E��ЙZ���ҭSҎ�W�����z.9S��V�Q�
�:E�����Wk5s-��<J�t�.�� U�K],~A����0��{���I��j'/CU5����蘗�TY�v��-=�Σ}o3�3�8���=��*QF~>U�
��O6	e�H� �[��ˑ��Fb�xZ��'�7�t��u�6l�`�7�������_��8��#����(�?b*3x��!ن�{|�֠`5~y�0$
�^R^��S���� C������%�p�s��y�3�Lg�}}}��r0���+�>8����=��q�ZG{�����.zs�p���WKl>�xDo3���d�Vj��C����Kf�	+ڬ��� ��<$�V
�O������r� 9p@.oݺudt6Ż�>�'K0`����S �F������Q���Oq�<�����z.#u獯��&q�Q�L�ޣ~������% �S�'���k��������I6Q�9S/��
[�+S]�HVs�.u����5�f��i�"H�SW^,�]��)U~E��{ߜO�_�N�[ &���0JI�@p�1�h@�K�.�� �"ɩ| -3�:�� ��� ��<�l�L	E'��A�ai���Y*G�K��ѣG�[�In=	��9�$G���W���X�pR�P1"tF<�. 	����W`J���/@O��ɩwtb�M�!�q#f �2�]�\�|�aR^7�3٣�4������b�8}���ŋ1�?��?��m:���#s���q��~�D�#c³hO?�B��	U'��&�7��N�B��6o~	,��߷�\���9r����L2ó��t������UP�"����*RT��}�\�P���ڕ�iNr}Y�sA�ch��Z���U��#��v�:>+ߠ,��
��^]�����r�h�y�*�*��e��Ϯ ��VJ]z�sx[ֵ:"Oq `���p ��rMF�g���ڎzJ%D�ٵ���o,�x��JnP��EB�P�X֜��M���%<�r��5�\&ΰ��C�q=��+���СC������Hf����3H���Դ�_�:��~�D::��e1�>��g�� T��)t�n�����d�G{k+N���o�y���������K��l��J�t1:��
�c66ė,F;p���Ęc[E
�(�	@P�RX���?� �`��j����`���l򊉻Po�(\3�ۭr	3��YS�j���U�U5�U��.�qh6!�A�6y/�d�]�h�K�i45u@Ԟ=wr���3�/����h���H;��C�(�h�NOg3���]]BlV0
�CF�Vۂ��@�.��F��,�QM*9U�c'1S����u��)��L`����*}f;�;��b&�',+��油�Dtvr�J �x���'&��wff�l3.)]A�ꕺ����C{��9�L?�V���S�N����U��<����`�W:l=��Y���M�ݪ�(�m�؋T'��R)�Y��)��J�T�!O�)�����4��b���Đ�,yk��&����/h����鑜���J�'&'��`��~^���!6��b٬,<��r��?�0���_2�*	MM32��9��7��4K�"�=��c%������̙3�?o�6n�(˗/���XTn����!��%K�`����[�ft�'N�"Q��R�����{�;22�e��Bu�歃��1�3g��t�u�w�2��,��2�� �I|�?>�gϾ`0�����xc��I�c\�X4��n�2����<yK����{��~��q��3�dGowς>�hI��m۷���e� 75=�U���%13�mnm���I&�@����B����J�E�}��<�\�chr|�a�RB�3�����=B�½m�;�UF'l���ת̷�[�_u��f=߰�nĿ`����Y���J���_[.˯�v���0(�JY�mZ��<�z>�R�1����ͬ�ɬ<���VЇx��Ȭj[M<&g���`��m��=�|���?00 ���c�3����'3��8>�WQ�Ј*|&vrzF�(��y�$<���I��=hi�F�d�g4�΢AJ��>���[�b�]Q�$#�g>�9��p�7����O�]��nD���H��������;���1`8�md8�AV���j�{Ȁ����\|�V���QLQ�LV��s\��0|n�y�m@���4|�ąH��TH�cǏ���#c㬠�c9PBs �p³i��e˖a��*��z���6��p8�x1�E`Z~��J�9�	����qI��2Ĕ�^�A?*䊯3Sgǅ���]�~-4��+WJ�y�[s�Xo�F�r�'|�<��N*UCin���UX�D����}3+����ʯ�U���ޢ��'�W��#1mO���\2X��b���\i����⫥�"K�8%�=;iЖV__���	������Yo>U6��/�e:��0�����v}��\�n�_��_c%����tkkSOOW�`��O��{oii:�����,�2 J��	rA��à"P�ࡾ���ѣ�f�����Lc4
Z:v��M�6ś�ɺ{{��֮]�jժ����ٳ_���a����<��#��(��m­���+�!��e���{�O~�i�_�җ���z��@0�_9���-]�3395Au5� \���+��� ��.\��)/���l�,Z���W_����$�;GB���F������X[�=����F�� �ZQ>l.B*/H���[�D��2��cC�o.'�T�������C�-p.���iݘ�'E�O�Im�ЧOl���˩�V+���u��8X�5G��QFT~jн�I�:�I�'���a9�.�x�[�F h���K��2LU�T'�����}�g��+9Kn�����X����"'<��s���Z&�:u�������ظ��-����}B��@^k���#`��]��خ��)�0��HLl�b9C��QK��\��0*��`����?�:��pr�GƖ-/?���m�|��G�����g��c�IZܶ��/~�w�H%�v����58�b,^�t`dx$�I���|6��Ҝ񟲢�F�b�Fé��b҄Ն��6�8�Ccc�=}���7/�	�=�/��x�8RI�\�{�b�ȑ( k"do��ba8t�8��L��F�y���8�޸�545�i�iin�zs��	���r�
���U�'�Z��
�Φ�Uԫ�Z[�h�&�����yT������.7����I��A��0[�xKK[W&5�L��I�+1=9�H5D��djo����n��f,�����ZL\N�HP9���I�W��Ԝۜ� ��ꂹy'�'���벵^&B��齃�k��d�C�+�8{��+� ��M���|ў�M�J�D�ڄ(!��A�rl ���,�hr#dE%�J"� p���8Ġea+�TCCbjj��͕l	y���g���`��ӰDH���OV�d঵���ˀH���;22�@��BO�L,�X��<KC��]*$g��K[�B 3�#h����An��	����_۽�X*&S��B�����6nX�׿��G@��m�׮�������-MM���?�������������o6������O>96JNo���.�EO�B@�NLO�v��fF7~�������oQC����8C�'==;w��dɒ����(lX ����F�_����m��Ho_��ӧ.Z�D��'[������TN4�"�熢�<B��Y4���\R{z&KL;z�OK��떩�JQ;�_���ӄV�6E8��q�f�
ѵe���hU:O�Tӎ��i�4*2��9��/C�|��M���EM����������嬵eqɛw�Q��U��*���y�~��2}�W\$E��Ff�!�ypp_��[|�A �={�|��߅��]J�t1}8�R$> �N\dp=��8d :*3��W| dQ�3x��;�.��Ƀn���ŋ�<yr�֭gΐX���C���Y���K\��]/���ҥK�z�i~�+_~��o�Ζb�۷Ruv�r�A(r��W\q��p�H��,>����c��g��_dy�+��3�y�CaW��-�I�j��ы�U�Icn3��ċ�q(��z^>š���������Y�C@WE.��<�q��K�{�'*N˙��_�_rb#ɐl�*F�ƞT5����~r~���WA8�f���E!��	&e���@�F�j�+m��y���~�u7ܰv�����ɦ���(�0+�$.�0/m�Bɱ�+����sߺ�
2��(�������2C�j��޲�)�4	���̀Қ��	���yll����̴p�B`)�^���,�F�*�e6���`:�8W�����L�!x��ݽG�EW�n������/�˒ƶ���0p4e��.ޮ�+��""�>�@�nj��\W O�k�rhj�Νh���e͚5�=�<�PU���SH`�ܹsWmڸbŊӧO����%K�}��_�|�;v��k����#�^߿jժ�=��3?������n޼�Y6ƛef��/X�P�����khx����Z�~=u05x'���1"�, �fO/^__�x�v\�����������o```���T�[�Fp���9K현b`���+c��x���y�M���[,����4/�o����ē�l( �ȇ�o���Qqq]�֌W���t�����CaC�^�s�5�/Y՛�}�J1J+ɢ.���J�y�h����P*��zѽK���D�$j8�{2���K.n�D�����iWDQ���Э7���`���]	�	��G�e�	�A�^����!�����d^����- ��Nr4y�d-��T��d���PX -fkg�o�ǧgD)�O�&�-��l���`p�с�e3���`���$�l�OӞ&ęi�]���{��z��
%�w�,�=Gv`�q�R{{+nN����Õ7��w8��	�_ܿo�/����ĉ�|��qJ?�x�@1_pJEӵ�.hnh,f���{7��>���{j�4��P�r�O�2����C�VLz��J�i��<�a�<���#q����&%'��aL�N��m��2*�G��WnJG�8[��ϾVm9�*:SΪj̱;fV��((k�￸?B1��)ryjr�&�r����Ǧ�Ŀ����Œ5LN�onmjk�u�q[���⭭�����¿xE�!#fc�2%3�\�$�Y: �c�c�8��;�J� �Z�J8k�Qu����n�x�z;uQH������i����0TZJ\4nNGG`��7A��씨Z��5��O>��g����۰\�C��lϠaR�h���|9�VS�~�Z�;Ct��!>�U5m\�B�:C���\UM+gJ��j��M֊�:�ڦ=4�gm�#!�%�(���m���$�M�۵%6q#�LM%(E��f�L��9>>1��Քͥ�3�S0x���:;� )d�w4�L)��Y���4��%���c��̙3�ݝ��~�ڳ�5��3��r%�D.�I&ɵ ì��b\���I%�7�p��}�����{�M��|��D�ҩdSc|��G/���b����E����fg7^���,LoG[{4y��������9Ɓ�
��Ǣ���G���P�����믿ԑ7���|��]w���{z����k_��v�ڗ�dm�hj��c��4�'Z��|�����H���7{��+��><���k6�hnm>w�AV��3I�����١��A.����W��E_޺p�ӈLc��8��k��Iph*����li��!�Z\��L!!�Ȅ_�\�u)ٕd�r�xS0��'��C�e̕�t��] �*���f7w\�'ӧjO�׸xʳ$J��1�nU����u�x�⅓v�
@R�g�:� b���k�2V��ٰl-0+2�S)�tYP�&�~����[3�+s/�P�
���-K:���y����V�HՄ�w#b���6��#
������=����׭[�gϞ]�vB#����E�^a����T�v����������=�go�ϖ�J����L���#��G��>�߲��7�<:3�jj��\����XLvpX��߸�r�d/��Z���|��lyT���놛n¤�LMrV�%A�P�M�6a\�)�Ƨd\ί�]�����2�W-����P�Z�b��^�l`^���������:��`h+��Z�K����v e�$�iii޻g?Έ+1+H-�������_@�VJ��k䊮xS���~b}��_%i��̘f%�Ah
����Q�ʶ���yyJ�M��ҹ��[:�.����5C�t,��HAcb߹s����-��r�7N���� ��hKs9ڿ҇Fz��{��,]����Q�X{�|�8G�L.[h��Pp�TG4��
B�t���X����J��N���\R
OMR}L\r�t�MM-�@�T�q&��[�Z ]�R-0�!���{*����?~��w|����;�&��AS^t__$�(��x�Boo��{��r�_�z5�>|x�ڵC�箽�Z�-[� ��ލ7B����I�@:�A���K���g���q1&���x��ŋ�/_.3N�9���W�2�����O���F����������{�'~���ڵ�СCǎ#u(W����%���4��M}��_���'?	L�d���XNL=!;˘.
�?th��r�������L�+D���xQ������-��� �<W��*��0E��p��J[���cn�e8��Ϣb���gs���5[�U,m�"�ŀ�ZfUr���s'K�����7�^�i�zGVt�I�2p�@�n�Ɯ�S3�S(�ӆBfz��1�z^u���<]��\H�CB"8��{�޳�
�l}U.&$}xaN$#6'q�g�^�
`�n w��_�5.0�`Cs%B�d=����K����5\�N�!S�g���ڎ���L�*��#�7��Z��eFi�EN<-Y?�Y��$�Y�?��O \���
2���S�N���a�A��Gɒ�%�L�%�����"�B)�^u����;^<�q�j�1��\bz�����p��hcSkKs8�DBݝ`��8y�ڮ%��>I�:"��.�w�0���;Wr ��$Cs�e��/�x4���*ҝ��:���Ϋj�rI���/r($�|ە7��Ն���}e�3�tGGW���Л�������^n�
'��xK;���ag��mD.�i�j��mq����v�JVss+�.�@(;&ߤ��T��q�-(8ڕ�XQ����91�Eju���ܨ����0�	�K"i���8���0��R��;��s���y��?�g8��r��(h51�J�N$f2ł��5=���|��C�%	�QhO:��oU�ϫ�v-�U눕?�.f��y��Hu�S����Q�p���d�
z��H����W��-�D���0sPFksK8(��v�%t,*�Rb��,g�-�!؞OUcc�HNfEH�~L�/	ʴ���S��������{����;�Z��5R�tks�0z�Й��t:��Mp��ᎎ���[�PЯ}�kS�/��|6�	�XC��>7t��W�LMc,�H&�\����P o����*㼟~뭷n޼pG�;���z I`��)NQ���k8y`���F
�:{2�';^�Ї>�8�o����ۿ�ۀ}���g?���J�̜���=���z��'O�bT�2�1���x�|��V������4��������)�3	���c#��H���2�Bww�0�۶m�o�V�X600r����9�� �h�@��9}�l��C�ܴ�e�nzer�8s^-Ȳ+��h����Y��s�Y2�E!�2���,fo%`�R���\��-�fY�T�ٺ�1�tB��r�}��Rq3�_��[����U6	W9��Z��PΪD�~^��u�K}V�u�'"g��v��S�!��E�֌@��k���=���<Y~�3y7���2�m`` �4���z�����͉�M�I�;F~��<,-��<N�O��b�Qג�:����	��D8r��ppp���_�2��;��Ξ]��p��ȊЄ�9::
�ҿd�iK�<T�[n��=�9�pll�բ���6m��HZ)�m��>�k�������Z�k_�����,>w�>�N�K,k,�j�1�֞�k�k�s��S�V/�սK-ނ3����e(L8v���_>�2�ioiYC&� 4SP�ٰ�֋������6I(��bѢ~��xM�?��󳄋%GlLBQ�|�-ϭ|˫�r�7k�H�ʯ����SW	s�{G�_��]�YL�b�*�j�[�Y��9?y��s�=����{ Fq�L���KezQc���u�5>����F.��.�.���A}��ӗ� T����0-A?�����`���[S�IW�]
��an���r��*S2Ӗt��-�����%&v�f��_?�������l�ވ�$����$�=1���.�uύ�t�G#���@``��n�|��@�Kn<��_4uM�Z��]& �p��k�D۱cZ�뮻��_�շpz2�:�d?���)|���{��?v�UWI�v�ޱc�� $6����+�֭�C,Z�G����|���������&�SSɾ�-�HA��O�����?��c�V��R(�X��*� s�gΜ_�dI6W���8��x��[��.�ݻ�/Z��I��゙��S��\U�GUdVE��W���
s�)�&"HJz�~>�Z�R%�MӬ�G���˽�'���e�_uO �e�zv�J��/�gjLNR�>2�S�Z��Bݑ����3.�.�J�F��9�`2��y.�v�|H&tB*��b������2�
��}��Ӓ�J�+��KǏ^s�U�<���G��`���=�=d���s3� ;�ۆW�0�d��t���"kq�8�5�+,I�3�*i��l,jȲ�_񁀗�Z��&[�1E��a]C����k֬����K�,��͖�f	} b��Nok�ّ���?��G?��@0lqp�5�\S`'���}��W�޴iݚ�XӠ�B56Ĩ�HCF11β,`�"d�B�ӉYL�������(�6$�d�� d+�U<ԫ��Hm��Iz�UJ�b5�U��I�|++���	*R<¡���P�HZi��1���]��+�_|i���nM�u�ʚW(��m�T�A+Ȧ)1�%���N��A��K�����T7����
 �d���RFI1���|da!�e���QN�[��Dg-�p��~�j�~�z�J�V͒Q)�M�:���>��z�^�̒]*�(� �� y�9�U⺜BK&��Cv�JC6�'���Ώ��ŭ�S���y7Pl8���Z��3r��\]EU����ʋ�2í!bo�Ü�������ݟK:L��箟�V�(rT�5��:yIL,_
y�M�RIg�bf����}s����C�4::�  ���G������y�
�$A$a�y��l�g�H�耤����7^��=����W�X
P�&4"��4�Db&}�w����ϸl��-�Fx��m��Y�
�uv�OOO�����xS�����0mа�	`�����=�����,^���?�1�(��$�jjj9{v���2b&3@]���/<���drúunG���d� 0�U*��F����s���O<����q�����\=���@G��Z�z�_����?��o����?8ndff2v��d2�{ϡ?��7�������;�Y*W�Z�w�n�e v��eK�7�[X�r% eWW�/~�L���l*y�M7-]�����l���r.\�������9�]*��*��O6.�����5�����$�\vV#�V���2��ja�)��.��lj�2��4����s]��1�W�Xb�&�J�2/������������g�c���Ǻ"��,zwk��/�q�:���ק�.>�dV����1#��P�e��ů:>��c�غ��"�����I�/����?E�?���~��x�	,A���d,��A��m��Y�Sr5˙��Q��>������|Ӭx/��՗p�//�L�*��$���T�����z��{�����Ν;��>rL��:^RG"@i�����ݻ?��6Fb;I@M����F�>|��'��z�z%U������<�w�b� ���$0�ů�h���؞�����뇶���|�2!%r�[�]T�j�K ����I���2y	� :;��2;���\�54����k#�Q��۶��"oh����|]�tVҚc��ƣjU�\�Br���nr)0`��a�{q�ֳ�R�W]X�N��#R{���T�O�����_�>u�Ѽ�����.�\?���thN�N�U�S������@r:��G���qP1���/�O\x׻�u�uWa嘜��7�������ȹ^�YyԽ����&ᝋ+�������64���]�%2���Ǭ�rN��H�/$�Q�d2ﴸ�)<b����ȑ#��X��Hb��Ū�46<� Jeg�tL�a;��{/���?��^�`yq��r�:k�$�C7l�p��ׯ\�rxx��<m�B�m߾}�K/��˖-#�) l�#({3�:��q/�� �|�S�;<�����o@��Ν��=~�xww7�$tc	l_��RqQ�����B�� No����n�cy���=��m�^z�%�RH]��?��?�v�p� 9��+�����O���/�����g�O���.�}�駁������]��fvFg�& %F��چ_����z�����I��dI��-���`�����j7ٱ�J��$x_5�C���M�!�-}�ᐢU}]��s�e���0��K�Xu�2�;�p])�/ܦ�*�g:��K���Vs�f<&/)�i$�2	z�ڰ��fs m�e�.�L�Ȧ�%���hr��s�YvnS�p��`��(�0�I1�K����޾/}�K ����۷����	p�261)�sc��3��x����]������Z�E��\���d}B�l���J��]�����-�,�iN�!�A�|����������������H8�RZ�nI0K�%
��:�[[۳���h����������믯Z��?35�%IR���bNbQ�E�1ls��?�Nyu�X�/T~rl#��
Y�|+�#������.�;.	=�a	�s0�.��7�oHs=g��)$]�����7�Cp��M�C������L��|)��cQO����l�
�44�햀�(w����ٔa����J11IL8;��qD��Jb�:���/��)����z=��Q�Gj��Q� ����U��?�ނ����r�L�%���׸��W�N��SȬ��Z���_ر}��ӽ����Z8f0U��^�8/J{�p���¼v6�W^r6"/����0��{J'�ŭaz���xF?J�]0`�l����� �	2ĩ���sgfg\J�!CI�R��P8A��������E�	D�����J�Cɠ�Rsɡ��$�9�"���w��r�-��}��Q�a�����|��
�K!#�3w�qǃ>���_��ɟ?	a�5 �ࡐi�ϡz�p1� +�ɤ�I�����#���ew�y�;�)���z���~���R�I����Х�]�2 �v�ԩ���G��������k�Apks��֛n}m�k'O�a�7�r=P�?��߯߰vᒾ��G[ۮ��k~�����W����X��F�'v�������������aaz��_	I"��c�%3�}�k-q��bR0љL*��ݳr�r�ƑÇ׭�R����̙3��������$-%<q�ą�aq#�Ģ�ʢS)�`���z�t=�\+�TKi~��LH}����#K���6�RN�1�%%4�J�*i��<�*ᠯ�^k��dU��Uzs��n/ֈ�h�����0ܥ��U]\w�婩׾.mka�a��];+�?��Uq~C�B�U]�h�mT�_�6C<x��+7~�O�����3�<�oZ�`���6��>�*�ֱN��[Q\A��<4UŻ�*��?��R] �m.p����Ѯ$U��Tڿ�	B���ċ/�����Y����D��Y���7���.�548%��,c��?��Ow�ܹy��e��.]�N��M�	F):��+i8}���'N���u�,��
(g ǰk�^�ݲ�Cj �@bf팫-Ȇ��͚���L-��]&���D��ǔ�Y4�����
�% r<�F�$�D.���Â�N�'RO���	����a46��X��cq^��B�T~J��I,ָ^R=�I�d�㡪�:1{H�2#Iy�둽��j�Z���e/%t���m�½x8��5��N!���Y��c8�������E��殽�*�/N�j�D5���4��ZsUk���cE�(_ޡ7+�M��YbZ a�D�ߛ�]�%$EPX�"Z\e'���dâ),y��v�ݐ���w��1E���e�d�I�c
�"�dt�Q�
ނ@nزe�0BKK��*�N%���sh�
M{�ڵ�>�쫯l�<yb���C�w�e@:pY�P��
��Y�j�h�@Z�	B	��]�z xd���W\qE�!�k׮��;w���<������x0W6l�����o���	$$x�=q�y��A<�2�i�[�n]�zQ]�����駟�я~�bŊ%˖��ٟ� �{|߻~�7�����.�͜���+���o�f�;444==�q�Ƴ�O�?��3'��'�^vZ��y/c�WO)y���SSSTŋK�0��b�N�2xЙT� ���-��w�@,G�9��(�F'Tu\�L���厪SS�}hਮ�]��~� �؞i3O��!��ٺ�qƥ�5�C�
�t^�*r�rЬU�j �.jk�8�z�r�PtO H8�-�A�\C>�_Q�8d	���T�tͰkڔ����S�&�)c�6l����+P�"�gb%-d0'�Y7�a��(^�7i���[�-b��e�`��ųT�b�ˀ�D�T跹����2��8d<��w���>��7?���G�3�4�K�2n��"��2<3�S�=<��7��4'e�A����{X����^�Т_� @	+����Ŭ�l�V�����䑲G`0H"
=�q�zsN`���G��Z�~��?�� �}����]���#�[:�`A/YR��G��u�ݸwzj���]
,_��s������n߱dɒ��wƣ�L6�'�����$?��5+�=|p`a��S�b�����ҷ�P��Zh�.�i@��Q
�" �eK�������0���Y���L6|0���{����t-B�jӷq�,�r�2S�G��[y�(E(�Ϩ@��8aJ>������n�C)�=E�����=kNX�+���NϠ���Y���JF�d��(M�Pr򥼕�xG:��v>�Ƨ��@Bf�l�ł	)����N&f!�:ۄ8iq
F$��bCav搚��"�g��3P`����)�������i�\	�7��U��4]����Y(h��"k����� o�S�E�J�h�Aζ��&%�����pZ�1)���G/!.m�#�R@�aQ�2�)K'ύ���_���u�"mxz�b>����������f=��39ש��&mZ����+r�i	���ڦ,��Y"�1��(���e�/1�#0hs��l����ߢ`� i�EBu,LMɢ�;#��\�2�l�xo����v����w�	����'�	��D#��Б��mh��ϔ2�������R9�k7^V�fSىYJ�U��	�H˴�P��饐�����l�E�/<�o�3v��&G�e<Υ�n$�L p�V����?=x�D1_:{�}[�j5��h:rC:�a
���~�����E�'�f�E@'�dә���������Q�#�f��鉩L2}z��������εkV r�4�K����XWWǱG�����{��?~����~6:5v���,[�\�Ӟ={ ��+,+V����2�ГO<]�; ���WP���pv(-�:�>�T�p�!gٚu�{�C>p���/m�d��.�ڟ|�)�����n�--����j�YWlؔ��d/��>�ho߹s��ŋ1�@���/>�D��=;���R�I��J!���٨	rUJD'��!BP� Z�n��\'L�������0��0�2�p�X�����ߛ������6�	�{��B��FIs����۰�Fr���cK�6��C�[,���d�u鮆p����'�F�_�-�y�����:8���iV檽��2�BX�;z9��:�\ʳj�G�?�	+&�ڤ�h��̪���H�*'���j��q=i(9xD��_��z����C�s�>����5o�I���e���xe�S6����?�c�Ilplǯ��0�J�ɽ��%��m�WK�b����a�;�v��x���}�U�~���֭Xo������`���9"�� ����s�\s�ş��)J�v�-��r+�K��PL��TS(����,��ٷO���nD �ٮ�"'0��T�H^VIqB7�)D�v|�K0n�R��?���0ݲ� �L��s�M�pFٞA�X���c�q(�s�;ك0��MW����,>~a;y��7v|�N��嫂De�ί�m�^?�c�_��u�T�jȵRW��
uR#o,9����#ʩU`�$�vf�\����ozY>P�$��<��������+�<�����l�����n�F��=��V�'�3wk��l����7��`sb:<�Z�H����GJ�9�C(��%6�)3p���I,�i���8��萿����+T�	t����ӧ)�ޤ(1 �ii%�.0n]�z�7����'�|�W^Y�t�T7���x�>��?~��-7݌����y晅���ɓ'���W_�P���l�/݅ ���m�r
�wl|���o?q��ٳg�-�B�A���w>���t�M���W_�,����Kw�y'&�СCgΜ^�X�Js_���l�D�_�u�]�9��
?��O��b�)��裏~�w���� ���'� M~�S�
F������4����z�>��Q�I{���͛7�.	Ք�P?�U��ɱq�BgWQ���T�uЭ��/6|;���6d���V�i"��cG��s/�&���eW��I駲��M�S�Dg�ą[�KScVj�sm�z����Ǖg���j����I��k�1/`H�ams:����+*l���ir�8���@V(~�N^$��[&8	J�l�;�M�d,�/�E�vq^�~��wߓ�d���<v|�5z��̭ق�M�pIZ`����BY��ʨ�*�V�B^�+��e����e����f;�5���_bTjj�;�9�MuC
-@t;v�P�5���p�5��{������SO�R�����dbx���G���*+���Fca����]�����?v�����w��N���I�@�]�l$4Q0v�X�h;uf}���B�C��;���8��x!x�R�XƷ���m�W�$��z8�|^2�I��2�ŊT�H^K��b�����m[�lkjk�#F1϶����4p�Y������_T�_:���G=�s�0�|_��ї�H�4?U�����('{�\�y�PL=�d٩~O�Q+�T�e'�z>g�Hq|������ܛ��qU���:=�>���Y��X�-y��l6lc0[�@^����x�$���@L����@�`c/8�-Y���Z�]��H3���3�wU�眪��=#ـ�ԧo�SS]u�s���]�Z9�"k;�LV<�j^#���Պݔ�+d鵴t:�����J0�C>��U��2�?�����4�3u�_�)��_0����U�(K��+�')Y�wWv��Ry�P�m�VVV��J(����9�f0
;��O�nd�E�4ƿt�|ͽ�4��ýTu�J	+���_c��f����ɪ�
��r�cm�����Q���۷K�"��1��U�K��E�?�����GO�8!�쁟�zz������ֶ3�u��]�����@�A�b��֭{��gΝ飯�z��gA㦛n*)�%�)��]�����7���EI��4��ہ���?~�É>�a0�
��A.X��ȑ#�@�>��/��* �u�^?a��o�_��~����N�ko�0�]�d����r�\{8L*͂e ��HJOO�_u�U�Ugg�o�)��r$@Y1~�,�v+�q덋�Pw�k���l��#���иe�!�^�,9��{;���ْ��������u��������Y�4(�*^}����o����o�x���[DsFԇ|�6���&
}X\+�˓ ��I�VJ�͆p�Ce��\V�F� 09d��b� \(4 ���� p/�D�����Y��r�������/��η'iZ�-��R9�6E��@M��U� �y1"�+4���`r�JO����g[^�x�]w�{ｸॗ^�J3�47�|׮]��5rp�s����,�g>�p����;v��r蝵������(���J�2�����_��m[!]?]9���UhO�j߲���qI�:k��Q��x�j�s���q,�Դ����o$ٖp�I�� ����$��3�������|��p�r :lQ8�\���h�\��^,7����挪@ađ�_��-��Z^w�Wc�X�"M�
�Ÿ(u��~�;>�F�����(����6W�q�qz5Ty.��h�����6�OuM�Ng�.����n��Qf�0�Ol�����p|JN�5U$HcWD"'��X͝�t�%q2����{�	��
�#�5�4I�&	^lE�\�@�(3��x@��W��|u��%J�,�)	Ĥ඾�@��/��1{��_~y۶m0���ǧM�&`⁁��z�{����<�� V0�k���̓�<����f�� LMMc��H`�K/�t�m��\��i���k֬�������A�bH�^����>w��w?��PYW�^�	�1@޴iy�-����kx�z��Q|���+�<}�4�+�0k)�?c��\Q���O��o��_����3���/a���w@���3�dpGi!l���0a����ӟ����q���*���#�J��	P��HR�AT��}��Y��,j�wh��a
��)>.�2��z����P�'}V^�V�]���w��(��Hn;�oA=4���r
A�y���8�������b�zQj1�َdZ��t�C�u��B�6;+����|��Is�1�Vr`bۻ�Ĭ۳��t�4�G��@ �E�-�2mꯟzz������N�j��"��q߮.�g,_�"_�Og2�������|��o=`�	��ʙ�WGϛ1��XdetGK%�X�N�-����DцA�J�-��j���)hW�@l��ח�"��g;�/�uם_�����,���L�57���FK�`ZL\�:q��S�%��R��������!)�,Y2a��T6�?4�B�Q�eÀĳεw����f �7��@ҩ$tk�Nj���!�5B�S����!�Ίu�E=�ӓ�[�j#���Y[p���Y�#���9�g��)�>��yE"%�t�4(\쵍[~���]������Yn&�JeQNn�0%?��qKb8��jL�A�D }F�xK����` 
��%U<��B�����tϭ�{��t��.�U��1Zn�C�4ߛ*�q�w�_���h~!��,�9�����j�.�'�*�kA�2��5�\ƭZ�fH�
��dKCO�-=�C�L+G������#���LB� ��L���Mo��Np�.6��R���g��M��h��Q�Z����=���Z J��,�~�5\SA6kK�&�V*S]SSU]12��#	��V�5���Cǩ1yζ� ߃fH��0�:
�^g�%�B��s�J�.�W�Qq������M7���o NZ��_���**�`Ǝ���<O�4I�g�:�ZYY��6l�y`���練�;v�Rz,R���`C}&��X�d2��� �y�|�C��n��A��+p���	��<y2ntm���nڹs'��C� �4/�r�#w?���=��c�P��p� PڢE�p�7��!�׮]��/Hf���[qOȊ믿��{>	�����9y������o<��T�`�n�ׇ����(3����ĉ��h��Y+�M�
%p�P��&�ކa��g"d�������9z�61\-	a$��.5G�ڥ�"�4w*�F���%���n���G�z`�,Bc��3uga���7�B��	�E��;s�:V5m���
����Q�X�`W+�<Ē@ۃ8;�W�<N��ݞ��X7�V�pEM�!Z ��m	�ʞ={$�I���\��ܚ� C��n'�/�r������G"wuL\"�Y���B�f;�@l��e��X!�_M6%*�֭[����?�yp�ƍO�h����apˁΞ=;~��L*��S2>TYSc���Ǐ���;!k   h��9l����ɓ� �~��3��6Q��8ҴTF��O�p|�c�v���p�s�iT*�?s�
��h��fA��*�a?�Լ{�z
��� ������u��@'��U�;4Ȋ��)��I�QB[3�(�fK!47��4��|�J�E�p
���ld�o��K�Tj��b�֛�A�`�/����D�A{D
���dR�s	��tKgr�l�rP��]��<
ԔX9X[c��=��K؜Sy�b��X
�^�Z��9w�L�+�N򺺽>��~���Q����wPh_z r��HZYs�U*���<���=b�����g��'VW�BG5��LE%���{���K��HƇ�gXk$F��Y�p�Ӗ��S�q�� FQ"Aj�y�}<c�]w݄	Tmu�QB��֭۵k�@٣�4�(�@�N�4i���Jj�-����<&�"���q;� ���˗/\�p�����"�<�������M�2�,�\�{����L�\[�l��Ǝ�����566₣G�B�.X�@�Ѡpy���F��o���5k�H�!��}���㮻��?��?b �ׯ�9{�=��SYUN�7�I��ꫡ�o޼����0F�ׁAb<�9۔��9�0H�~h����5(g�Vј��y2��֌w���(��ճK�u��v$U���F�^�G�q���~�S`����7�L"�t���HH�h~����QQ]�.�ݢ?���O�[����r�g�b߂�ģ��"�J�������nJ�d�)��p+U&��0)���Kc08Vf0H��P�d:8�"VR��/uuu��:�#�tp�+�[��B/j�c�un�M�Bf9�6��vI�s���p<߶P�{ڑ-�m�d�tl���/V���
�S]MԠ��V�s\b��mF�:�WQ�$L���,5��s��3_��W��v�w����W_���Ne�y��s �8r���+�T�ȵ��r4�`���O�<eڑÇ�|�I(�X�l��;G ��4���2�O�D�H(�Q?JG�8����BوhIl�;H�2;Ec%�l�ܙ�4�6��b�@{'�&�ʮ#�1*��[��YhJtڊ2�D
r2��'�<r�$��L�r�PԲ�k� vu��L�M7��x�� �2Alp�˚�F(�l��!�y���P2�vt��+{fA����x3�E�58G'$NF�&�3�h���
����U���U�t[C!3ؙH�C�� 8ˤ9�D�JME��[J�s]�s6gbQ���U,4X�s(�tu� {߰�ee F:�=q�ԋ/����7.�x)��ْ�$0�w�.���j�3DZ���#��%H��R��V���q7.�jY�5�5�U�a��p�Bw2����Lg�k��6�r
�5vE7� 5`AWw7�,*�d�D�&d7�^H<hs}� �Y����B������v��J��PUz����q��	(���򗿄 �mqF��uuuA�Us�ܩ�o�38�����C�����PV�1M���L�Д��W��F����z�NS�h�΃�p
��oɒ%@Z�s�t�Ȇ(�НMSaX�@��P�������ǎ_����@] L�mj0����n�e�muu5;wno~swυt����>����~D������}��������5Z%�e��O�:u���߿`��O�4jNggG}}�<����K_+��� ,�=π.�SMϹ��"�
�I[���N�8�Ɖ�t*�5�R����J�nj�S Q/���?�:��TU�Ѽ�(B;�oV�R2S���
~�Q7	��L���u_ʷv��mJ�"D��%��Z�I�ކ/��5*��T��|�+��Z����*����7���o׿��V�_~��+6m���%�=�W�ر����ߓ-�L�s>�.�dSܘ۩�gt������qBA~�!����>���1&�|������w�!��P�]�E�JÙӧOC�~򓟼f�|~�ɧ�F#�  ���F��lh�?O�H�_�җ�����;���ph�s�� ����3H��A���5Id1��1g��8��y˒�
$�$��U^�m�������Q	��9�ɢ�FŲ�^�l~�(��WhVT�L��y��g�^ ��˩J{� /lAT�,I����z�`K�ȍ��L�8���-��P�lW�>�b8��'z6�^�h�dG~��;��)~_EX\�ka[nǔ�FK�C�<UyUu>��q ,ݐs���Л�"���.W�H���l�MBlG�K��v����j*+��I�%���jl^�~y�����&���h���(l�^��JA��̮Pt�u5.�SI��J� v W��u���� r�l�WH�蜴I�R}�A�/%,I�nz]^,�][!i�4*���P_���^+W��#{쉻�xk�ƍ ����8���fΜ	��-Z��BpQٶ�r����; �7��x�b@��f���5kֲ����	]I�G�;C`B�R�m�@T�.NR'�v�g�2���#G�Ǎ�_��r���o��؞ �%tϞ=X�'O�1������/|j�>����ޯ��x���׉��YxG���Ũ:::�SV�4���Uȵ�\CX\)�@oIT#o?ﳅ���Ñ��a��Lk#w1��[���m�l2(�h])\��,��,<���S�ೢ������×���bTw���Y!xRw4F5�_|AG

�� �mu�n�.T[H�*J�a�?×��S��K��ۆ�F`��"�\O�9������'JE)�d"3H��3�#0�/�l�F"/�%,��H��9b�^�je����^}e0><uL3赮�l��"�.��D�-��&������Y�ˤ���D��t�����r�P�ٻ�O���P2ۢ3�����/t��^	Sy�e`�	�4;�{�|sc]������ܹ_,�����QꀞJ�1�����ȟŶ,�e�P0d�e	�MM��/|��q��������荵51�T��T��Jh����e�
[+���+�/X�����/��
>TWQ�CAT,&�5���Xqyo_���?��8�����	hVt_�K��BնW�2,VSv2�䨿��Z�����;n���%$�2�<P'y����~\t��-�F�B�n��d]Ӱ�H�V鸮2WK��`ٴ�A"wu�l۶����t�HI)����UTj�q��M�D�ި���d�s����0��iJz�d�������$M��$Ճ���`H9��o������\��}. &4z��8���@�i^
�L���R�9@�PQ��W�_Z�9RkѱsVV����e 9*����>j'��deh��me���������E�{V6�Q3&U�5�0��`��鏖ƛ� 6�ŭL�B��M��ݲj�rpe�K:�T���T�!m�^����ڢk�ϼ#��Z�ޖ�����\{|�_�kM���p�J�R�����4Z]Mm}m]yIIeE��p�0����o�njl�`��0^�)�{�-(e5U�uu�e�j����W��KE����t"@�����OZ&��������n^Y^AMR��S�z�`k��p0�Ii{v�>9��T�7?�����W��x4<���6  �+�� ԅmbΜ9�g�� �n�hJ�/��s�e�iƔ�c#%Ѫ��x�������G�?�jժ��g��8�>u�!�9(̲e1A'Ԩr;�@v�\:.����m��]���^y�\�|�J�Z �1c�0�iӦ��}���wDK��ώ]%��?���?vݺ��������7��  �o��o�h
d�ۋ)vqbl˖-;u��3�x/\\&$�=�0G�ӳ��2pD7S�+�A0"�7vJ�c�-��f�";�0�t6
���/B�P�@�5�7��8o�HF��r�O�4�1�Hu܍:�b���W{h>w���( `���G�!����,���1uf����M�j�g�	t�_�;���_$�Dp&x��� \'��)�^� >_:�ř��A`Sufr��w����O~u�H���L�C�7s~uZ�Ũ�W<.�Qc��7�,9� �C��(l�Z�44���1Q�,�Z-IB�`��^R-b�<V���B
L�<uÆ�h7���XF�.�ս��wI^S*M�j����>�m���_��7��ͳg�B�ںu+dD&C� ԅ'�b2�a�� �ӧ�z�W^�����kqs�����h[ZZ�++�����z���_�9��^���0]��.��*c&{�}�y�w��o�P��-B�R��s�%�c8}��; 1e�)++Q��SKf�W�0��LT�Vzy�%Y�9������:��˖K��B�g�����d��;��Z��-�81�y	&
���ߺ[�в���C���U����s�a�3�)��� 0�Gc�\[�M�.�T)ڭ-��>zt#ߨ/QsC�� ��"Kg��E}]�D�ɒB�HH��J����|��8�d���k�L:h���2�hQ �e�´aҶI0}	e�(��t�:��}� s��8�2��$��^��Իp}������E�I�m�M��K��QD(����tM�/�����dy��W�_�~��e��{�=��/�`l �� q����V|���x�w���O�8�&^�8��k��;wn��y��R����͛1c��2ʦ\}ŕ��O?��|�C���=EgK��O}ABa!f�A^�!Tڞ���4i�$YcIK�ˤ�fz�UW]s�5��οb�^�u�O9v���Gp�ÇCnO�:�g?����;�Hes�7s���t�1����E@��� ��˗�۷���s�>}zii�jjj����Y�bj�\�K�磺�S¯I�g٪d���'%���ŕ����u���y%��y۫���������7��E�v�?�Q���[w7�L:[�?h�����˼�q�m]�cꔽ���ۦɭ�%�M�E�dST�B*t8�BH�w��큁�ʚ��-^�z��_�c��hi��r���:$�)E}ٚE�D&��I�.��e6W^��\���t��2��K�u�0��C�9\�֭��K ����oI��XI�,�.(5eQ ��N��'N�gn<����b"�Us�̞5sfyYl��o��Fg�9ȝ�r7�Ls1�!�z�0�w8_OÎ�e�(sP�F#��p���`EE͝w���O���w���~��'�X�z��9s8p!8n\�l���$ںk��~�/>�����Y�<��X�*$��I����VVU��� .e=,C�3�N�#^�%9N(J 7gQZ�P<np��"W��i~+�y�;�>�_��s����u�i���m���[F�ĪF!4����[�mܼe(שo���&9�&++���.4�(�m�Ӧ�)����b��}�L�R�J�"�V���*@(���I|8+)�e�E(h���N���!Τ��i�0�,.ف���!BxC�$(6��B��*j
�8@;��`QD�Bۺ^l�T�FA	X�!>�Wp�XA�NU2�W�T��ΒRnJ7
����H��/���!V�b�L��\_�f���mIum]M���
(Tx���T(Z��"�A�)��g����)X�K��O���K{����׎D��b��Io�1��H�hjlX0�Ⴧ ������'c�U�H4�L�1#TR�0�k��4$�H�9��lg��	��e���p$J�x��` $fQ�l��Y�l �MsY]�����vC�[�n��@cӦM[�b��͛q��ڀ{������U3�or��2i����~��'��� 4}� OS�O[{ͺÇ0Yv�{���ؿw�W���u9z4���\�nh�gΜ@�y��:������m�pR
�RKۉa�s��Y�d	�d:>À���o�����~����A��uu��;w6$}}-`��`�D�|���O����O�:��������?L��n�u���ԩ> 9Q$JJ�}}�P��D<rF��Z�,��2�l�M��z���i��8�'m��3}W���O7l�jύ������P�\.��@�wU�5���3N�#2��n���^*��/��2;������Q�����W���qx�h(~�t��}+�&W_��Jk�p��C��lLbj��	��캗����%�r$�s^N��YH`���k��u�]���/�՝�����lN\%�LD�=.���P��L���|e���~!��Z�8�å�~SV��j���u5�V������(P�p}G$B�$����1S�L)��¤��?@mmtR(��m�2���@d���$r��6xZcI$�iӦ�+����G{��W��;w�K�}z!�,S�S����];vJ�8�����ζ��N'�UT:t�{�����Օ[e�\�G`y�Hx�:�x�X2��N	v>f��#7y�GAr����t�&�Z��Jq6�={������K��%�3^Z^NUZ�/a:�c�-v8�"V��W)�U�J��4)(#�8ō%�R�S
�=�b|��(��*'qB 	��m�$Mya�3eI6d5e�"qP��Jb�U5|KWKT��j������n�K<HF�x554�����g���Ո\xu�(7avL<��X>y�d	��yy�X[�C�8�J:N��ޟ�ax�*l/�[�5E�R�À��^�@=L��������֏��*�\�%79|��X��&*"�|F�"ay��W�N��{}����@E��x#x�@?��A*��z��ٳׯ��s�=���9c� ��0� ������>��ŋ/Z���W_�A�k^�t�s�]wΘ=������{��---�Ƹ�����ѣlǥ�6˗/ǐ �$�Y�J��u�	S {ؖ3�
�I<w	�sxH� K@����_��ז.]J�)�AI��6�8ۃ��n��6?|�K_���_��X�o}�[X��3gb�R��'���{��]v�e8�mvS��l��?�/�c�sѧm�ت�P�ɏ���Lik�Y�%����8�����k��y�uI+���W������!���������y�ת��H��.��������p��ܩ
Z����u�3T�j��*Df#�`��$BY�$%�!=��;��Wd�e��|�g�v]���������'�z�ҜҊ�T���X�v��)-5�:�8͔�P���5�5��L��;���(0�i@��MJB�.A�?6��y5�ln%�p5�����?R� ͢�ڥ!峧M�3sFMM��ͱ��������P[ә$Xly����8f̂�7e�4��ֶ3౪�*��D|rA�먁���P)��l�m��������[��N��Y�g���H8Ke���g=']z�%����@Y���??e�d<����o ��F?�����j����q.٥�|��j�XDθ��$±�8�G1I
�jof	��o}p�_A �_o����%z^��E�=ؖ�<�?r�x8?n"����t.�L%�k������F�P�b�VR�-Ͷk�)�N̤�+�����1(�A���l��Ĺ)�[�Mci�^�R�U�%g2?�ZK��UI$Jwwo�`������0f��\$����k�X����d�H&>��E���`�w6R�jV-�e1bURح\"��/�n�W�9�Q����a�S�U���Q� �O�$a聓'ZvV��Jʠ��m�����)-��p6O?~��S�Ȥ
):���/�G#�K��&�SP5��`8ZUQ����]�d����;��UUW%2�P"a�M���uȐ���S�Ng�����<�9�n2 '��Ҙd��C�|��\tB����d�%�K(`���c�u��Mc.\�<s��/���]�v=��z`2pTyi�A��9�fO7�<:�p�?z��lǮ�}�+�̇��e�׿� 8:0�'h������۷��j�7��mڿo��4%�(3�Ei�ُ$D����D"G�v$.�r�@Q�����%���k����	���<����5����O�0�c��_~�-�y��]���ﾗ^z	�~��������|��ɓmm�)������}���U������I��M��_/��#�V0�u��c�H)p4-� �<�� ;�	�wj�RJܪV��Ȗl�����睡
����s�EV���t�: Za���0��O���|ڠ�.�^z��]SO��#ݳ���ǋ�qM�����B��C$��J��Z�� ��<�z��i0�{����O<q��A*���n:���n���8�͍-�#�$5Xc�=}�t�1���;=�+#���&�،� ���p�j�(�<<C��t
�Ή' �$�\�Z:��YYȈT:���0��m�h��R;`��ٚ��DЩ�cBtY�?��q`�Gyd͚+n����^{Jd]}�766��b��InF��M_x��p���ٳ�@ ����e˖A�UV��|}Eྶu��D���Zd�P� ;�,��ş�s*�cl����L�P�)���ş�y���Y�dõ�����}F�x�Ѓ�2�7�cS��@ZI�3��_|����0��RC�\
�|H�2�vX��h>l����L��L� 9G�*rt�T*�,9�2� ��A�d�����w�)��2C��-�"�%�N�ebuP+ip�M%[��3��ً8D�1b\��lw�\3�?�����KkF��F+�{�n싕�˩�����Ԋ�z�����T�E������EK�0~�bC%���m���^�tٚ5k��?�l,K:9�W_VYA޷�Ѿ�ٺ�K[Q�)��ҋS�qa cE�ԅo͜9|��B~x���W�^�v�O>I�29�Z��J�SӦM����tȻ�뗿�%^b	��� �h��.1����:�������(-��~�Q���WL��_��q���d2-�8�)c���,,=W�b.�ƋEK|������q��³ (q�-[���Vc<���#G �1*Я�fb.���������FjQp������}����l�����ӧO}���Ŗ!U�|�]L���]V�5r;R����ό�%]|~�Ų�^��/�U��
��N���|�<�m./�I�M��uF�n\�A/���k�<�G^pH�I��.~���ע[��ʼ���%3|��/�\�g�cP�bҒ�/�:�X���|`GZ�|���sO��B��8��kQ�Kj�B����j�f��e�bc]}}5e�F�sg�9ph?;SS#�a�d�=�̀Ial��s��׵����k`�x�،�K��u��r�Ç�::z{z��{�*���xH� �8�J[�"�ۻ;�MO�<u���˗]��ot����QA͕�Z�H�0���������HMM��{?��[v�C���l�} n��榦�H$d$+�c)ב�V	�jժ/m J�7o�ĉ�}iY��R\94�q����F�djr�a.�S\d�[s�m���� �EfrYó�\�C�0�?������\#LA�I�� ז��Fנ(c�����M��{{�5�f����T_?�2@
}_H'�Ȥ�6C�H�������N���ۉ����1�G���AX��Z^/������F�z�p!5U���6�� >�mClW�Ż��2�����YR�M:�	(̗��˚f��FA��h)K�mKt����h�s�a�t�`w9�ȳ](������JV�=/a���Xn��|�1��&���c�ȫq�aĲ+��"����(�]���gBP�B66N6g���N�HJK��w�̙�h	�@R�\�+k�egЭ�]�A(�9�:����@8�b|��8����\7�2��,���"PnCpÉT=6�X -,E����}{�k��j�ƍ�����믿d���O8p�_��رc7o���'V���
� ���m۶�A�G�|�Rno�i��;w���с�@�?A��N8�p���W�կ<H�{�R��!�L�ׯ���^\� �pg)0)&S(�Rϟ?_������p.d�瞛4e*��#G���J �������������w�#��ܳg&8vܘ��ظq��I�W��m�� Q���������Y6|2<+�q��@xĭ�)���|Qe��gؑ�:�c�K�-��b#pcl���'��b�x�#7��yw8�҇ajE�И��ͨxy��;��Iq��r˃ ����6[\�β��8(�,��G}TH?��9	����흝��ܙ�9�]���5����b���ݻ���L��*?v�Xk���Y��i*�3�}I��v5��T|�.&V�ʛ����sd�۱cǌ3�/\�4����{r�&�����˩��I�&a�X�r��' S2i��Y�i�s�;�0B��B!["�x�!e(� `B}Ĳ��G?�C�B"@�;w6�����҅J�P����Z\�mӖ��~��˗����L69
� ������޲��MV�!���i��r��B̞���#�?�\ldh�
�	��1-�0O^�A�̕;��� �,� ���u���[<VE�h#�S�n�k6��>����4H��3%%��La��ɫ؀"�����j�TO�'8f�|�l%痞�������[�3l�991K�ɪ� av������N����4ݛ2i;N�Y��{(�g!|��?>s���;�X�uN)�?�<x{�ܹsslS��\�^Ѯ����]�B�(����\s��Q����64`Y 7lo%�i�`�P�e�k�XL�؃���A>dq@B���d48C�Z�S�|�|Y��9b�[��H���Ѽ�u	UUU�]8 ��C9a@?��ͻ��^y��3�  ��IDAT��o�>��� :!5�����gnE�� ljh�:~<	�����X�8�=�{>��3_����X��u�&<��vȦ��f������9K-�`(��׭[���/ax+V��C��8�� ��ā8qg,62<���l��mK6u��+���l���A����/0������y饍��eX�?��?���,��C���~�H���]U��ӊ����vI7E>�YC�bݜ��4����.��ċ�m����\^7�t��8u�h��w���#̀ 'e� q��u���c��N8�o��
�3��z��(*YD�,��w��Qa`*�^�/ϔ~]�H��$ӎ�������nB���a��H�h�)N�.~X�Km�x&Ew�H@� !T�ڡ&H��p�����>�矆���7b�����[iA�v#<H�z�e"%���R0p�ԩӦM�\^ٵk+&�V[���6}�������|i@[�tIUM����A���W%�9�(�0�@i4R0��w��;���4��`� ���}aɒ%S�L����銔�������3���01v���.v����v<%ÒB�Z�x�ҥ�4;Q��0Ks�N{[0@�2!�o�`��Ds�u�w(.5f<�i��ܲuǟ}�������O=�<�a����g���@BJ^��ޛnni=��O���z�/(�����D۽c��5W%��z(942�\.�w��2WҭKw���H+��1�וˤ�L��U���T|�Q#���ei�v�0G�qiU0��t�xMgty��hO�7M8�0m�OnȨ�g�.I6���6�l߾}���өL �n*�&\|(Δ�����h���\�+0�kr�_�	E©���Y&Q���I]VA�"�t@�\�=hG�a�k1l�`_|�K���-spx/�ԉD���f�KB��!)�K59{ �U�n��b��͡�%�0HM��-.�������e	q-��<Lֶ8��� }J3,�4��0mn�`mǑ�4�bM6����1١\���s�nq�td{��s�s(�"��`!f�N>�F����biM�u���Hl�9+�����uæ�/��K�@����H�q���R=��W�b�.�X�r�
[�i^�Z�.�v�CIr�����"�ł(u�8���bؙ!o�"
��9N%�u9#��_�����>���qJ�L۹�S~��" �Pi���*ޞ�&2����,��l&�+dõ3i0��s��|2����`(���<��B{��8o��={�l~}�'>�sg����P2N���{����ʞ���'w��5X��[�w+.�H7v��W7��<f���e�-�����0Ͳht���{v�H�O�<���!3,�b��2���}���̩��W��@�fp����`���%��p\0(h�%a����u,��[�c����Uf$�~�s���c�Ro7
��t2����\&��<sƬ�s�?�s���sf͚3�׿~2޼E��]ؙ3g��_t��~�߾��˟���K�����oƌ�C�C��U'����}�{�i�m�4����I����!�i2�Q+�B��4`]�z�0 �8�m�'�'�~��M�%Y\,��&1"���s�Q���X6��(����:v%3(F�Tq��H;������Pм��Fa����W���bm�����S��,%q��c]zPUD
vׂv��TZ� S{7���cT�Zq�VhQt-eo;�ۇ|���X@��3	$�.E_�ʦ��t`��9��Amz����k֬�4i�֭[��ڰ��G���5{��tQ�a@A�Vв3P��c�NC��4\p��)��ҥK��M�0	;�P<��xK�C.�a�t<��f ���uh������%*�X�vmMMM�]Ee���H(O�Mz�N6���J�%�@�0tG��w޹w��M�6��0�m;w�%/G��iIg�T
1�``�>��ĉ�?��Ϟi;�aÆ��@�WVW��T��%�a�u��[�lٴi���;\H��ѣ����u��pcc�]���QUZV.�V�1��۱�ME7M�B�+2p��f�w�QD�E�y?�\K��t��.Ն��l�/�`��H0(�hm7�����d�p,��k����G.�	_VV��z{{�>��<��I� %�Kb�mR��0y7��#���Խ������I%�:�+ӝ�����bg��h�-W�yD%�������*)�WB�	)%%��	��,_�]�����ROJ��/n�T]>��q���}TY�~q��`�j�d�R	��:���ѿ31�߅��~ռF�BZ�P�RMk�Yr9%5�]�!�	���6���M�:B o2
d�#�K�~�i�W����:����Q��Ӕ��!9�KC��V,hiig�}��'O���F,H�";��nV��W�޼y3��u�]��O�<y�)�?��O�ӕ+WBC����0T�s�Α��Tl��\��0-�	[@O{{͘1��ۿ���N&�q�36K�=�7��0Tq��ĉqg��N���G5ɪ�un�+��3�Y����
V���7�x#�����3g�FH�p����;����������~e�>��O}
(��W_�24Y����bR�Q+��GR�."`�Ak�5
6����YE,�tu���NE���d���_�:�"��E�>�KR{]� 掍�2�vKm4�*ůS���A�B�i>@�`��o��ȑ#�ׯ����`�l��͝H(,�A:�I���G��H��`�=�&	;Yee�0]4�拓x���S JƎ�Ra��~�7: d�HQ�M��ô\�&t�p@/��0�D&1���b�iiY�Ϟ1���ӭ���K�\�!V�	�3<D .46R8�
���s�Nȋ���|��l7��(3	B�����	J]L�$7Ӊc'N�����k׮��{ꩧ�/_~�5RR�,�"�V�B7�t����^��9�f�v�mX_w�T��D^L&��e�W
JCJ�����TᲴ��N�V�S���
���F���(%*�ĉ�}���N�4��49)�n.`��'ܜs�J�^fõ����C1=v䨠���F�2����1�F@��jƣ%���㜴���q��;iU��RJFS���R]�|�*���-J�W����U��q��adj}���
w����R�CG�x7��V�L|a�&u��}�!�pP!��.z����N�S;�y¤�7f�Zin�y�i�����8i��>�V�Ƚ��U/8��B5A�3'(�D�o��lԔ���%�4� &M�h�l.#t����D:��65< 1&u]����M�R2n#f�:�1�(F�0��ĭ��| �#���z22���ax(���sߕ>�Ғή�S�L��{�՗�f�̙s��A�	 (Bq�TP	|T__/������P���D7���+�H�[�����İ���Z�R��||�dOC����sq7ȇ1cƈ�رc���4����n�w�b� �ŰA��0.�͚0S��e˖AO ���2��m�n��(�]v�g>�'�xb��7D1۱c�) ��]�t�*��b��Z<��a:TE�e������cI�z�QD᎗+����ty������7u�)QA��r���9�"�>�枖�S��'I���2���w�A+�R����[��ޏ̼u�_Pp�0���9�#�B�Kw��ݷ+4
B伡��S� �`���?����S����.��+51��Y�&L����7oxҧ��G��2� ����>-lL�k��+R���q�БX�,s�
K��Y�f]{�G�<�DE�VWS�E6%���ec%@�I�b2���۶q1��b��A����x�&SI)\D�ڜ?�v����^�*�d&kATmܸ��#�m�޽6���O664`x�Z2Cj�S ��A:�c�=��C����]xKƎ{�X�ĉ�$&E%�з` lz-��d0���� 5?�S���?�x���T����
��.B-�d�=�in�a2I�M°���jd�E��@l5�a��i@=��82��Gc%b'����j��eT���dM
V�g�YK�IAf�#�i�	L��`�*�KM\/�Q�uP�Faq�W�[-�_��Xc/��y��<���� ��/+�7��^��g ���X���#���8�W��)���6�Ű@�J40o�l�!��$/��h��{[����6�)��h�t�^���/�ZŜ	���)`��V@�  <��ٳg_}�U�$�!	,���y%�K�K�b����
,�H��U�;d�M�q+��w�G�p� ��L���k�j {���'O��k\����D��d"I��B����W�R����F����{HD"��MЪ��C|5�o8���C~�h� �\Z� ��c�zz1H�*���r�U��-�*�S�|�'O�ǚ@����jc��:��S���۷�`{�Ɛ�2!���,�L�82{��x�}7߂��یǽ��X�Ʀ�q�@�ڜ�ʮ*��O��Z�r�߹YD�~X,�e�
FB�"����p`�}k^��x���<��Ǣ�p��]<�k�~|�����B�ܵ|�QI��4�Ϳ��A��|���A1t��%�pA��P@Φ({�@Ow�i*�+n|�MM�cy�Ç�ln��>�J��PX�[�P�0tS7Av�@0	�o��څ�NPyCC�cb�P�D7��IIj����֬Y=e��͛7C�a�%!�����2�k����44�����]�gKc�[�s=�x�����V.#��M� �ZLn:-�r���a`p������8^���?��_z�1����2%��P8��܀Pw{z�qg������tvϾ��V�����o���mۯX�j��a]ǀm�5�9�N���9e1"��?�1�������1ͳ3�P0�x����a��**2�+�p4�%}*Si)nLeϢѐ�g#9��@m�����q��}�v�{��2�Li��ph��=�穻CD���cPo�`*�5��T2�͈��--����8n1��0�?[0b��'����V9�^��+�M!�yA4��q�tHQ%�@oR8�����Ν��@?v��4����A�.֚�e���v*c����"x��ShZ�U���h���)>��.�-�\]�E,�� q��'C&�nrܥ�ʺ���"w�b'�xTAN����z4�M�Z���y�k����ǎkll$�pp���Fޱ�4p1����#�w�n�n~�C�)�-.o�-��S�Aa�g| ����h���h���m��0w��������|Bn^���(aqC�|ְ+�9�@�ź�OY��[HH-�\����G?���}��ϟ�d#_)�$��ڹl|����3m�z���m�g�d+��4|i�6Ę��]�0��L˙��$g+�,Ter�����h4\V6��j�a*���@P/�N��9�����X�P���cy���L
#"ܽg���X��h���c=���}�{��e�ٙ3f�m;748ܖ;;}ڌ��tuu?��S��צM����~����/0Z
|���[v�R� ���fJ��*R�T��+�_YV|�����]����X��!�%]ɚ�q�v>��2�ȫ{uR�-��ZŴ<��zޒ�B��_I'wT��j�J�a��O�P`���ϴ���o���^�O�w���W��jl�\|������a@;)�샃Ð��=brP�����A���+��8�z��9�K��g��s�׎�,N>s�,6��S��[�ϴ>|X\K``0並1X&C�8	~�y�{��B#ϒZU�J}G��8� ��2 *���hg$�ϝ3gV [����5.�M�E�$��jj���ü�	����	z�3�<��|ٲe����C)���D�c�LK�
F���O]]TLA8��B��j�Ք�'/'�F���G�J;���ҟ��L/���}JK��b.7�~�����F�_	��ˤ��ґm�C��5&���T2)N"I9��˅���5�tk(]������p��]�K%L\��ʉ�:�"KT�F3�Zp�{$a |`�Y�h���@r�U��ְ�Ȍ�Q�O
�(a�wnj�P�Lv\��vX4��A��Z�$@���+ QS���M��Ȗ�E4]�冠q��l!b�qM�a�Ɠ�j#��չ$��@9�+ƚ�[��"$�O�WR��㿭sIۘ�{����",��IYh �����$ ɶ	{J�S9�Z��r�����[ L�?gϞ�����ݨ�uz�b���S5�� WFt�
)�w�5�/��R�e_�j�������^����o��o��0���fC��5��PKr�1M@����I�&�HW�릆<K�G �I7�Ag�"�oM�4o�\G;8Q���/!�˘�t��y9����0`0X{��=�:��w>��~����Z Q�[g�� �y���>c0)��R���L��{�nܧ���̙3��-[�=ڂG@D���s���xB5�5����?�߽^υ�Zp��u?�t�-��6	Xѧ"����8�_w|�ܢ�]���50rnnӫwϦ6r��O�wڡ�[�'�I�XA/���Z8�|%ǳ�j���6���l���DJ'8ƿ	�&�8��/�`$L$Ree�P����p&Ef�!���+��Iw�,��WW%S�S-'�i`�"΃jKJb,���!��i�S��Ul�v�ls�e��7����Bg�'���[���IP�@����3c�j�y���'ε�TU�IR;�$�-�R݈CZ��F��<�7�cH��������n��m;v�����O�<6��z���c5��T0�;y�'���=�I�B�#kj����G��drk��v��<�g��v�څ�a*r�Q��\Oo��>�g�p��?����m�����W_���݇+�*(Xoƴ��_s\�3H�Ǧ,\��%��OA\;vN�S`��p)����gzg���腍��xl+O�@��{��t����emxBٲ5�/?e7�)�Dג�E�����&���	�]����i/Z�D�d�֭i __�f�S�B�DI	e�BI ��ث�UK�"������{Q���f���
�B��ʇhn^U>�����ɂ�A��cCC��
��d;�Ś��
���v<�AW����7@�cS\i���h�"�#�BE��d2����?�u��3gͮ�����Ng�ԍ�m���樼£x<����H�b��b�Q�|�t�R�oe{%�鵓�H�Pj�A:���1 ��ƶ�dUuum}]k�����>f_���R�DD�a��$ ձDm&B�b�bv�`� � ��شi�ꗿ��|�+���WǍ�X6�a,���6�`��9XiI�����K��P�C6;8<�70 U�����$KYi>NVV�gө��2�ó�l�r�s�t��!�S�d�Jrh�<�(o�J�D�R�𱡡�����7�e�����=���|����?��� K�̛��������6?�ײz�j�	�Õ���=�1_p1v�%K��q� v@�ǎy�G��}_���[��IW(L���w;�Y��b�^H%+ɺ��4F"\KsԮ�~E�N�<�
�<�Y9ID9��}��0=a�?	�f.�%|$%��-@��T��g���J���|H�� l��
����F���
�	�O�~6*�+��2E>kg��9�����ȧ��29D;q�V�Zl�"����ʱ�@� c:|�0�v�a_��mmm͍�Ü��ԬI�n����g���t��!�e��5뵼枢%c��e�"8�����ٳgB�k9y#�����.ҙ�( [ �8��C�I6g�� A[��'iw)�0�c�]zb��y��<?k6�+p�o�!*����'���	Rn�$�f��T��2���j뤵V�|��?��[!�����ꫯB A�4Ij/ �Ν{��7?��}=�0�2m�4�(\�`T��K�8vu��
[V.��Wz��9$�0�ha���/�K��;���B�xi�r3jhh����c�$L���3���
����){.�xjU3�c���q�9����x^�k�@���4&VI��FUp	�K�-�9\����uHv*�#f���Ã�Ϯ�UCjٌ��Eo���y�w*w�k���>��+t7o��n�guY�[�S��d\F�j��������X�'Z Y��Pv���)�uQ(4D�ڭ�Jw���������u^\?�����(�����8�Hȏ����k��� k.Τ�9	?�L"���r]q��7o�����޶m�=�MgH�����}�������*�g���*�\cRl�eW��7�p>�_�D��o��_��g>���>v�����ՕW^	�1D�9sF�x���2��4�Ӂ���w��Y�- �F�۰;���[Z_(?�p:@�����t�{�Ͳe���A��8.��=� ��{�z���k׮mk=�+=ov��-1���3fA>��:C�Hl���ý�ދW��7n��00�={���w�u��?~��i�&HOty����"Լ��_��t���"i��,A��͜�;\�(P��~����e8>���o y��D��[�P��ǵk�:�+�VD�$a���)���K��X_��*�@^�3���8;���;2s슲� U�L���/l���rV���6lb�C�9��/\��_�� �������I�h1���1i�.q�%1�#k��A�ݝ�񹱱����������#�(�
�UN�^t����6�fL<�ޡkvwwW����N?a��i�Օ������=�1�J�<A;wc
�J"��I�omE%$	��l-k��fB�d�l��ʫ�������lW�YM
k$+�H���1�j)���7�_6Kj���ϥ�jyO�ٷ��k���?����'�=�k����k֮���3�D����6��_�h��?�_��֖�}-'[N9��uw�⭕�Pf@���%Q�y&�6�a.N�S׬�y6���	�ق��Fp$�a1��� E-F�}�H�y��3��ĕe�d&B�|G��u�:�20L�>����p������4R�[cJ�&x�S�AhJ?%��O�G[.\��"H<TYI�V@�x�  H���ݻ_�Rۓ
�9Z��Pue6��a+��Z?c�t����bO��G���c
���![�x/��a��&��(ǃ�jؕ߭U^����tq�JB��������Ai�)�X7I�5Zy|�����}�u�Q�w��k2��i�^X�4	p��DT��A˛A#)}��|��3
��&��3����^�@�pZ��F������{	���h;+����G%y�� ŁH:CP��u�K��8z�@�F�q��z�����v������2f�z�*XP�4�g�$�\�J'(���6T��T5�n}��S�L�w�щ�Ø8�*Gb�~���˗�ӟ����n�J��S'$Ñ�2ܰ�����U�K^��'�Z0��_E���P;Ν�����J�VX3A�	�SH�4B�*�[�n�%4�W�!��M�T__����}�QL�{��_����+W�,-/�]� ^ [�����{��D�b���"��)_��W����{�_^{��<���$줬,�'��'?����q1 ,�飯�c�p�QAYh���/�J��d�86��
P�l2EM�쌝d׭�e������^�4�a��E�Otr��fP����%���Tj�s�0P$R׊}&R�o䑏D+${�����Hs�� 5N5B/A6�����>�U�
��Tj���X7ߪ��Pԩ&P�/��_aH��A)�vQ�n�y�b��ʍ�kBR B����oN����Ȑ�s�ڛ��H�[j���b�T#���k�:���"i�5�Њ�3"�%4�՘�/t@0��ղ�if�)7�;��A��N�N��hii��$`�ذ$A�V!P�/��I#y���drP|dд�ý��K�į�ph��p�1t��;RS�`u�<�sد8ˎ;�f�h`�<�S�
�������a�+0�p0�bŊ'�|R���O���g��t����Ldsn� ޣh��L�xz}�d���$.|;��ѽ��ڽ~�닔*��WW������'	��
���)�&�^FWjw�H���� �Ks� 3)z�\�1�I���r_�đ܉;�]w�R|��_��Lri�D�~J�} �%� p�w;uꔘc�~���psL�0r.��'{�FU�ʊ�ao������Pɴ�tј�i��p	ht��`��&ۡ�6��C9��#���,�|j�@@��Vd����94�T}Hm�|�c���(4���f���NAu~q�Ι?���DrCUr�eҶ���F�h� ΁�@�n��ӧOCĉE�� �R@�ƍS�(y��OE&������E�/�ph&� ���)���an8(B�
����b�r���[o������A�\�cHQF��Z1(�π�t�����a��
`��	+a"����g���;Q��A�j����ʥ��P瀇N�>��gM�0z�c�=���C�m��o�۷m���K�,���֐�,ذa�46}衇n��x�E���֯_��;v,�$ll�U���/���͙3��I+i��`$��5�q�O�
���1(a)�v1�B<G����Q�>���I��8�b$�W�^�T�37���l��çr���Vhf��0N���$!��6��źe�<)�8�y_1�p}?K�����D2��DF��X������j��T5�ՔR�3�(;��g���T���;��N��Y�K#m�� t"�	"���P�J��6�� ����#Ln�l;�0:�����fV(N!�T?3DŲu.�X�v����v�pmW��^�R�p�Tʼ�54�Z�:���O������ʆ�H$���q�Wc����=���ѐ��⦥��m���[�p��I_;~��+�l������C2^v�e�'��^��h=�cQ�l(��F���Ba�w�t l0���=D/wJ�$閣�d��H(�������KP���̗P�����Xi*p�ĖXxD�g�EC�_s�^��Covt]��B����i���ɘc��F(�h�a	�M��ٳX@���EM�ؔ���QTR��2�0���	��#�I��Y�n�]gϝe�j\��d�&ˁ�b���J�l��N�\��Ԧ�G�@�T`�z_���Z���@H��9�\ݚg���{��f���f��	���8݆��ɸ��x��gd�y���7�^E��dB�r���N�"홋v�+^���BmK4���g3�ؤ��? ��;g&��p|�1����63�(I�oGϣ"ݷ��۹�r�k��� ��]��K �T2��E�O�@BW��)�i[񬆂����f%��t�Ьq�!ĤT������͛7v|�c{���)���ȑS ���'���}*+˩��l[�j"KS�2�t=�H��I�����y~��I�0ӌ��qm	Q�1�U?h�N.K��*mZh%���+��{/tCE�9m:�, ��3g�9sf��i�Z��\G��>�9�����ɓ�Ϝ��v���G}t�ҥ7�pï~�����C�A%>|�0F��3�&��T��ɥ�[w�z���@7ݴH`B�-dl���xH~��'[a�EL<������G����,vȶ����6��.6!�+���}���nm�9���yN�������<DS7++��9������;v���1���a�0�׮^�+aNB3���:(G��.Ֆ�(��V��a£�HJ`6sc���Tj%H2u!z�_� ��3N�sE,	;����+�t榍���//{,�E��Мd���<E��0^��?�̓P�?�#2���5�_��V���.���P-���6���j��,� ��(a�{��q5.%��U�'?��ѣGaF�x�8�tU$��4������e��5{��0�*R�!_�J�#*!�b<�
���د�E��Q���'�&��
�����]6�&c�4^s��|� �y�
%��q�t�M��7���xj}:�}��Ξ^��M�U��J�*b�uc�@��Τ�	�6�%����֯]�e˖g�y
�])��B&b�O�:�q�k���,Զ�k����|��ms�D04�n-�O����@�<� �d����t)��z��c|5��keؖ	��\�>|X,T�>�G�|��o�	
!K���%�q����e�����z�U+@J�@�gT��d5�(�?�8������������K8�Xj�+�),&��T˄� k�)�*dddD�T�ɸ��&Eո.F����� #G�pG��#F��A�)�Y�5�0���ia�l"F:���(W�eh�82u�:Z�jl���֑�U��_.�M�7�xc횕�_��V��R�ER�b �!N�xl��K�O�M�K#Qy5�,2Z)���!���󅒴[��i�{��Ifs�dhkk�̀��#d� ���L���L3��@ǗI�ep�L&K��pӋ�H ^�h�ex�3�<vÜK����W�W8#���A �C(�ىӨC]�B��۹�'N���"����e%�S������"M^J�y�,K��l��� ����1� [�?����߱y�����!4>����}������/|��Wu���]�v�W��`�A��?��?��i���?��{�;vlÆG����,�]0*���?���~V���C�*�N��U��K�b\�ŵZ����󥨵h�y���_5���s�/����!5}��@[���0���	U�Q���L��r�{s;E�Xy֙��&EW�%��dR �L���g�9_�$�
�h_�T)Q��ӷl���?� ���S��J ѹ*.�J�c�驭ۯ����v���鱗_~��g���e�IO� �cȘ�	)<N:ɨ�	I��+!�X�P��'N�Z�|9^frz*��.������W��7���$W�v	ո���e��*i�;��;G�(`b������9}��>F?�;{�f�Žo����]�f����!�I�?��Q<�,�Y�S�06s]B��s�cG�oڰb�2�1���k�z��%˖l۶�'/��^ZNa�~"p�t;pL;�U*� UT��3�6z�%S~G��`n@�iđ@mYH~����4/�.ȣ���.��+2��f>��B�2�e�����1��K����#'���!T.Cg�D�A�aqϟ?/m$N[�8�Ȋ.����+TS�%�;MUWB��u��R�g����)�Fb�ؽ��Ny����	8���#u�00��8)��c�5�z���3i�_
�G�i�HRt�lb����g�~$�5�͈jA%�AP��`���c�����ȗ8�6[�gt��#�M�($����s#I��p��=o�qÍ� �.X�[e����0}�Ӫ#�g�Ni��m{���HW3�H*\����"!AZD��a#�Mi'ܠy�1+�����)�W�f�Pj\Q�-] �!�attRb��/��/����7�8�!O�8�LR�=lT�V�4�+�H��U��h�T���"ޢ��)�> <�\�����M�
���\U)�Q�fXc�:�k5
��"��֖�
��� g fH] ���Q�	��x`Ŋ���������o��;��o��O��O�{��P[�j�1&|��ݘ��Q�����O��?�sgg7ƀy D�-��m����ϱ^�@�5�\��o.�-~�U�^I��[K����	��
�n�݋b�+ղdo��u�J�]��\��c���ָŢ�mXT�E�����t�����C��(��w�"�X�d/V�nG���p-K[��;-��3����c2D���.���1j9��ʏm����	�ے��@t�S�df�3&�c��^�A��9:*�6R�9`��y����,]J1����7��7�R���^9!vl�A�u�ۤ$�)�+`���X�=�F;VC+���RP���q�H̑��D�َ�IQ��Lʘn�G>�0*���g��5�7m��;v��lc��$Z[D�1�n�ԧ𛊑�R>��]�zN&b7d,��ͽ;���	k;{�,d߉c�aJ�7�3�LQ��"�8`b���.��W�B_$=*5�<!$�m%q%6��%��a(�Jhx���֓�#*Hُ64Z�A0]��� .�%긱j���ڨ�Yȹ��I¹�q\��B	�c��LH�Dr��2>D�Y��f\�Bug{{\$SjP�W��A�T�9pW�+�Q�	�2�U�ZiAfF�:�Qd��Ǧ�a�W�1psq�;�Ѳ̥���cU�~	u@}�øf�=�ެd�b�e8�#lZV9o{�i�������������_���#�7q�K����C�,��u�����B*$cq�E���e��T,��[,P__/������
�Ў��$0�̣��be%E�̼l�z�	�01J���rG{;��b /���8���� �����߾��/�={��oo+�
(�(�G$��Ed��1q��0����YqHvd����V���Ձ�qw�����(R`+uAh��>��$:v�8d���گ}��_}衇p�'~�����;>	��w���0�A*Ƽs�N�������W�R,���.^���>��_u�U�|�ܙ��A"<(v�-��K�ȑ3���ɸ�UW�#��B�5q���#�_�ieԽٷp������V��X�s�?�#�.�}eskl�J���Ѯ��t����[7z���['G��`��!�h�x���{�ǣh��O�u�����NS���6jz�#����bE���ĵ��K�ׅ�?155�Jf����J#�o;B�s��\��ɭԪ?z��G�ܽ���������?|�@���Js��`@���/�� �,��&7�����ʤϚ�⌍NL�3S3yX6�7��N�3�T&,R(��)p��Bm�*�L���q��d�Gx��i'�0�n��}��/��K�[ܧ���o�2m�|���K��4n�Q�:�ū@��4��/?N�@���7����w����ӭ�;C=z ����@r�BݮڸzG.���F�u!SSV��C��*Wh�p:�tA�s�<DP��J�.��Y	[h� �g���l���$��$p&2NNH\���DN��d{hɔ�\-����kr9���]#�����)2(�]��s�w�rqd����z�[��q1W��N�V%P[1��������J��H�j�b�99)����h�Bn�NDQ mbb�ff�BJ�L�NN�Bp&Ȭ&q[�zZ�^�ٳ�@������Ud{!hn~��7_�u<) ̌I�`X~�|v��Woټ	lb�!Ϗ�,�,I�ޥ��iޙtޢ���aS�ҩZrX��7�]Ȑ�T�[N!�J�	~��[2�U�^�l�xa��)KƳ���3C(����Q��,H}�t���/9'Z�f��?r�n1���}�/��/�~ Ź+<�+��M[MW��\����s�kP��0!�¼dj�+��L2����քvl�
��)�j��K�.��vfZ�f͵�^{�4�����g���}�������K?������{�}���W�߯�$L,�-�A�G�^@f��ԧ�n���?�1漫�J���]w.+�L�6S�C��w���� 6n��z��~�:o�i�`DH`�tRm�B^d	��������B��GS_]�K�ybѸ}e|"�ڿ�Y�7�� �sf�7{��]޻fK��8�6^��/��3OW�R���q+>3�vp�밆p�}phVH
c�84ē@pK�#�
�xo���^a��'�Q�b&�.�z߶�qmCW�q�u�Xi��m50�w����E}�s�70٧~��|��]1��/��/$���_�D0�aZ���]5<)�	c�G@�� ��W\����&$�� ��8��<%R$,�2��d�~q���y��p�(���I�b�
��Y�]�]x\[�m�ʕ0� U��GW��9��^��Y�uX�>���R/'e��k׮��������ܷo_-�1Oj)��dw�c�j5��L��+~��9��Z�5ȗ��,M��בd�ɮS����z�`٥�&k��Dz�D#�#
S��+��e1�P��F�03��b�H�GE	�����!Ô,f^���j֍"�A2�����]4�/���M-\A02��l�W��A� 2	��cA��=n�))��j �FazZ_�5�8t��r��+B�{,�>�T|��8EѪFw]��S��m�af��Ǧ��|��޵�Q
�e�fG�X����F8�q�Li[�J�r����������z�T8��l�/������Բ��}rjv�������Ii��P� ���cc��c��,Ɔ�RcRo� FG��.!�[�Z�\NQ�n�+6z�sϜ9� g�&� ����\��H����f�%���+�vY�Q\DD�����	�@H��rf!r'c,G�7Q�bɐɴ	�` ��� J[�~���ǟ����t��A<�ӟ���O?���|e������K Nʕ��Js�Հ�?��s���1�����7oƴC��0�5�v���x>��nܸ���^��O~Mz��� [1i�0Z�_�a���CK1���n�ex�.�B���+Wl�����n���#�1�W"1������<��PH�)R-�2~Zո1�D�+J���x�TVփ������aФi�=)7��e��<zl��C:����jP����V��X�9�3��LPS���2	�^�\�ס�׸�bTq��K�sՃ�j��U��E���:3�[����[��Dy.�N� y��Ly�\`Tj�湞��o�9`���;�q�Pp����ЩF!.��A�-;:9*�p�xC�ҿ|��?��?����������3�������a�Lt�<q�4K�qT*�s�3̊J��Nf<�%���vO?�+o���'�x���#�C�TT,�X��3�SR_�B5]*��r�J������r�(���R�W�ڻ��/��c*��׍��l�T��T�:���-X�߳(�)��T�Z�)���+K*�,JI�U)5��|�k=��prj���c�6m��i����؂8`TAI ._F;��*�Rm�Q�Jy�Rٙ�97:J_�p�q�T	�U�WSlV�J�ZC)��ٶv/������T���%M2��M���W5�?A)��vUeTZ��6�'�$������#)�H�vsj����3g O�Ύ���$�vOW�C��R	ן+Q7t�L�O%Hy�OO�}	��/��e�(&��S����d�R��F홤CqWjv��^ʣ�$)HtݺumT���u�9~�tL�����+��&�%�6�J^q�DGWw�R��2Y���Վ=A-h�*á(94��LVj�us�c��-[���ر� �	�&!Y�~`����(�!�HЈ2�C�|�Urm�8<4�c�S�T��=���\��e�G)�n�C"Ћ�jD��b:)���ߕ�Wj;�X2Eku
�n2q� Z�0�Q%IF�AU��J#>��h5*4�'Q�aV��gΟ=GNn�G�I{YqQ�
id��EB�v�-��D�W�����J>�Zk:��0#���W(��a�%=�X(�%K�utt��{����G���~�˾����_\�v����_zig{;�������@��W�䰃*�=�e�w���|Q��Z8e���� ���/�Z���=vqljljժU�m�\�����ɧ��򗿚��+������}{��?/O;���#C��&����l*���H�o�e\*��K��� �hG6�ue)B+�����A�6�N<7��>���dɚ��J$3S3�r������J'S����<bv�	�#Ï?��5�\321><>6�d����1�+V�<y������u���w�'����z��;�����k֬y�G>
���SOB'�$���[�x`vvrzz|�Uk7�{�'����>槒�p�nWo��|��0U*e�֨��̳_|��������9���l�k�*�[��g�:�F��:�#5�MB��W�B�R�3?"�Ip��g`����u��q�^�j HMJ�Nd7����cW��U��D�oI씿-��BЮE�"�'=b��,C�#��1Q8����q�d����g,���u{��������t�IcW��1q�ƒ0'���A���V��<��A�E5U >�}=�={��õ�^4[alb�t	u��7aM&�t�����.�B}�G�����on{�;�m�v���og��>��B~V�LS�o�]��ʌ8�)�3Qb�I�i)+%���"��8 w`���	��(��Yq峄C�����31���M!&-����v���d�P�'JX�К[�n=y�5��;ԪqA�u��pI���A�.�F�z۸n��+N�8N�(��q����t�ةR�UXc&Rϼ�;55)�̩��2M�a���L����l�Z���in�#b��wq�B��K2��2�d�O�b�4�d��8g�}���Z\��r�*%���*����i�5$���@9�&���G�[�5���z ���>��@����j�ʜ������)�eb�	�+�x3�sY�L{�"[K�U�x���:��J�R��sAx0�df�-*m��D��xg��_�tE���q���`��5��y��S�g����i7ܡ.�.�_"�t�N����RV�0��A�JT���hS��Bp�Y����'��k:�d�;�kHV����O>�$��W8L%,]���[o�J!;v�ԩS0q<Vk@� �|>/��`r�\��Z�%v���n6�#HV1���58����M���".�vtd1p
�tC��`//Gٲ���
u�8.0��zl�d�O��aY�(���ぼW�e��\,P�ҝa#�����hz����/��իO�=u���%�B�/��a�<G�<$�`۶m}�w�q������3π!�өԖ-[��W^yE"�GFG/^,�·O�J�< ��կ~�x�UWA`-p[�?�/�!!a3�Wz�ffq��u�IJ��&��� �z�r}�����l޷��m��?�i��.]v�*��tv��o�
K�p���w�����iu̵��y�����S��;��@WCP:k]T�pq*2�[<ۺlo"H� ��o�P���H�Z.ɶ�#�i�"�����(�X.�\��w͉a��S�8�l�K�	i�[A�|��߭V
���g��/�f˵�����>?9=�Lg֬[_*��}``�:��'���T�
�����x�Y�g����t��Q�C�W�̀�H��aoW�L!OV3�ī��d�����߸N�ϕKKڲ�Z��ݝn�N�LwvvA^�\x�M�r��E��óax��V�@�5(ĆD�{1#x�U6n�x��!��Ϭ��E��y����,'��\9
�]>3�����8�^Qd�U��j"�&6^�x�_���oBi����j����"�[z�n����T�ê�G���ڲ��)��Z�8�#�Se^�?L̙$��� 4��e�H�n��hI��y��֖�HG�U�Vtuu �AX��u8���Q��������bר�}!�U�N���j���(�X�k�Q���*�xqa@ٔ[��P¼��zUY^|W�˰'�
CV�J9j̇�?�i�+�2DV�1�o�x�g�I��k��V��I-�þ4�P��@ܘ\��aB`m�vK�0k��rE��L��؎��-��goU{��66\׹��J:�qG{%��N>W�;@�����r��:�KwQ��]w�	�y��	6�8\���o�i�}��l�*���;~�����_�J#����`��}3��!�� ?`���鳀 }}��xjdl��ر��c��<�ů@���.��qc�z6y;1�#�ё�J�p�'1��Ą��P�믿��~�{ߋ�x��^z�_�W �ήEڕh@q^E6���]EJ#��[���\�|bj���:�7n Ą�dy��y�j�h��|��[n���?�>�(���ݻ�偽 �?��`Ν?O5Oc���o����{
�T��ԉ��w��`��r,͑#G`���4(Eq1��QD��Z�
5Z*P�rHn��Ş`B��*�6>��U+8�a�X#~��j�`�e�44Ao��Kйۊ�.��g����u�a�GzK�ե�����+qQ���(�1:��D����ZF�-���{3c��	u�?���%ƨ��X���T"W�Q��4�Frq��yG��5A$!b�D1>�W���@Ҿ}����o��+Hq���[�&}�s��ܱc�6��m�i��S���fE��� �+$M�;���V+Z�Ġ����L�uu�J+Sd}�P�`J��-�X03ً���D.dD!��g�vR��i�#��f��,~���0a)��K����6[��	��z��GF��ΒXg�.59�xڏt��	K�*r��\���K��:$�2е� �`SC̉i�����*�������LuJ���Hs�m�;(pM/��4��U�t1'�ϟ��7����(P�c� gA'P�����5�%��eP]\o�R7���V��H�PH�!�o ZЏ�Iұ	��8�D��n�ԗ�ԧT( �hJ�8�r����J�٬N�W��	������������H��Ѷ�X1vѶD�Y�Z�ĕ�˪e��>RJ
�5�J[{�#�m}��ݿ���W�;xeqw�Y�[.D.0�FuJ)5JL�.w�|ްaP�Ν;:DE��Յ����A� �|Ų!�vժU�'(w���Kn�l��	B���"M0q����/���(���s!�d���f�Z�{f���ط�;��$f��s�J�97�����l�(L�gI�,��
�D��lZ�`����=.8����h�ө{�*H���2쓦G$S)H�	j�L�u�
E5,m�ⶀ����1���A?���b�@��_���;o���?����ro���{���7�x��'1�f��`||�n��n�ᩧ�5�1-+���Xgq�.���gi���oE�Ca�����U���J����	�N~A ��64����LP�!��J4���ø���꤄�M���I*�T���b&��h��-0�il^�ZLL�qg��2G�SՏ�.�q�����>cP�{6����L,ey����il3�U˥S�N��a�\ys�>��#ɴe:{�'g�SS��[��H]�r�*KO�����]��}���:;ڻ:��F��������Է�C;������7������>t���v�T�yN1�P��J00��-$�#���^64��s����ʕ���cɺu�XT]ܵk^�CA?�҉d�--;<�5ĭ�^2�9q����XO����JQ~&%X�M�z��]����'��dBt$�B�qUnޓt���2�~���	&�ס#G�>qk��&���Y 3ll�0��Kr�qWl'WM��0�x���nV��\N���4������*Vd�N4v潸�m�p.^�gӉ���jWW��˟B������i)2S�|R���Tr��v��!`�U�옌����!�V�Iχ��m�L���SV�}`���f�E��t��3��Fq�M��@��	�(l�SM�4�Yh�X\,e�d���Au��T��.[�r[��a߶���N�q�q/��L#Ĺ�e=�>"7������od�o}z`ɸ��e^�o��J�i��ti%�b����cGO\�am�\Id����Ԉ#l��yW,x�,d֪��V�Ui��Ǭ�S�'�f�\}a/!ߖ˨�v^�h���m||�̙3�d�>�~�i,�M7���7�	3 Ёň�:��O~sw^�? ����W B�4 0�+�-Ί�m�}�:�m���g��I���5�IZ�U���x��+���۞>}:�D�ďOL�������'~z|�bq����͛a���c�(�|�"|k�,Ɍ�\.
j]�=�%H���[vi�;�9�J��L	)v¥8{t������,�m�z�1��!�ggO�<i�|�2ߧ����/�}�݅����>z�7�\9@&��h�\����ҥK����\q���k׮�$�^��'>q�uۿ����>q2?=�'��0]�ܖ�u���t
�g���=�@CI�FU�b�R,A��=�Be��te(���k&0|s��.G�����}=�s��E�[�a��[��>��֌�!����*q4o�8R�V(C���y[�K�|4ߦ����r\�}�e�#U��� ���#�t[m�ĽT]ݓ@b�2)
I%|��1�Pa�������'&&$H�%�֌�G"�j7��8F�h�n����A����h?{���?��O��o���~��������=t"�M,[��)��}�����;��8��B�ឹN�r��%��������b�k�:U��+hw ��zx����g��X��j��J!m��Բ����{�0��L��A~-)��|r��)�(f1�$=��sY�G�J�g7̥��̉���gn�z�	����ZI=���+d݅۝�t[3�&p��F�� "�Eٶ#�f�ę$nK��
�̔wb��+,(*���9���� ��7�\�~=^�P�p�c��@\�R�bŊ���Ǐ� *�јR�U�ɛ�¶u獞O�pW��xp�XJ�3��!{��JX���B�����B������ԅ<��-q�&�`��A�`d  �Њ0��mL3��, ���ǉ:�ۀ�؏��Nb��y�rA㮇�Ƙ�`P�\�d_�s��"+7�/�1e3�je
u�k��P-�e�o��c�1���T�j񏌌H��_�׍U��׿�Ƌ��8p��s����D(�]�� B�^�d�|��E��$�8Y1��U�Va2�9L[�i���I�%�k:��v�a����`�q�<�[�T�#��l�N��������;pfr��vuQe�J�\�*l�o��T�n�<���%�@��?'gy�e�Y#��]WZx��!O��V�s���[��p�0":�2W�l~bǎ����w��ݏ<��}�W�, \\ �o�!pϕ+W�J�_��_������tS��`HX)���l�M�p�u���a]�D�cGo�7�3��W���f�S3����&"T�nG4�GY�ms���-Hn�k�����JDQ+,t"#+��1��������EO����1v���_1�2���^���/-�%���-���*]]I�	)*��R X�
J�X�BJ]mTS��j2�Y��ew�]�T�[PS=��΀�;Kuu��:s�g��z�-�~�ؓ۶m��~�?=�3َ��7���7=qbٲ����h�ԍ6����Y���l��<wh��^�����{U*�XIf��^���uCb��(��Mc"2	Xl�ZЛI/_����+TA�T����3��$�\*�j��n�J-Y�ޣ�r��|�Ҝ�f'rCp�������
�3B�@,_��"�Nz�f�7�\GW������U��h;��"��Jp��t6%u!M*��0W�)y3�F6ÿ5.��4�f^jw��������m2�2�(PL�������$�!O���^��;:r��Sc�'|,A{���3!L/?L~�2�U�|7A]R�2�z *��Eű�)�+�΃��B��\}
�Jh�@��Z �
�\N={�$cz(�v���Z � 2��	�!~)׉1�x"O����f�{PZ�ۻ$�T�מm�7'�^(+���>W]��4�0��c�	/���v�c|���:���$�xN��ƭ�/0��V���6�,(3S)W)���,o��xl���hм�S���oEطZ ������i�Xż�P�=�Y*�:{w�%f�(�o�}�����E *��/�r��W�g2���I�kKֈ`}iy(��A��G�kb�Ž_S�t�Ob�A-��꡸��|-�/���ʧN��57������9.x��i�!���a� ��coj���bG��H;w����.]�����ڵK*���Ig˥;v�ڲmkO��-[��4�B�R�" w/	ր}��k�{��%�.]��fJՊ貣Gc��&�0Wz�Ă�1!X400W���m����~;n�iӦg�y̅��G�AՀ�#&��s�ش	k���L�ڡ�~�i B��'?�I`�'N|�k_ú@Kb��XPFc\� j��	~>*�+��5
��`!U��J���I�C��8�Z�h���T*gl#7�.�L9��0v���~p�#���Y��o�G?w���T#�����G�8q��h�J�f9B?���ͮ�XuZ>l�d8�ޕ���:4n4=�����5�mX�ulbf�&��&yԸf�D���\����8�!uM��W0����1������ʙ��Ô����G� b��_������?=���uk|����F��c�۩���rH��xI�@G�����F�:� �'�EꚮQ$2�b���666��rb찁$jk��Eؖ��ٳg���ЙB^RG��x�"dGF�!�$y�f�K2����xs��_}~j��JE����R�����Z1��1�&8��)�}�(dJ�%���-̬�]�cy2�lY����E��2q��i����N��Z���)����)+"���*U��*@�)�+��,���o���\��r,z{��pR&$��O�J�
� ���BB�����
a�D�F(�@�A"�B(/��:��i�(.�I����� %~����>'e𦪑l��d&�6���B�2Q��gZR0E�G���:��?�5��H{"Z)mR^bsS5
��{ƒ�����1�}����,��e'r^���R�����B�W�������e�ڄ��I�֤-:Μ?�����6�X@ gX�����}!*]n�4 �N�����2PJ���9m�F��"]�Pl �ƙ3g����tK{��$}��}���[����o[.�~�����?����o���Q�ޞ>� �K���8�!*�%��~����ԧ>�⡅�,ס��j�Ѻu�V����N�:*����p�􅴍� �l�H�[a@�����DI~eEY��`>_���Pr,��0�Ύ.(8����_��G!���� fa�p��7�,ۚx(&a���R[���k~��� ���_�F&R��^�JI�����r�0Rq���,]Y����|��s#��mBruQ.��t�jhߡU��I����K��yh��Dj�����8\ť�Y)��"�� �FǠ��f�Runc�t]Qy���Wq|@�[�H1q�c�)����`1GK@'�����Oǋ��yRf#�E<���.`����\�=��B�~����,Ȕ�PW ��U�ģ�� ��O+?ɣMĨ��B�
�_��:ڏ�8U�T.۹{�?�˗~�c�^���޵x�2�g�}��*U��eLl�d�M��M�V,?p�`�@��8��"���E����x�\�+R�w߰����ϟ;wa��U��X8226;S��b�1�?����3��C�i?l�jժ(������ܵ���/X�+��ONL�VB5�����Nx-���l���ɓ�U�\�Β�,�AZ4�p�����#sY2�:�ޫ�/*V)�r��:;�F���q�H�xWo>Z�Bb��٤^�\��G/�D���ldI��o����Wy;���&���05����2��;Hk�ye�*� �� . �
4��,.�5���N�Ŝ��/��n(��RB�Cjsaw��j:Cᘳ�i|����0�]
�T0�����▣�O�pD�éj!���L�b���t�!.%�E�=�Ǥ���N!g�I�2�[�3�̤��.��S\�O�fAP/�����o�篎&�8ʅ-��E�V؋ӖΤRi<��Ŵ�b�Pl�m&�T�R��H��l	��d�FX����cl|bdtr�u#�g �%(^f)�%5��'V�x�w?ԡ�B��`�p�UF��&](jq[<'m��թxrw;��U�0?��L�
�ޱ�� FY
� 3,RQ��~������@a1p����g$�E����L*�h����x�+Ɍ�V�z~2���?����{w�k|�3�9z��q��ڵ+�c!�;�ɦ�	���l��n��_��Wo��Vش'O'L_�zg��,}��w���k�o͚u���[\v�J��JY5�<�n�aT�6�Cۿh�l��v ţG��侀3W%$�ٞ#ӽZͦ���33܀�w~�s�c3��O?�&�n�馛��>�y�Y ����-�p������z�@�҅p��1�0�'8O���~7�ݽ{7p3��J�24;�A~����0���\o��x
u��Dj������_b�);�AX���9�Z5��D-�$�o;;2$R�Rn}�>=��7� ��R��k^�6/���qFSH��?ݨ9�E>K�D"�v������L����IU������� &�~*��n��A�Zi�H
i �و�f�h6k��GQn}K"��G��0�V���0�V���w�(i"N����#�-����?�h�b��G>�P�D�v��B�T���о���У��#�G�������9N�P(��p��}/���w�~B�LaD�XTH(�'�@��-���0)��Z5�jXL���o�A ��ކ�p�����6�ծ�&��3��!>8P*橶����DҀ1{�e�������G��S�'VY��d���
�[�w�^���a�e�h=��P8�o�����Y������= `��JI��]fCЕ:���yp�dE|���ND�bA"�L�V�Vwu�B@	X�G�����&��ɇ�KƮb�����zM5:��L�V�M'��3-�b��N2��{"1o]�[�r׬���6�a���o�mr�OFJvZ)P��7-z�"{��n@�ѓ��� K�U���Dz:��ltqIJ�9*�{�4Qo�bEoݗv�KW�}�����M��K�����V���\��	�HP���\�<�t]L��2TN�R2�'"v׉䇸��`.цf߿�
���+��1���~z�����{�Y�x�]�zzz~��{1��}�c��������P����9z��	I�?�H��%����_�妛׭[711F޾E�ۛ7o�\�d��q��JS˙�q���Ҳ��s��|�;���Jv����o}�[5j���U|)�Meq�J�y
��|mI-�L��;_^�z�֭[�����Nb0��`����)�ꫯVb`��<��?`�~��6H�)^������/�t|�\�h���Q��R?�S9t�ʺE#\�.�Oc.{���w).(vY�_8q�{RM���Zc�B��Pz�U������j8�Էum]�8�j=Dz��x�{y��%I5����څԄ1�ߪF���Pᾠ�(�X�I|L2Mp�L�n�8h�Ys��D{ŕ�aۑ�Y1��d��R�򭇿����	��<� �R`���HWNc��%0�+�!�ehg�V+�����w_o~�/�3m�m��s��!X㝝�J��R�N����ρ���	�\�;��B~�"s�{ 8�R���W�>yW�LM T��wNMM&����~)~}&&iAA�2�p�b�*QGT�#������'Wl'�l��d\r����d;fq�s^񐺋�j��w(�U��\|����^xs��e��&f�Sh��������;�4l�D[��b(��k�/����Ju|�RNv��if@'�H��l,��%��m���'��J�H�劤�cC�#�)���M����{���X!ʪ����T*��e񸙙)	����#Q�r5�Z�v�fC�:�rD"�o_� ],þI3��w6��\l�أ�5����B�$[.UE�gS|#�0�B�ճ�S�O3f^�3��G�Ad��7�i$'|=2:]�����fO$�	�mg�:�1Ǘ�m���^Tب}#���j�j:���3��N�vw_s�����<�q�W��#�1:�y��Oq�R�X�	?�!Y����x����:��Y0;;q%p|��E*u[,���\xqt䟾�/�+���C������?��'>�������/ }�KQlܫ���S���ga���� b �`�lٲPoxxX�^���M[�\�O)U���/�ʮOx&���R�x�;�%Ԕ���lQD�e�s�t���-a��#CCC\��� \/����l:E��D5�I64����\,r8t#\�icw_ot�ę3g�gg � 
�
�n��_���Ƶ۶�x��=�$��w�-��ݻwC��fo�ڵ������
�L/�z�c�H��D٠��Θ�y6޲���(4���Tt)��+u{O�8h�Di"e��H��#HYď��8�����3M̢�A�q	�\6�,��4��i�����6�a	��c������%�CGW����]��g�u�P��K��(bWNr�M]��z쬋-{'�=a�Oq��)�9WP륾5ݥB~�Ν����r���?��c�v���l 'nx �=Rmy��� O`N).�!c󹫷�`-\�|�P����Z���d>N+�bB�*KA`�R��y�#��lL�[XQ�s;�� �$�d��t�/Y��CQ��#%16�{FJ�!�,v�0��c��ơ.@��q��)��g�a2r�m�x����q�B�!l-d5��Qt���6����R�SBmFGǡ *�P�!��U�i����>5Lq<�����C�&:���l,�C%О���=���P?CCKiúZ]�t)��4�t9�W�/I�c'rmr,���M/�����8��d]��Yj�[J��@W�����n�ϔ�j��j�C��eM].I#�>��d�s2��R���1/n�4EnI��Vb1$M���J1���۝s���X����4Ɗlm�jT���W�B��r�y�i{@n�*�aHM��E��!Q�s��߱D"�c�21t+���D��w�n�"��H��L)�ጹ,yԸ�d ;�@W�'�|�4��%��O>�X�}��;���>������׾v������m۶���z��7>|	O�I�ժU�e/-G���gɩ�y��o���G�c	#�┒ E����k�I�v���Π&�V�$��)q-/+�k�dfϞ=�	f��?�14���<M�d��ˈ���?��u���ݤ��X�"^$�����D�R��,�$���ZIh.h������tR߭�b����=�i�&is�yɸ��/�e��}�^L��rct����>h/�A\�����|ȷ�j�-���a{��}�)-pܵ���*4jXK��&9��f����Ȁ�aT���\.���l�� � eә9�>�ǉ$F(uG�e/P/R����Ӗ�)V�K%}<�R--Y�W�?s��-C��o���K����|s�ܐ@R&K�a�-�X��n����ON$R�����ŋ����Gʫ��)��T2=;SL%��W56\X��e�_��ή�j�]�M�����<yJ��S�n�I*����,!�8(�'G;:rSS���^ ��'�よf����Xo����W_<�!w㔼w����=�[�b��0�M���"^e����Ed�p�w+�
E7(�H�A-�7٬�[�6�Y��띬�x^NEk�7��8u�$�2��@��+?�/J������R*�
k�Kk 7!��0 H�P�|+�G}]{��;��}}=�(���T��1߁_�S�Zٍ&�i*ZE���ĳ�Rg�ZG:�I�dn���&	�~ՙ+��U�c��lXh'��j]_��x��q���e��!bܠ��'���Qj�I�#�W��`����e-866�|qt��%~���nYK����o�H�
�&ҹ�W�o.����A��m��$�O=FE5� ����ٷ>|��=����B���I[U��w�ѩa$�q��,3Ɖ���Ia�i��rO����&0B!�:.׵����c�**�֬Y���Aei}�7�x�ᇡA����ҙ�wܑL�o|ϭ�d<�����/ s�>��ŋ���,[:62���簵�V�H�D:ә�vtt�~��./9[.LN�T�A*����K��������~�)��3��8���=J�$ڲyk_��7zxzjV��q[-�tQ�f���dL����� 7+5��Ϝ9��a���ٲR�Ǽ��W^ye�ʕ�Ν+��V�[{���5*u�toX�hs �n�:����⶷�hJQ� aC�� �=��gJ���0�-a��c#�&���[Hn('��k"`�OM'�A����5Z��;�<"��S�:��փL����P�	OoВ=��o��Èǲ�E���l-��m�,E�\�xOd �8iB�s�J`���in#���U�L��?�|��r���J�����
�3��:{��믿~�wvtf׬Y#�8p����4���k�8g˖-8�bJ���c������h"�2\^<�>-W�:{�44nP����%ө���g�sP��r��ŋ#Q�L�[@N�޽{Ŋ��N1�p�H�l[�q+M�Iy�\�Kͯ�8��0G�.�U'r续c:xH���zf�gt2i�){��7��h�;���7���9���]⤭$%�:�>)���.~�J����r+����!UZ*�� K1��BDsRЖc�e���<4�y��| �{�^\<::,�� s�-ź��'�``2�q}�Pg7�f��%&�@(��U*�6�MP����zV�MZ����F`aK�Hǥ)K�^�3�5P�_��d~���4ܖ��b:��&�h�{���XED�$�ـ��i���2��J\����hꊏ�ů̃wtpwl�sz]�>Z�՚����@v
xe|&<b��h^R%LyW��[����-�$�|�>y�����YF�Y�ɵI�@���7�E���%����|�����{������T.w�5������W_~�����x��YJ���Q�
�["��s��W��H-��"��+����]�!����[)A�3�e�Zx1_X�d	.��|<�H;�i���@`�ÿ�/wתU��.[v����>�@��;w9r�+�_���g��Dz���>y���7�<22"�B!�\�۞�X�ʗ�|u�i5�<���ir}�\��>fc�>G��#혿4Uۢئa>�l�_���7�ҿ�����2I��&"��v�G�@��%F�OѢ��.qf�x���3����A|�rL�nˡ+�p��d���Qm� RA���E��f������j:���!�X� BE��PT~X�\%!D����Ӑ�˖-�:��`�6��˗/����c�t�±��R���8���3��.@�S���LϦ��H�U+V�x��
�mmp���e�R�L"�����{{�W�^�ʦ85�:k��g��/]"UH�b�-+֮�Ʌ$-��$�҇��FQ�����+�B�P}i$�J�-���8T]1��z�ި3�>)u=� ��N\�_���٧,>l%B��̿1>��XVG)�o��/M�6�-�X%k�3bH���jn�����v�29���8"�ІH�8o�s���3��MD%�L�p�9�^W�c0j'�z�!�b����0$`���PHr+��@U(����ס�cf՞�H�9��4�3K���|k0�}C3���yQW�2I؋��.yxLT���v�
MFQ׼z����:v4}�犌�HDWY%(V�Œ�%���[BT�0)�����-��33��'4Q��qYjWC�øNKe2�D"935���:93y��a)�'�a�Y_��f<�(��z�f!L��m���Cn�(�v��Ij�ԯ��2R��+Q�R�45;��Pwi��L��$u��g0#�,�_|��ѣ�:��ٵz�����w�|��90�aÆ�%`�i���z�3�S'�Ps�����]��N/������̤��L�c��S�N-]��|rj&�yCˆ��A[�'P��7�ŏ�c 6�3�� T#Y�t2kJq6���W��Jڇ�]($�s��q7��q�&LݦM� 
|�?�(��[o��~������M7�>������������?:<�_�k���b�TߦS�G���q%��]}G�`��&Š�q�?T�'t�L��&�y	X¥�ϰ���w�S�,;�*�ԥ����rB�X$�DSI5��ץ�h>{Q�$��=�]��ً���@ɖ�����V���ٍC�c� qH���L��h�h�6������\KV�ڈzÿ�ɛ����@\�~��XP*'8�q��	3~�T_�8~:g ����2J�xld�|fE�A��r� �����sωՈ��-�����������G���۷��w�O|�������Ha�7�Q\�J���V�s�Ы��cn2�jtu�k�2���2�,2�RF5��&P��vA�`�(�#�˕�#��%O�;���vv�dh�p�3�_l�G�� XO�Ҁ���I�Z��X�Tu�Ҟ.,�r��@nA)0 �����H��1����P$mg.^�(bu*�V"�GK�g�A�F`dC%��Tu�r���37�!����2��sb��>����7M�z�aP�c��;=�����C5U�
%\V��G��?��_+6��,��)�:������$?�}ٷ��EwX߅��Ey)0���t_�ҡX؆V���}{�pm��NܶAC��eR����K��Ui��r��g�r(��3>>�nK�Y���vx������
�r����k���I�3X�g�}����I?�e˖n|'w��~��|�g E�����������ǯ��z���!��
�F&8=�pXGP�ᑑ�{�>����'N���]ݐ՛7oƿ�V���H-X��,'P�66q8��pK���MC�C�{\�s��:t�̙3x_���m�vP�l�ڵ����O�yC*	$�y�=��Ϟ:�r�J���̔uje���>�6e��X�}�mM5��7���Յ�L�y^�Bŕ�¥�+9�d�}7�c�\�k\$��/��n2y>�l9�%\���?�q�D��V��͂�	��u"*����uY���R��=�q�-�؅��WU=�__9 � zՂb2��s����@��}o�23z���p�.�Q���3�Qܶ�[��������\'�J�lM$�(����^R\&�D�s��T�5���L�3יN$����A��
�<eG�����w�x=�͕�����d�\ݷo?�5*�Ta�-Z�$?7�)�^"t��Ξ����>��Q�p��@� x�ر�<�ȱ�'�����3}	v�UWm߾���Kۺ�^}�՞���%�T�#�߶u+��{�����~rժU���$gN�]8{���ͩdʥ�p��E�����CS��`.��Q� ����k3�9��<'tc����α��~.��;��
.��S����ZX�E�Z��O�G�i?�����JI'�W���+}.ŁB)�J���`J����RÍ� L����ʠ㜵&�*��f��%��D��i���cEνF�ĝd"E33�מ�[֊�Xɠ�$���~� �I0_�D��T
�����$>V���*ʉ���H*"��y������)gx�-`���ꍨ�f'lo�a��
�H���*̞�V�Z�ҳ��=h��Ea�I��J��'m����Z�2��#�[��W����y�b�;Ա\�x�D�5
���b\D��Z��3�g����dʶ�ż'���Y�P6�Dt�g4��u�v�.���R�h)1.1\�L!���$RE��UJK�PF��P^N.;51v��0�k��O�NgoG:�Wj�0¢��)԰\,U���c�§bU�L�\ѽ^������C�	��Z�b�����4���A5!y�Amfj<�A��:��g
y=U<bj[TX%��x.�z��H�㈠.����0��i9_t3r�sOj�K%n���'̶k�9r�ȉ�T{�!Q��B��L����bG[gP	�{��l&791=0������K�jo����j��Ӌu̦�셛p�ڿ�Л�v�}�����������/>���ׯ����8�n�l����K�;~r`�R�L�iwɲ���1�l:���V����%<���^;r� "��S�`��ҝ��뮻뮻fFg^y���Ɏ*K!�Tʲr�@��i.�V)�!8�>a49:�u,LL��:��V�X+����'Ϟ���������e�/���u�+ ѠG
��C��G���������ɦ�����e���AAu�0Ɇ�bY�ś��ǽ�S�4m��{�1ED\�P����KQU�h��[ P�Ў�IE*�T�ņ�U��3jO�(_'N�{)fnO�׍7�-�O��(C����'/h�s�-�`b�p��Oy�0$B61`S���l�y���X衆�n�,>mq94l44]�Z�ĕ�2U�{3P�D?������i�I�u+�X*N��o�%6B�������ccc�sɒ%Rr]a�Xڻ���c�RW-s��86Ko��a�-^��/�+���z�y�mCJ�cr=}_�����"�_-j�C��l�F�v�ڻw�w��_��������z�8?>>��?���7�p�?\S	���ay��x�AI�9v���j:�JY0�Hd�f�dV��7�Y��c�T:�I�5��4��&���j���YlXS���ua���dfI#�����G�&�)�wz�	Ս˂zJ�;���%j��҇y�!r3MWB��9���0$�Wj_�?����)�g�-�j��m��F&���\�+��g�|��k!km5Z���	��O�{�s|�no�s���k�U����:���"�E����/�5��X玵M�u���h�e�3��U���C~,>l�5$�.�~��8�g�i^Yq<�Pɔ��x|�ڵ�R*$��Ca�ֹ�[ۑUoű���?��n��t�$�+���\�����_��K](xT������Kl��O!/�6��9Ɖ��d*#b�<y�9����RW�˖-���S/J��ꆛo��꫁.�[XJ�Vjvz���ûx�<�wU�ٳg{�	�ܹ���)���F�:�+���{�J�7�়��d��н(̼Ez�zc����Sʍ�j��G}���^�۾};t��V
@���c�vظq����$�3��w�yg:���8�����+Z)JY;$��[�+'3�B̖��P�Z�=���JYY9�~�#Z`Wp^`�$��8Cs���WC��?U��+=�a�^[�ه��ys�kե4"�.�Պ�����M��Ny .5@�>3�S2��0���t�W_T\��Њ)Q!U�En7�(�������oo��� k��@4�qI��w��K�2p&>�X�bh��mm0�(�?V�^�+���|�����5R~�R����?gg禦f��<u�į��;::^x����ͯ���t� ����L&599>66���`���I<oQB{�NYZS�@��|L("�
×�exϔ[D(O�QZ�G;j�(��Ƭ�&��5򓼗O5?�|��EM��t���'Ӗ�+�:T{��+k8R.��f�G����"�ЪMZNK��K�F~ȟ�x�D[�=LQ�}Ϥ��H{�S$���jY�8'�:#�R��5&=(�&�g��Z5/�+B�>���'�t���bP�c�u����ڑp[$)��"�(�و�7F�l���g��� #+|֞FeI	{���3r�C�X�]L&̈́-�/vX�^�����B]WS����mS��z��Ȳ6�Q�P�O�~;����	���lI�oܴ��4�oބ��M�q�JTbE��X���$��|�\���:!�zɀz��dFlQ����q�ChUTѣŪE
,���,��gUPR��!��7���tU*%H�d:�S�B��ŋh�/��PL=N�kԙ _��9��c�,������X�g����󩧞ڸ~�؉c� u�G��ޖ-[�/_~���z*OM8�q� Jh�d�ʑ����eg��ࡘ�u,\8w~fj�r�.qX�|��t�l蹪�D��uD|�'BcZ֮_�y�极��_��?����_�;��{�޻��_�:0���F;֖۴i�-7݌w����rY�b��?��#n(��`I�q�1�|dJ�ڕ�|�ϸ,��gMZq���̢�v�����1"�'Mw���g�e]�;D���9ߨ��@k�-���cN��i=Z����dQ����"�o#e{b��[��T�uf�9�9Ggf)�a�����ub��(�56==�&���4!��ɤ�O���TUW��� O(��տ��o�_���;�X{�5k֬k����x�����Z�tn�gIX���ʈK�P�(�g�<����]X�d�Ν;q�
?�gH�n�a׮]ǎO���"�{�z�����&L�FT�ơ�&^�zM޼r%���#ri��4ss�	�։�0u�s�J���H�8��0z�����	�=��zB���Nq��P��~#]��z��&]� =/̐6A�� l�1�4��^T6jR�M�s�j|���,���Q�Jˑ�ߘQ�	V��Z`�F���_�i�0Ƹ@���D�N������Fa��l�M2m^�h?�餭��w�4]��1-i��7���f�@��G�w�[�t��taq��N�,䖦"��������-�����Gqr #i���6n$���8Wq�/�XǜyFn�A�a�$�l�(kV�JEzWD)zzz��'���v3��S�NAPP��	I�� ݄+y�T2-��5���N��ln�O��"6���^z��W_���>+�B488�q�)դ䑋CNq�XWOoP.?��#������H<g��=�q+%ݖ�&<�@"�6)#*�o ��=k���>��ٲy�֭#�{�ܹ�G}�w�x��w:t�ڷoǟP�;o_�>�s��-ܾ}��ӧ1W5N&�A���,������V��ňj�g.h"6�Tu��t�%�fڎo�<���VM+��o:��5ц�J��;?��h������F�[`Ʒp�Ա2�͡擡��oCD��R��*���w���Qn{`K/���V&���l�x�ZP��$��wT����*�D�8��QVz��/���S�U�5;���K��ڹ�����%����)fz�w�<G�S%~E�_�Ղrqn����cn��^I/>�܏�a�� ���Tq\���D.���Y�
O�˚�k0�����J[O��kxx�ȑ#�|g��e��J�ɩ�M��8o������v��Ê���,B�
���r�T��fQ�&�(1�J,Z��1;M�u�A�$K�4���}@�Ȃ�i\�p�����;�]P��[��
�Fjr6�/�\?�j{�l����a�cޭ���j�9�e��Pfdm4�;5�v�Z7-��|f�&�,d�a��Sw���jQ��=�Xj���P�R)���A�fB�I
���F�%�x�q&�V6:�,�*�������/&Uc~E�Q�c`s���?�}�VBO�t�R�Ľ�]Wu6|��s�jf4Em�%˒%��l�M܍mB�GH�!���<!!_����		�yR(IHq�p��"���zo�2������w�uξ���2`8�3�s�}�^{�w��ֻ�3W��pV�F�+*����M2�����;��^ ]S�_���"O08<�ܤ��|�9��)
�w9:Gn�׊_��>e"`�2�S�U�5�ι�js�=�6G^��D* �8�x�;}�tSS�ʕ+�/�ŭ���Uuèl������T|Ba�?+�v*:?��\�G�����'�767����X_�Y��f��!��Q���O��8ght-iH�Ci,^���{�2��,��166���b�0ZXZ��E����#E>�N��ك;g��L�,ŚЦ��:�͐t2Kw���0�1�0���8�Gg�'ZBdf��EJ���)��a�L#aZz���dY��5��C�"�ZvI�.Z�����op �_��irr��g�����o��&��x��O?�a�L2��#��Ώ���T?���j\2��
�2��R>a�l�������X���0���A�p�
���F�x�ē�E����0RN��?�j�j�`f���jN���/�Eo��}�ey=2[qȜt�0�*Ǧ:��Tj��z�6�S��G6�(&O��I������i*�dv��_�饖(� ��:�:q���XKY2+,�2����hj��\��mɀ����H̏%<n���%��AK%�X̫%����@��&�922�st��c��۞�b&��֯_��w��پ};�k:M�p��	�12�Q�/���A5.�����`�V(>�����s�H9_|�B�����ĸb.~j!Xɕs�,��f�r�)1�6�z��T�J�Cb�K�a�e5Ɔ:�<O~��)nޠ�"���V��b5���ØE񶊕�L$$ex�r�`�<Z�_��iE;$@	��E&�z���`����h�����(?�֡R��b����\�#�򚱨������1�#��C�9烴Yy�Q�]�����UFsȩ-�g�'̤��\��<}5�.�r&q�
dw�D����,"��^�.���d��ޣ3K�P�tg�S.�j����-�����@��"<�����k��7?�񏅙L�={��5k \�2?#���Vkc�Ϟ<z�a�|����2���'�������^<���^����^E�������33������-[�xL-{�x�lȸG'��2�y���|�����+�*nQq1�!3NV)' ���cy�24
�}xxhh��K/]�n�{��������Z[[q	����N\�j�*���/>q���� ��N�	�o������<K�jjT��|_s��愪'��Z����}�P{�\�ǯޑ;�9J��K�b痞Rw�*�AO�����<�_�������ċ�)� �
\�)��+�Ð|Ϛ�
ߛuپ�Ϛ��c&MK7��ck�hdﬦ�~T�k�9 `���X8~��ݝ�I[J%�-����ڿw�],�&jS���=F����ũ�I2E�<�<y�wǎ7D�P�Q��L�g!��L�0�9ݓ�*��-����0����,�m@f�⫏����Q(S�߮�LMM�߿���/�m��%�NGҤT,!\��u�)�|#.����R�n%�4�9�`�l�t/�/�h�t�vBS�t��r�����=�v<���3��t:�n��z��ϕ�i3S�S��X\sl54!�U���FF�f4k�(�C��y~|P#	QcD>����gb�:6CR#���-:MX����)�H��e��R/��0�ߏXo��hs����/4��&���U�pr1�"��]��Bc�!�I�[���YZRE����>��M���
a���{ʁ�Xe~�*o+Ud@�C���?�=��Wܰ�)���Gy���J�[$\��NFO�1x�@�����Wb��#�#G�aV�l1R��'�=��s^�-�5��!����T���YV=�3$�l ��I��Ht,P�[ڈwiC-##��q{�I&t��\j!�|f�Tmz�Α�;�'b.?ӳt�1�	��BK�X,�LN���Y@���I���
~��܂x�4-2*���n�f�W���^��p�S&�E]�a�F���N���������|�]]V<a�X	bɄ��n!`�ރ��55�OM��y)�S*���|.�\T^�ǐ��ؐ�3W9�"!���K2���C0���QÝD��I<���a��0��x�K.����/�M~�����_��|��W�<y�ʶ-�}�߸��{?���N���]�n�}�{���߿w�^,7˖-lD{>�=�9<�#֜x��>Q�i�U1�_���n��p�x�٧[������"Y��̍p�T�jUǅâs��@���7��֛���z�~t�?+/sd6��P7��;\WhZ��Z����_���i^e)ՙ���s�'���1ô�*�=-��R��r�&&��j߾}��~;�| ��������$��F��(o��a�����C�w��*��y�D'-��0t|;��Z<OR D���i���m�L��7���1��a�r4[���[��r:x�`C��YQ,�nmٕ����3��p]!��8�d��2��������}������{����l|��,{~0R�+NFWtw�Ϥ-���l'�܇�9��P��1�K8�tNU����9�0�c�E��R�Gc��_��ۚ�g;�?���q"���HY3��w�+o)���^IR�H '���T� �
S��}EK����f�r����zd��"�:�kr���j���C���1�,m.�R3��	��#��ڗm�?�'�H��4c��$���d{�!e�[=j4�6��V��Z�jn��6��H��w����ى�\\�2��53��ܼ�#�R�T�X�]!חW͵�<p<_��΀fc]gu�,�`˗/G��Ri�Ds1�ٳǏ�)e��I���p���:/H�2�����~�����C�@�K� ��3�<��݅oz�-�Wq���l��#?�я��� 4���f A��哛)Hj��	Y�Ą�1��ׄ��4_�B�o-�}(�� еk��M������_��_}�'[��{OO��M7�4x�����o~�ܸ���W���;�c�ʕh0�A�`��O�b��>���9U��
���f�*+Ww�e�Eɉr���譄|�����c�*iI
��?�m*k�5��c�̾�m���h�d��#z��{U���nq�/\�-�Y�H&�	����'.�Q�D qDI`��[,f�
.�������`ˉ�p��(�<� ���fHYk�+Q�L)	 1�Ԑ�fR &�z�$b���;�Z<|zjJx�E�h��	��1I1]<.f����k\�JИ�3��PR�JdQ���Q�T�X��� �	��R*�W�����L�������11>2i�npBE�jR�ܓ�KB�D�[�N�c�\q������2�K@X����L!�H�2T,����Z���g��8v�+����O	VMMd�Ɠ	�Eh+���&'�$����GN������?��X�X�uÂ������7^�h�*�j�rm~U�v��a.��l!���i�&Rq��|/�/�&6�W�%�'�C�Rï,�5�	"���94�f�h|����/�
�(�̴��E���e�u�Ÿx���$">)���.=�:`y�=%�q������D�p���cF%]��3@,ôB���8m!�R��,'�(�H�6�qb	����|� /;==�������Xt����Ĵ�x�<��P����	*[������Dw�T<쌔���gR�Ր�6�J���e�ΰ��:0ENq��j��Y�f�.�;e$R�hlj�d�Wz���X�7�S|��.j-��:Z2"�ԍՖw�4E�2:g��=�W-߹g'�!f�NDqNKc�@�H^@�&5�&�=� �H��X�J�B�����SF/�djSm�����be�����6	46 ���.�;-¢gP�
�<J��)\�4�wup`!X�l�o��.ۀ;��q���xbh�XB����X�b�
�688���
]$�����w{챛n��~���LF+�'��w��516�I�J$q+Fy �x&O����x�`s��*���m@+<*�20	����(�	����/�0%�Ѹ�&�m
�A�@�>z�=�yϫ���m�s6,[�z5@$��iӦ����^�|n�ӳ䮻�z�Gpնm�N�:A��O
�ă��KWw7L��q
t��;�C��D�2d=�죣��a%)^���ҫD�cF�h�ΓE���#D"�l6t��s�y^��~8�p�$�]�)�1� �y�f�5#�t��)�A����G��,�l��/`���;��U�\еj�3�%Yf!C1i
�R����<ӂ}�9�??�m�<Hw�H�gI�i%\70�����Vyɸe
��Ìv1�?1-5���ӧqS2�8�X�e�j�sE⊄t�_�� 3<�Oc�&
������Tt��Qǉ���5��c�1��}�����9����D+�������r�+U.�+�qe� 4���e�����/���p�J��:ߠ���d��S�_���;[��|�L���<�B]�JpJD�W�;���?;��N��P�jz��Bg�r�(����,;�l���|q�za����K����˓��y�U�Rŵ�\�ui���܇�{P���
$�����R�ї�N:=�!�rs��%�ȓ�Fa�uv�*�ň�&�8�r�X<Y�c���2�T�H����]�u�~��C'��R�0�"o�����C�6� _SzI�*1��<=C�D)7D���O+����!�b��-of� A��"	�����N�6���Q�52��Q��<�?/�ͣ"t� R�X�F����t��J{��j�C���Q�f�R�*OH@����.�A{e�Hj������'d���d"B1���NHث4ƈ&��W\I��w��V#Lޒ�k���D��q��ȑ#x.�
 �?;Џ��q�p�7��g˖-xq���e˖���a�Z#D����U�X��{�,-1Ć�K�Oɍ�ב'{O�(CV��O��d�_w�uh��O=)A/+W�\�hѱcǞ|�ɋ/�'�۷O�.��%l�������w�o�k�.�0(X 8\��FҎ��(}��Q������ľ}�≸�>�92���.�%>s���s�Ω]+��ӹp��t��!���熓�\"�~9��ؾAM�f�\7�����f@�$����dRN1���*��b'�V�S�-�0��c�����sJŨY�����m�5�1IB�a�skW���֚�����S�N����V�Ψ�u��	9����i����V/�.��j��I�&������"=�G0��*L Z��{�' (1�/^Xv)�[��R���bH�iA�{grOϵ9���M> 'q3���oē�B�|��i�l�4��/�vm�5!=L	�|�u]]!�1�Mi��u*M��
�"^ƶo�AE?�H��,����JL�.`���5���<�C�"�Th��lO�a��*z��{ʳ��b��(�4q�I..K��	���L̢"�%����".��z>FUOi�\�Q?�z;�J&	�Z(.�	k]�lu� 31���13�jf8#f9v�)L�>=��iZ�p�{�]3�D�t�AY�1˴|��~k
)�uyM�Tf@P��0�V!��tK<az���;j�9a+�`��c�8̌
5a4�b2u�qRI��-3(Z�h��}i�B�?�@!wT=�9S
g]]�>��$���:�O��h�/�:܏H`�ƇRv^�K��KJ���2�A�%��+�#�ĸ$�ȕA��ɭE��ȴ��eW��j\����#G#����w�0344��K�w�,ɟg!�\�2-�ؤN�i��yK���c�m����}hdlrrz�N���nZ�?U֊!y��f54d�.��/P?s����u��T&-�)@`��{�b�m�pI�P�MS�
�3<2�q�0��A��Hb
@�Q:BX��K�5b�-��) ���6<�06
���m"!���[#C����d<>00 �o���cc��-ӧϜ��Z Q�.�����n�z��pg��f͚g�y�_s�Z�����=5�������z�m۶����kk�xuM�MI�` >�{��	 �Sgq�d]�����0@���z�Dn��SK�I�S׆��k�"�Ԕ/�B"�=U!��/&E ��3¢T~�y���LHVu�=^��5 �fuQz_]�4������
�H��6Kg��;s��-����L�a�_B}���~������\~Z�}�ww����eX!m�M�rL�ё�!?��M}��=C�`�I�´�>�U؇ !�Ĵ;')R��Y�>���C�������p�k���t��a�edj)����W]-[zC����	ʢ������¯�g���=9n�����ˠ�N֤�0�1">;�pM�]�fX�Q���$�g����9�]s��9�����+{U�`�Di�xU�*idC%���OB�y3��/jP�H�D�x������>�s*�!���Q"^I���4� ɰQ�!fH����Gr�dÉp� c�1�J|��O�^|ɉdZҴq>�Gy�5-���~`�u2
b��i����3=��|frϨ���
+��9���o29��7Я�C�
�5���	X �`��)3S ��d�HW^Y�ʝ+��s�v?��ʰ�ҍ�&�lT,��}tލ
ǔ�-̼`��7�yʅt��+,bb�Ȉ>c# w.�ʒ��FFX�T��q فU �a����ǯ��J ����
�+$ޤ%x.�GSjSQ��رc��w����}��8p476��3566V�uy�Ze��r��&�#��(x5<��(j�ΝK�,��� �
'�[�k�F0�BW!Q��Z���ٚ�---��?���K��x[��5iI~fF�mP��[.z��8���]r�%��N�.��R �����7�x�׾�U�k�������x�7da�[�vٟ���/_���[o��u���� 0��mR�s������9[׈{�M
%��V�D��W�xj����#�_�6ã��QT������$J߂N'�$+��)t;����?��K�m��pj��9{擞�����
I�KD?-��f���qr z������R��0������nQ�D]S�b
�Ԭ�le-��g��B�E�2vi�ⅹ��cǎ����5j:wO%��<�p��@���i\f�8AJN)K��r:�����v�t_*�����v�l�J����0#��d+d4ź���ljlX�r��������o{Sz�O���A)���R����D)��(�m��V��f��UqӍt�̶gʎ��2o�@����2�T,�a���[߽]�y��c��x�0��nT�,�w�T8�<�M6tfsB�
��C��Vt�8�LO[)¹=�q����֭�ar��Wdr�YM=�b&�Ϛ�X�N6ٶ�@�m������l�a�\$h¤h���S�('()�UX�5_�"��]��#t`��]Y�d)Bfȓ$�Dȴ��RI�v!�wmc�)1Đ���v�ŲC�<a�UvʮME�L	@7�{�J�R�)�	P'd�Ӽ	^K��&�b|���)ǅ�Y�/�kAv�D_��*D"�3.q�鬄9�&�W�r�z��x#��BG�)�P��� h�j��F���(^���1{F(�B�vU6FX�XתBf<? @�@���6\]�0J�����9r���K��h��%7$�9��� =�Ӌ�e��!0d����3����xc}CSC���[�MJ�%4�&MNO��<
.yWI��Fdhd�������ݝ] ��������A�B�t�Yڱ5̙�t	f�cclD���-%���X���{Asc��!twv��#ƥ�֖ŋ�����m�4V�v 8�rz��@Hcc%�5C5m|r�s>U��h3z�p�F3kdr�m�Ekѷ{��������?����Z���������'ONL������q�ҥK�^}��y���X�>{��Wa��\Н��\ŃG���u��6mį�V���G>�s��'N�M��PV������.Y�!z�E�����)�+�T7[s��<$�ܛ�ѵ5@�Gb��[�am͊`�<_�̜Z}�{&?��A�� Z�c;�_	V�'��f{X�9ԗj�����|
�n'����T�h=�Es7��|�c�|���za�MTgE��3���ov���V��;��C����t�`K(�A~5}"J9��[��<69��dWe2)��K@Q�lӈ�I����)ѭU�u(���6�P��[n�e�ʕ�����˿�˗_}������WRid�MRZ�)|U�;T>�΁GȰ�)F_�}cE�$%J}����!:��5��1�v7c�c����/"C��9jW�Me�JDB��sG�屘-5O�
��F��-��%�x�<?�א
*�s����)ֶ�S�sH�X���M���.�S.�Y%�\ 2��V�IH=��2W�R芸�9~?؇5c�E
r�N:���d-��(�B=XFT�|�F޾����-<^D�U�{�U�}c�x2�P��K�R9�*�B�+?,W�3ۻ�I�$bq��Q쫇�t�'��ⴃ�J�as0�Pe��H�'9۱=Y�	[p�3IЙ����ٙHQ�� ���*j*����_��)Z��@����BE�<��3���w��%Q���l��izR2]0^��K�}À5��淶���w��Ԃ-⡔O�t��GB�*{/Jk�� q�H 1��e+.v<U�>�d�D�=E��l���'���9���+N�����g>s���Gy�&��q�2�<Hód�ޫ��"O)N_��"3�	��e�]v��)���>�KS�����jhX�dɊU�������D����¤He2 X ��=�ؾ}'�iH���^�`��Ĭ�H)^���:~RMw� 
�M���.�x���Ӄ��{�>� >K��}����i�&�:gŊ[�lA�ѓ/��r.��y��$����/�d��Mo���U+{�����߇@l_�ݞcd'��3l��[��Q�ω�pgL�����"�Q $�^���Jv�\\�o��V�hV/a�k�'U"o<�����W�D���C"�?v�T�q5LS�� (��������X� a�תؤ�{i�����Xf;,��u�����ڨ�"�/ig�:=I�L01�-[�i���O�t(Cދ��c�5)��]�ⓓ~0�����XC���ݧ[�իWc��V###�Dރ��y�k�.���>(��Y��&���j��?��d6��˗�R��3g��n���4y��Ze�*ŧʭ�P@�>�d=|��ԐNSڐ+�+�Yܗe�,Ey�{%ⴧ,��ušP�&e�����	�B���X*�������L�U�*�^���Z��X�f�t��\ǜ��l�(1gbO�R����z����$d�+s��W	e�
��.h�hmi^�p���V��"��r�
Z�`;C$
�4e�����*	�jϔ�J���f�Me^0�BA�^O��r�+G	�L��2M�$Ӭ�4��c�.�hɥm�X�qgy_\!oll����E�kR�
Z��(3r�s��J���\f�7G�Y�2�#�1�}!��*gB~�������~(	t
��L�^�c~'�bhdHұ9c�Wr%م�,��I���$K�_�W�����a݌
�^mE+u�+Zӫ�Ry�uQ��T:M\��g��t�W���k���"m�-������JDт�rժr�'�ڛ�!j�C9�4�v�w�{;v��&��4.�2?�����T&m��F4���G�������w���+0^1K��5�j\"}���� ���t���N�H��B\�Q�Z:g��tht�U��#���*S�:\���v�Eaޑ�<�2�����e�>{���ͮ;p+�#�K%�&Ʃ5N�B�s��.]�`A׏� �;r����_��Ͼ�a�)�W�Z��Ï�2ݵg7f����Y�K�w�,[J!����wva��x����ffvuo޼yɢ�/}�K��hL�D{���Uru�cSE��dϨ��R�>Xv��,�e�m�D\E2�Z��l��h��C	pԋp���`��D�>�V��Wr�^�1��*���+=���"ku��[�c�{ם��S���h�y�#�1��F�,!�W��D�UJ��\��}���k�^{�O=�#�����E�q�xY�t�bA�ǫ7R�+tRY^�Z�i^~�e��f�>�o����h̐�G�G�!�-�!��5v�z�h����1�ک�ǂ��K�o��}�0���Y;�r+(b�㤅�U�@'���%��W'�VB��8^>	9i��N��|����GG��d����h���P��\��Fί\^#�s^����*+_K� �@�`��3�0�%SO�p�.�;PnB>	�����*;AA�J��u/d�8^��}�P���(������ -���������T@�e�$�T�:��p�c���0i ɜኊP�����ɰrPz���\�hnn��.љD �6:�5Ke)h�rֹ�)Kд�d��2{D2�,�aEW�
�F�X`�|�9CXO�	����<�V��͊���ȋR�G|!�TB�����P�<ˌ��V��f
��p�l#�]�����;��\�_���Wn�ja�D,�F!�C��5l.!��4�fL	ym���vԈw-���g�_ko���Vd�IBa-�=~��%7�<y2�i�����gd,Ay�`_B���G+�&S��?8�$�r-}�7^q�[�n�q�����,�S�r8���ě_(~�_��[h��L�8,%�ʰjh���/�\|/��H��L6���S$t,���]]]0��*�T)�����@U �$�l߾}Ǐ�*-Z���������ܹ��ѣ7�tSk{�]w�}�],
�����������
�R
��� ��1�-���N����v|s���6NF?�яn۶�����`��|�͸��Çq��?�A(���)�]�~�z|���pP/e�cv�ˡ�+�l�6���Ŝ�]Ӣ>�d�h樘UUV��$L�#,&+�)A�?5��}(c�)f֛~�.xI3����e�q��'�N�A����h��������������j.��0�P%��P^=��KQ&�ۛ�x{wLA$Bj��6�V�r洏�q=��2oS45ԧq,O��C�x�$z�3�� ���yG����[��1�4�v����m���Ð���	 }�%J�9� -�"�tq��I�r��	��X���إ�7�����.s���Dym2���H�Kv��O�$"�@h��_���9�nbr�J%�]�Y���[n��ګ ���N�΀y�9��֌����ӳb������$L�Sb9�~NMM����8G�Y���.E�brRp�����.Y�Vs�lC�]v�������wܡ�9)ɡ.�$�����tʱ5�JNqr-�q���r��gQԶcp�4�z�7�jĢ�i�l^�L8�dE`�#��o��Q���$3�Jk�唩���$Ƃ�Isdt ��.���,|���EF�ơd2�a^%�F�D���!��TۼD���V�W��^O��z�t��`Gr�����+��qN$K���'�h�H�bxp��4� �����n��e2O/C�YZ���L7I�_�e
���\ 
�A+9���(e��s�Y�^�-ęb�RL}��� �`\,��D�'�|�\�\r<G�*$�JX�rْ	D�7R,y:7uv��)aC��IQvr�Q�����̺B+��Cj�z�
,J�{�ɉ�'!{*�8V���!4?<�.~h�	�M.G3�x��Ș�oNLL�]�*��a�(��OO��`�ļ:oPJ<%�"Ҋ��[�aK�<��$�T���Q�*8A�ˌ9$��"0�'yd�V�Z,��ӆ��%7���gyZ�u�%��A��诘Pf L���4���2�ʣ��PP/xU-�$�=|��f�Q��$�/�&�%ߋ&A��,S7��d]}���X��E ۶m]�xQCC���PE�tm����Kft�I^*�9&�(�
o��T��/�>WO��<O4�Q�xy�7�c.����xn禎}�g����{�sA��Aڈ@�SD�g9Ű`(E�G�1
2#3����u��W^G�ꛒ���S2��0�b���hOKK�u���MO�~���|��ĭX"7(�Ӧ2�x����&�q�?�Κ����\>3��<�7(v榍W2-H��w�e�{{O}��/������|��0��0/���������#�<��#�oO�8��X��kz����+�57��c{����w�3�VǵW\�u(��'&�?���_���,Â�����w>��Ǐۼy3:�v�k;�x�ч�{�u��D�\�R�;ڻ�,�ܱ�xC&ݵpy>G;�\��\� �r47�t�"n�,��DԦ����}K0���u��f�㖓�d�T���Ud�Ry�%��`1��<�wUUM�`��z�Q��(���LQ��p�
t���+ej��F�2甖��n�L�\��4��Ci��ӓ���[9j���V�͞�z��T�'u�zY�8|�&UJ=��K�tY�{�����2yn�T�KS�Q�+=�a
��=�p�))�����$?����}g���?��Ck?��CG����L�6�x�)q+�V>e���b(V,h"́�y�7�p����oA�OO�=����_zb]]#��^�dzzF�u7����x��wCy�ݻ�D�1��lT!,6F��4ٯ�0���ž\K����^��9�驧�~��Gm��G3�P�k*�<Z�Ai;-���ÎŨ��CϽ�������C�O�y
T�-���;�_,:R,/(��<"?$��&��̀�� �ߔ�It�,텂-!�8qd��� 3�s�L�āT,��}�c���Ѐ��'�D�i2'V�P��SORq]��d#+�H>���-\�O�����]�/��	����	)2&M�����)��*Ҥd2�{�E <�G�inO1��$;�qdKM*�r���E�TmB�zL57䈱=q�T`���I�K���|0ZH�f�)�Ky�G�}tL��5�cٲe@�p�����+�n>�\W�Oӥ�c$���%c��5hͣ�����2W4��A5[ɘ��:��_0� 9zB"�^L����D���E��E@BR_؍ЛUz�#<�#jVoV���g�c�u^x����`�>��3�C�c1���ǭ6l� ��y�2�$r͚5��~�?t/�7o^��#��LYY]�����ʗo���~����8q����iT��JqɆ�Zt���к�TzϞ=�[o�u��������]��v���������_|��+V�ڵK��W^y����e���.{�=���{�o��� ���}xժ��_~9 �k��?xd۶m==%����֢����D�����@@�Ѥ���z���ǏG�6�m��O���/�ᇪooo��;v�X��|�V��d���ԴL5L
Q�c���p�Z���0zfTH�q~���?����M�!��a�R�C���t��z%�{��AD��U|�F�GF?D_��m��ƹ::z�ܖ9�|q�����p�o���K�R���4�?+&C��9�0���M4r�Q8�x7S���(H�ur�`���a��&���Д��>����{{�-:;pz��N�ٲ�HG!`&֤�A�dx*��]�P�t*��Xc���>��{�2=�k�+?�o�Lƣ��GG�	*�b�ʓǏo�l��o¼~��ݻ��o�
H��S���M��?�����ka�ٳg2ٴ�ꜸA�6-�P���O\}�5�2V����/|�_<~�d��k�ۑ��㦅N�Z�86�%N ��] �~���kE�:v�U�c�:ʾӼ�сJ$��DF��5�$p��2��7��2#�R���JxU���d�����m���������"��H��6p���d��K�����������q�1�0��g��WrJ^X�h��1ס�.G����W^{�w����4���){.P���\( s���i0~b��H$�6�8Sqc�k���v���F.Lf�v|�T�)�K���|�����q@��P bSC�ϑsB( jkk�ǡ��ȱb)��[#��M�j��%<��8q���/%���	.�<p�����S��5=3k~��7n���[�n�c�z�{D�.��w\��I���%���ܼ�<��RSu�jZ̟�[���bN<,�I-�5���A������d����W�Zb�opC>�c��eK�N�>S.9���!�IUa�r�Г�#��S�El�ò$��OV!�b)�1K��mgN�~c���[�{����qq{������PJ3��tA���7H&�	�}�M7�n?��C�[�<��$gU�0;r��׭����s������-��
�1�D!������E�Tb�d�P���{akk��%K��?ѷo���o��o�t�~�a4V��G�8$H� ��u�.���d]�W],�g��?������������~+�n������޳+V-�﾿8x�pޑ��1�� �aӦM�[gϞ}�;�h��~�[߂�ؼy3tΫ��*!nbL
'"N�|饗(�4Q724<9:�b�
��&�O�z*S������;�� ��Y6�3	��[/�6'xx���5���n���5�E�pސo0Qd���J&Z-X��H.w��/�?J}_㯊~�ȳo�U�*-��N�KV��ݑz�\XЏx�� a�HF�d��ө���b�,u��E��~�z����� �&�000��\��	�`n|�{�����W��<(��NӲg���äۖ��ĵ%�����������b��_��޽{w���9et`�9t萡�[[[1�_{�5럌;��7~��m������?�������׻:,X I��&�û�$��˾�>�w�qG:�Mp������;ve2I)Z �*��1S%�O8��y
���KK��̫C�-�H�/"�%JKC�TA��4=z��/�ye�V�!^���|5!��!m&ls-ݢ���K=����F��X�)�����1�@�ʧ]!.�'>$�@�H�s꥘�AQ���p� ���~����/�������rH�T����<8�˵����ķT�8*�\�u��x��Ip4E%s�y��z�&�*eO?_��b.kHc:44$abL��166&=S�k�8�}][��M���g��O�JxD�d�fbq��i�v"�*�B�z�%f�t��A��:�<I�����%x�Bf%�_���V ����xo%:Tۘ������2I���ο�ě��1$���-�C���e��6�}cX��n�lH2�Tz����#^F3�䣇.F=���o=∊�t֫�9"TѮc-�C)mٲh�ꫯ�n���6��A���j�vuu�S �N����+W��a�m����ܘ�� ���K���4ХбR].=)��ZX7����P�TS��
����'��Կ��� [���|������T<��g>��߷���U�V}�CZ�|9$v��=����� +��p&$�ӟ�4$������O�����M7 ���-����~����0�m�B��F���ի�o�.�q8yllB�GK����B[T���o]��B�����׋JU%-��g������*L�G�"��!
*�Y��%�5Ȭ�i@����1:<)BIk�!�3_�$&��j��J;jZ�m�9����Ij�h�zJ���$졢4�FE�U�N��8!�-g����%�D�߂���K��Ǉ���=mmk:�h��1#�+��o�,=�5��&��K�0b}�5��iDn�a���]*o�t�����`uuu���\!�8�L����A���+�TA��M.�-�V0�0s�/����}��/�C [?���\�-�Lb!��Φ�X�5�jkm���\a摇��&���k�����?xݵ������>;6>:9�V��=;���	�	�vR�`GG�?��]�<-�_�ۿ��s��g2��2?eW�b�t/�S�!o1�"�e1S�?�IXK�"֟�F��|�'buݐ�1L��/Һh����`#��I��A�����㎫%b`�(�W>��1'�=W=�Bg����#���4���<�,�@X浵�Վ1�5K&��t>g�������F��L��F�^�*��C9�R��+�K\�"n�UI����d^s�5�(, �E^���C\G���'`�ƍ!X���),=E�ˆ"�3���L���� {������dqj>��AC*Y2�cjf2���)�g����͘oxt��7C�K�R'));���8���e�=�2�����hXy|T`%��RIX���ը�*�&)!��9���Դ#�x�L߉S�� [Z��Ÿ��3e�Cs[�ғ:�#��~%?"��I�1C��@yB?sx0��zE&�H�M�k�9C1��V� y�H��/?��,��c@&;�h ���{a%����%	�=2J1��2��+���8:ӐB����!�13�k�T�=M��꼞��S�ݲm�4�s&<rQ�K1;+;��9�'i+��2Yt[f� �H�(�آ��	&�k��χ~���.��'>
�t������1�2�9x�X�¶�{��I��M���bɌ��ш�.p��˒bq�'�������~�رB����P��ʖg����1;Jv�ȱ�Pڀ\0v��y�%��\���#��o��V��K��
��x�e�{zpf_�U�\����U�������×��h<t$O�[ttt<��3�=��̲5k� &jU9�|���rVd�~��e[����~2��a�%+����VRRE-R�D�dS)�ep�a�1�~�U*4�W���7�e�T_sSGg�� F�RC�ͅϴ
b�BS�4ɟ ;Z�����;ף+���f�)�o�X�*�\u���z�Y������fԦ���
Mw�n���!�v��N�T�v�������>E�l���@��ᯘfX�8����l&�ЇȢ|#(#C�aE�����|�#X>�&N���$��kb�$��bY�=<�׉�_Xדi2�q�;^��"�Y�h���_�v�Z��g�y
7D3N�<Iiϥ�<v�o��E�����_r	E�{ƃ>x�}�56��-�_ú�XIE;c��
 8sZZZ�볌 �%܇9S	@��UɮDakad�+�D�W���U�[<��N�t�IXM��uKy)���[�xO�_�O��׊��[AT��I��T&���� aٛ�M�� �	
�2"�6�:�/ʖ��T�l���!��Q(I�u/X�x�-[ Q�֭ۼy3@���x���ͻv�ڷo�=V������Wؑ�����d2�<v��P=Z�F*u�� �z$�P�;qD�����`8ۏ��^�!RI�=#�V*e����c&�86�ǨR"WFR���O	�L�zUl ��!�R��pO,���&&�?|O��E�
��Q������ޚ�da/�ߴL����`\{�NU��M�!>���?����+ɀ��"u)(�-��B�yE-�I
 �Fp��ԴU1*FHbGM�7"*W������R�Y�\`
�4ϛ'�>:::61	@�Ɛ��ʎ��W!.�B��� �U�d�ٳga-Y���nC���/^�h��]qHc�=|��l\���p�:n�����b�(}(���Ɔ�5�4�@B�,�W�9��crzj��բа�۷>|���o���~㍝/��������8�����ֶ���>�ׯo�7����o�����˿���.��~<��'�ǋ�{��}�=�P�/Ͻ��@o����ɜ I���o:1:F����NM��5d�%���S����zd�m��+�S�_���&
 �%�o��L=ԟ��Im.� wn<O�q����(��Lx���r��X�.j-l��T�f��1E˜+��X?�����M
n2�4����F����1�¾�h�XR�sV��{��w���<X⤝��L:	�Iuvٝ��{T���{�]NlR�D<������w��K/�M,fۂ��]�eۅ�(��b21w�R"]�a����E-�gX���]P<𽧟~��l�>�Y܌7f;;�\n:�LIŷ�m��2�=1���w�b�`����!S��<���ϯXхk��bq�����r��W]s-:�vܣG��?�c�X�&���&�3Y��eK���-�{D��Nb~��G,����:����&��S��1�UP��ϒ%�׃b��[V,O�ߤl�FB^�3��t1�ԫ�{n�y賶��_��y;��9��5_UL�@=�Z�����%�B��D��e꩔j�J)K>��d��@{��d�b�
5T�X�ՙ̂�m�]r2�ݽ�ʪ+(/�\~v�!θ��ۖ.Y��K/�n��h��4�S���W�1������Mю���P��@��[���%�i&�ŀq�l�.�1��vL3�ҋ�ohj��H�ⲄK���Pٗt� ��`y��"g��\�d&EY1��.���D���2�	�	J0b�%��]YGMO�ZF�T*�JcJ���C���f0���S"�,
V �"3��$Zh�)1�&��bnX��tJ�)Q�%�x��Э�)Ll�,�ر'w�,M;�X�s�l,Ű���Z�*�Y�;m�ӎ'kgױ��2D��#���e�LC�|=��Y��.'T׾�C��&�4:D<h��i�����J9��<e.�
Y��m�6ϝ7��C~ʥ"��u��0��:42��c��S�����<��sK�-��0#�	��O��v���b��k�.d�3�,v�0�0�����M��7��3���J?�c�Oo�I{{;L�+V�޻�Ϥ��V���Y	X�Ų�s�ޥ�Wb�^q�U�量Ҷ�ɓ������w�ٻ������@��o~r��/��R�dcu�'�?}���I��뮿��瞻�;>�>��[�n�%���h���+��F��JΦ'&�'�qb}b
����X�ʅb�yc�#PD��I%xY�=?̣���U��辟|`���~D,g9�j0\%��B=���_"�����A˪�����M�P�3�ٍ%���OԹU�]:��Y�j�^xDV6�rc��Uc�(�׈d��֬�Q����#���*ڧ����Y�WZ� y��a>9�ݐ�Jc�=��4��Kp��,�;w�<s���U��o�Z�a{�?�裏��Ʈ�暑�abW�����榹!����6�:��^z饃��۷�!��"�d&Eۗ�#�ס̲��I�V�x�W,X��H�֬YSߐ]�f�����.ٸ~xx78C#1	�.{��߰a�'?��믿��[ؔ��7���;vH"�HQG�&9�v� �]��B�%�q0���h�*�"D�,ܯ�����i�L��7���F$�(>�ɩ|KcZ\5h@�|��7Ai5�{T�Y���(�QLF�%�e��'N�%Q�g��o�t����ն]�:��3О�l:#��������=/�	q�a�p2z-��Xu`�D"ԝ�tF�����	v����LԤ�\���-i�S�3"�L�f�o�*۴��>$��$^�g/i���L�%�'�g��~�ҳ����J��8rT�9��i�@%���;*ף�S2 ���q�S\�P\e�y*�[�T�K��WC�e�aͨ��GMj�VR �!-�%6����x����qª�گ�P��geH*�?$,	���֘�@C!uЄ�W�3ŝ��;�!�n�ui��X�cZvX�W�5jZ$O��E�K�;!��g�-���Q*��y���Do���򮮮S�N)�.��������ǟ�t����S��/�]"Ô�k��8Ɖ�qa�rT��咼z�����|�;q<��ȋ/oG��?����իWSBI�ٵk�inn�9$�b�}�Y����l��Nkּ��K������������'�ׯ�xݺ?��?��W��{�������o}��ȿ�˿�۽�����f�K�.@{b�i�)��h[GG�����C!���2S�q�E��M�,&r,&��%�zu����u�,*�$��#���/���8���bQK!��\�lQ@�/6:9T%v����C�ʒ�dy�2#q]Q�Rӏ�����I�W�L9�;�DwF�?�L�5ާ8$۰+��L5"9�B�U��+�X�,C�t��(Ra�xD%<1��aD�{AH�ϨAb�E,]	`�l&�4�OLOQ�_�|�A��Υ	����������a���?����ﺽ�m������������Ǐg���T<����e���q`?,D���%�6mJg2�v�-hfZ����~�Ⴧ�c��P:�#d�`v���\��]]{�;�����g�tww�q̓��05_xe; #4�;���/}�/��������t��7�����Ɩw��]@z�?���o|�|H�b��c0Km��cM�?�o���#tr�"F�D�h�2�Lϐ��z<�/@�Et8�?p��@�!,�L���S�}]���ڔ��������	pр�EL�p����"�a�pp��$vB��'�-�G5���lj��޹��B����;;��`f��D2��aY�pԡ��IY��?:)�2I���ʭ"��tf�ӝb	�G��P,�A0\��/��-�₲eb򴮎.��&���\����F*�ohj�64l����]?9�GF� 	������m���K�*�ƭ�����a�z�a�nnhĻ�
��lCb^j=�L564b0pN2K46	]���4��XV��'�0� j�R�(z|���t2�H����0�a'�����W|�-نEEZ�	����l]��%	tt&�Kr�R�/-W$�S��u���.�d;n�)�Pr�vo¢g&��,^V�&`>
�~N��h0���8���)�L�eB����B@7�s�.A��M�8?31+F��zɱF%�C�?ڬn�o�Wރ��*p7�9S��dj�;�z�la۶�a��P66�OMMĘ��LU��Y�%`/)Ē��:���K��Qy�8%��9��+�P� j�5�� l/Ƚ�D�7�jA� @�Q��N��^�T_�9�{bp��g�S'N�67�%�bN��FF�uYJ<�uƔ鑑1r����܄W������a�^y�6l�����UW�a@-�R��]Tɸ"b��HPL�=<�D煘L��ۮ]�Z��䙟ly��14:2�c~O��9t�h�� ���Y�%K�?O&:�:�s3傽jժ�w��ݹ��-5cŊUTҠX�=}���[�-�Y
��'���?��?|���v��Wuuwnܸ�844��w�0���>�9���/��Ǣ��_�r%0��A��D���a@E5�������KB"HڼX�[1�´�
41��L�1@U�Xg�k�A���0�D4Ѣ�B-��Z�bZ��

�vռP�Ϟ�Y�8����9��꽔cH �$� ~Hb/�t ��8�r�R�)Ϸq�	]U��s����a�������6
e˨���e���5��~Շ���I�p�v�Z�vw�TҠ@�/eYM_��i�L|H�lXH����0���Ác�֭3�w�}���_�җ���ַ�����BT�8���G�)��ѣ�:6m�R��O|�о}�>��H����bCw���y�XM�����?P�?���E2e�Er{���FkO��a9r�D�>E3`Z�w�}�],3��TGw�S�?~����=;��I��ڭP��*�EZ���]��	}��4�����wC�*MAy�� �7�Gr���`_�.2z�R�(�Ԃ�5W�H��M�Ad���������ϱOD �a@(̲�iZ����S��sK��A�}%�~V�%��F�k$�����P.M*In0<^vB)��!�X�ל�� c�OH�4p���vG�R�iJ�EyL�����܁����Gr�B�?qi��"�͛7��0���ns��0�%�[-��A���K%�R�Uܴh�x�$%Pl�%rY�yC���-݋���)h3NU��>�RK�af�0��Z4�0�HQ\�5I@����ȏ�N�|�]�BA��G��MMN�x/]���B`�+j�;�؀��(*_
JJ�.�m)b�0[E��)!7�<�
��R�w~r'�?L�vt_YѲ��b(NPK�Z����ڬ�eۣч݋�[�N�b�䡑a(Վ��ŋ=ыO�N�5�H�FD�;���@ɉ$Es.\�	����{}��E��:BQ�k�.hl<��ӕ���_R{|� '�Ot)���n�B�;�b��c�����3�&k�%Y��1=1� u2}�/_��"^�
��s�=�;��\>39��������M�C�z�5�@�x���C-Z�Z�tَ;��T,.��Ѽs�~d+�Q��bnh[�5�"x�.���N�c��z�;��&�j�9m.<5�j�3{�~n�9V�"�Un�k��M�p!/V�z�S�C�j�A��<D�Fs�Y}�|����2*�x5xͦ��+yⴲ�र��i1�p d���P��|����ͯy��~�mҟ� 0��Cǘ�� ����>�*(��c_�4PK�\ @���d̚��?��ON���?�����56�������k�Ο?jfj�X��L�LC}㼖d&}�u�X�l�#�=��C�>�:�s��#��@��.S�&b�	�A,�s��P.I][��ɴ'�YCk�7px�/��}�~���|�U/��`�c�L�ѽ���_��_��}h^�<YpO,�h��8x�#�zBi��@�`��,Χu�Pp(�hJ㈁�:�x�\.2*jW�A���Y���M|�ɋ��Lh+�[���{���9cbۄ?b���$�n�ݘ=�o"�r���.4")\2@W������MʥW,(�F@Y��cn����.��f��,MM�3�:ͷK׃����4��,u��%	������<��� !�v����@c�|��O�[q���|��p�ɩ��l}*CΉx�![/D!�aե3�|�0��S]2ܶ��y:L�4����h�o�z��)�
���:4:>.{~�����n��c%N�w-��t*�s�0�3s��/q+��_[�[������:���6g��y�=�",�"!�?>:�i�Kg��U�!��p-F=NիҐ��l��X�2�o����c�]Äg��HZdb��10�b����X�J�~�%�%-`2�~�G���ge*����� �K1�
2u�&X&łi��"*/�م4Ǵ(��S4)������2AZ��g5X�i��_��=1��ԘUt���taz�cAw��e������e����'{��쒝Jס��SS�r��F[�������LNN�8NQ���;�5S�?��(z���b?�?]B�t	��?��N'e3Z��)�,;d�q�L����j���PWW���=y2_(`��66�Ih�+�u�ha�� �,Y�P_O�8����3�y�Ru�%��山���z�����oB>?�� �:s���#'z{�@ ��%����yP����:�l�x���b��~�u �at��(��/;�wO/k����-��'���} 0�C�E���L���b���z�Co��k���D�#�,�ҫ��6		�e�-?�S�O��̊�l���O�WǙ������i���+'(����9f~�!
W�'ǭx�L#���k�:�B4m*��I�M�n6� �^�f�:<�Z���+��o;�3�$c��� M<�FÀ�(˩8�u��O}��+_���n���+z|����'N,_����@������]�����O��O`��X����	����>L$�:��%iq�iZq�T���(�4�Ց�hՏLR~L�={��<�s�wdw�	tf�������_oj�R�9^���aV��	�
B���5M敞Z�lYOO����9 hf&���U�+7� ��ۋG�(��*���_!+2B�Kɢ`3ԓhK���E6"�UBX#�~������`2�ru���H<����ҙ����ؓV]���S}C]����63Cn6�Z��];w������1�R��P��,�0��(���
`���rB2��Kixd�����G��M�T>y��C#��u 10��SH�&��%!����=^|hh�+V��t�M눊��$�ݥO�m���>g����E�"?�ʒ'�&��$t���'U�_��C)��eI��K�G*�=�)N  ��'w/\����B�.�)�E���@�8%.��.+�E�%�5%IVԂ�D�e"����scǓO&�y��kHNY�G�2aJ��Ib	�j����NV�~����1�\c��K���2F����%�����L2�I�R�)ᆲ=����-�I�]Hު);�U��FF�/�qY�v���<�������fㆀ��s���� l`(p�"�O�Μ����-�+m��m�eW�V^P�Rf1&�M�F��:4<<��$��,��ea����D����O���o�~L@ ��K�B�Z֯G�B��絴�*,���_!u�Pl���)�����}/.ǃ`�:pP�A%�UH|��w��݋�VU�WjP�F�s�A;�j�#����@&�aj�̹��j��kk��:�7s^U���`�9btP����<ݝ�*��-�~O�	��k�b�5�5J�e\�J��j-�0��'h������
�E���\.��3�3���K��<��J�,�ӡ x�� �#9�<�	qCNm��;X�俙"�O�]@��#�Msq��4����X���L��f3##c������O}��;�l�^p���t����wV���V�曆��x ��ޏ|��'���|vhh��g����0Y,��מ��$&^�s��L���4��bE_;z�����=�^!F14qߘ�)$�b�ݹc����-�<71>�;��;7m´�
���������M%����'��`3עiƈ��`�Gjk�)����ذ��˩��D��=
�-@�-�x`��n�}-.DM�b��Q�0��I`�#��ф��	�95MC�G"�L�	`�����lD�y���r�9�X���׊�9�|���س��%�,E��e��.�̆��B��c��%I�Ǚl]c���%f�moo�X����]�x{W�ҕ��_���ĉ^<��APo�@�M��ٺ4���.[�rɒ%�?��r�J��^&��rVz.O޸���;��676�L,>�n`���̳���3M-���cǎ�'���Ź"�v�M�L[�����N:�Ɂ�;c��������4ز�:;ӝ�<ݯ�n��3f� Ni[��m���������/U%U�ʑ򓥤�]e�U��J�eH")� �= =��ׯ��Ý�9;�Z�9��{�{�HP:����{�9����׷jW�^?{��c��c �7shd�ox0�/h�Y�噁!��B)4a��� T������ �)��Ĕv�|[Z:t� ,�.0��s�x
F;�(�x������$,%�zJ#N�Z����-��C���=�*T��������/� >��k�a�j�־}��n��'��ۊ1A"B��M��fIr��(�]�1�=�h�k��I�V�h6��Ƣ����}po<ū���W�D"_�d"թ�+�b�`����Z��%��aω�H�O#��('n5_������6�W5�sh�2.H'&�=(W%Q��+ͣ�Jg������>U��������ӓ�����:�U/fD=ς�����?�����^z	���o�淿�mX#�{/]��ǘ�;=�� �8��K��T����lrrZ���YY=�FC����J��\�+���(�#����!�F7���-.�����,���$� �5�u�im%�Z���q����~�sP�`Q`/` ��*@8��޽{�{��g�5>pq�Vڰ�h5Y���JUK%DH`����-a�B�#�-��G$���#e>;c�~/�N���I��?��m*I5?u�$��_`����'k�}��uʗ�n��k�R�%&1�^����y�*����Z��*�N7wM�J��K�������3�lE��B��<{+�Ż��վ��w+˼�Lj��9�Kqմ�E�:���~�*���ECCC����(�w~�w�����0ڞ���{�G��}�艓�J�[��֋/���ۿ��0��*\�ؠ�"d���*M��i�e���i)�3ZF�K��E��W+�4mI�����6_��׿�@��?�<4�b"lTm���뀖d����r}�=������+cb�E�ujZ���6�h7��J�mQ�ȷp���dtr�4,_��D}��OCN��ɻ��;�xx<`ٯ�k�v��:�ig���Ņ�I$��P����]��)e�"鐝��Z�*�	(ָ`mUZ��߿ffW����Xm� ��*h�����B?���LR��~�3�����[�L>0BP/n�G,��A���҅�p��_��_��-�b�D|���O~�RV\���;�$f�^Ps`��5�ݽ��ۂ���q���7�}�6^
7A
P�~�3����WqC�>;v'<#
r�d�)�����rE���:u���|vh��	&���U*<��p�%x/6.�F'D�P�9sfq�>v(������;w�LMN���[xML�.t�*Vgbt* �[;�(��B!��X�z^�}���q����2�1ua(iL�sA��[9,�t����bͩu���e3jr����p*b�4�Y�ɘ�
༌��<C;��SO��YT�(��Bp�g?�)�������^^�2�M�˭��H�Lt��>����~���O�}��ϼ�"���_��+��JZ��@�EŐN}�χ��]��%�,Ȇ�>n򐞶[#;�g6��^8|�0y;ΰ~����C��3�<�������w ��4ӕ�UV�b�b7�]N�>����/	�O>�$��G�G�O�:���|�j  �VIDAT�7�x��A�zO9���='�����wq[����'���N�����C��p�@�]������	u=�^�R����1b��x��D��B����hzoO&~��L��)v����:Ҽ�պ@��D����D;�đ��,U�M���1t��mS�Si��5�e�j�����R
�e45^ ���}�k�GGA���^��I�V	#l�FRo���`�����/^z��~�B����c�^�,�,���+�z�p�����`Q����b__�٪�o�M�v��F��.0'%0To�&^��)ph�|��$�DJ�T�����4��{W�OM��E�菾��+����rY�VW�13C���}��h�X�;48 ��F���a��SC5�����՞[@Ʋ5�p��@VB��1���f����~����ĵž�1�Z���z'��l]|�ç���];�%$`�)��(�S�=���F�Dx&�J}�*WB�Y\ل�?<];d`d�3����P�T��U��͵5��*��������K�.]x���N<*�V�/޿'�b����s� MЇW7�et�Ǯ���?>
�m�u��� <(�x�z�����+�������?|����ap@*�����}LI��X�ۂ�\,%ڙ�!�9�������o6�=��5}�_��/�/,�I5h�����i}613�g|r��H>0�����������րHc4���$�,�gb��>���;s�'��/Iw}?93��<rO��w�}k�
���+�������꫰à��2ʗ���z�F"�ñG9rx_��������dmj��`>I�!!_���8�(C��t$=�?Ћf��=�<1�Q�fq�|(0(I��~��P�VB���6i�����I�J�QO<�+A�E?��$Q�����Es^(s�R����\/�Ǐϝ,��G?¾�J47��C#�T�%z�+*�6�T���ͭ����ɉH��PY``���{���گ=��S�?��׾����������E|��*�hr|�J��'�������ٳ���Cb�fQo4����DZN�<�|���L�i�~���llttc}�E-/^���۽��^l���WP��z�l�J:{�����z���{����G�����JU��_W�Vs�V�ъ[��Ү�Lc[������z���?�D�b�¥#+��>�^����'�杸5����}7V�`��j2=�;N�eTW: nܛ?XEkC�����E��ߓZ���v,I/p�t|T�'vx6�^c�x�t��z��&3Qo��f^�������ԣ�%����8�M;�*S�*r%�'���������Z�|;	�h�6:�&˰�ݿ�w�9��_�� ڱgv������)�N��
��\T P6OUk�}E[��Ň��*b����.���~x�o3��O�!���'��=�A,ށԿwwQPY|D��A�Ưj[�x5�Y}�ڂ:���:���N�fS4��I������j�:��f%�Y/�E�j�^4�^(�|�]��!��Ϣ�}��nK�ԧ�1�l5@�R�t�^�n]P(�y�.�m���l+n�t�BT`�pC��k�\i`�N�ӧO�۷������oa�XQ}
�ֈ��\&�a�Y@*�#c������W�@��W$O������8ؽv�����*�v��6&uQ
�@��9��Bpc���$�b]
U�SG��FNB���d3G��5
���16�(���0 ��|��)�F�F�������{r�b�PŞz�)��PkĜ������;w��W^�I��7~�7���`�cT���:o����/���/|��P�\��/`ɠ�uՌ�O��&F1��V
b�}x�����EYwV�zg�3��M�<g��>q���U���V3ɸ~���S=��ӧrYsn�Pkw��N�y��#��n�ً�����R,�믿.YV���x�$k4�{�u��j��1�!��j�#���q��c`���8�?��Tů������o~�������un^�=11�Z�Z�JN�?����I ���P�Ѭ�� �nllac6).i�>��`�_b/�g9n� j�8!>���/�K_�������X°��A{�̕�%������N��$�╱yA�Zȿ���I���`�M����ݞ�N������E���O��s�H��#��MO���[���.�d�_�J�(�7~.*5��A�l��-d�B^�@������#��-JE��^(7�o|M%�1��a�U��$P5�X+��B��R9n5�p�X@�F%�.v�P`�D��[����G��h&�Bk�#`Z&Ҡ75 M2��[���L�7����6$��ui�.
��a,F]�l9q����u�3�Pt��f�a��&ȵ��+ES7���{��u�����P����������,��R������?�r�6L:VA���Z>�����D�����ͼ ���rղ��n�d�1��&���M����*7 n}'j��|_|�A����fQTl5*�b5�k1ȩQ������3;�w���Ic��4S��`���e2�S-T�1��頪I%^>�(�}���)5��#�#R���P� �Vr��}-ݒVY�.d�fR7�����jj'v�ݐp��>$֮|p*���}�VK���K����۴�Eh���p�//�JP��>1Mq�B�iX��_K����BI!2��Q(��y�!^P^�l��'N�
����=�OOL牭��υ7n�����ơ���_��<{`�������3�����{�lo��{O?�� ��}w�%�2�t>65mf43�҈GJ�۵���P~�o�Z�J��i���AQ%�<4�w����B�M��@�ꭁ�q��F���%`*=>�*��p}B����Q)������025��Ri�?6��R	4�l}��������&�|c��KI�r4��(���2�+�MM���Q�]�ֵ7L�����ڿ�4:��K�.^�833��/N5���X8*�O?��<��w�\�q��?��c">?{���˯���#'=��Y���ؓ��9zx��M�H�^��&�+{�\][��9:9���Q����h�-910�%xWO�C��DZ�װI��M�r��7�-oeL��H&ZV~���e���'�+��/<>�
�_"Ϳ�K�}XSq~k�zp�@0&`�5���I� k�q#�ǁ�󒊤�J�05 ;5����I�1sIu�|k��(�S�L��"I�m�q���r�/�G
��/]�כg;}!����ϱvk�K���\1'�r�O��Dˏ
E�qR�
Ќ���lb?ZY��­;����������={6
��={����_�/��ß��'���7~��_���� v[���k����R��8��9�~��R��v��I��,� J���;�Y#�cWo\�&1s[e1��������d�a���'.\���u�ak��3{�`�w�������
�ť{ T�vxD2����*�����'-�����/_�Zoİ�ŏ{�Ql��v_��[��z�r�5į��*mP�V��`�'2�Aj3�M)R����ò��%~����i��M�T���FO<��6�}��OI�ci$�<�˲B��[ ɰ7)��vR���%~A�;C}��Ǒ��<��Ҍ�T��&�'Q��S 6_�*H�cE9��}�cG������S�m�Y���d��&��&�u��+�u�����躳���h��~�����UB#	+Z,�j���4^
����v����8�w�w:����?���������N&�B����]���v�'��gcN�4N��=��F��I�:&������Ӫ��ȑ#33S�X	X���<d�]���!��s��Sv�����e��y%�#�M���dM�hV�,�u�(���9�����|r>$gug�FՍS����`<e����Uzxߺq��b�-���ؘ�IC\\,��A�)����o�=95��,(���0����-!�@�p��Ѭ�[X��������������;�?8�x���8���kx(s������C�5Ֆ[�"��+V�21_�o�
ak
Br�K���7>U.|%�\�F�z��m%��XeB�-B-��l�7]},���A��Gy���+�s���y�&!�y�����	w��Ҫh��ڹs��vP^q��x*J\�]��������<x�εKR!x���Q�4)3�+��H����K�ms���3��9����u�.�o�y�A���G�2��cc�M���M��EOn��&�%�X!V⪶�R�����/?5=��! �3{H{��J�G�φk��3q�@��/_<q����?���}�K���Y����g���g^}����?��k�4����cMWW�q�W�:Gc_�[F�w��8���Ɩ���|��O��������=�k���ځ �0ʍ�F3�W�^u�A���g"�1��+�yk��;ҩLAa�(;Q{����>:$��v�E�;)�����j��4{Lֳ�=��N?��;��¾u�~FL�}�>T����n/�Nz�}'�Ir��ي�o���DV��'0Y؈:�g:�;X�.8�R($~�4FI�Iߢk��ARf���AK0��i716:�W�ؐ���:6h�h~(�-�U�^1M�n�������������͛����z����Z7D߀�e�'M�rj�t6-��[�P���:��i�l�
s<4$@�G���o�lI����6�Z ��#���KE��F�^(���cthX�ȌTW�io/��33�&J;��!�t�N��|A���U#^��arV`YK�lF�+E~���r�����2Z���K���l[� k:�8s�!��3}�rbS���>�Ǟ8Va7
�J�ch`���o+��q��"�)6��{˸�8��4����v�]~���-Ƀ޻w�f���*�Br���R�2cfz��b��D�
��8[������j�!�՛M�q��S$��g���'NFG�5�Ey� ;�������m_�F�+Y��Ek-T\e��SǵZ/e�N{��M֔va�<R$�����8�� �_[+���O���S������0�
$�!�ai��;D
 ��{�(.�O�5<<�W �8�0�[�[޾��P-��f�Hٱi�lױ�d�w�E;	S�,�ȿ�2E�c�k�W�]:S{L-a$`��g�3!h՘&�-�h��C�R퀥��p�%.o�5�I�A
lnL��R��d�)&*���J��ѣϜ;���^W��2:9)��Z48=1%���f��5VO�,ŏ#�k�������p��٩��;��9����{sui��짞{��_�l�P�r���R��e9^�>Df`pxbjRB���駟~�G�0YM��X�thTx��cb�� W�D1Z&���1�����?���}���;w6��1��͍ͭ�PS�gg�����s�����)�,n2�-��8��j0����𭨉Z��	G��P;el�)����WA֧���EP�ے.t�6ex�d/��[�zk��G1�۪��q�^èK�����ߢ��K?3���ܝ��ϻL���}=��}&P36a��I���D�[�g-��ړ�P���m\jP�Q�j%�7�&Ƶ�&����������&d�(�z�����Ű��/�������&+� _]��Y���5�~�~FUn7��ϲ��b��<�S��f7��;�;�"5����7�W��$=X 8J�j���շ�#�D��֔t*U��3�k�N��k�Dm�Dn`۱�{}w!����Z#���;{/%��]���jÑ�m��Ů
]><���UAK��������ב��*DR�}<>>}�&�����.obq=�@�b�4n>3#R���{�FGǨ�`�O<v
<�>3j��[�O�h�{.���j��Q���F���e�E�0<��q��H��s�pCl��=���n
3��p����U���FF��o��[,l�vX�=������6Z�� �!�صª˾�b9��ݵ��
� �̍�����r>v�(URv��|niқ��HW־�ׯ���-0�U���9MA{�K߱�{7�K����=�Q$CSG@�����W�2[��:w�����+nU�C�g]|���fg���d-���?���{cx����}����x��̘��u)�iԚi�~�J�i,������3���\�ږ^ɗ߅�thn�cz�����}��k��'�{n}u՗�������	C����Z t!Cq?�<�
^!_,��ͱGK�T|5Uj�%1�xƆ+�9���3ׯ_{��q����^}�}A��|E�1���������onnlH�}�ο�_+�Y���><(�$-!R�)Hy������u57�|�k\ǁY�J�\����ߎ
���E��h��hl>��#`,iR4�ڒ���0�W�k%ڗq�겲��b�;��[��3�-B�%���uh�Zv���mr���ހIL<m�%�c-+2�)���Q�K����xzJ�ǫxL)�Z��"�S }Pk����$I����r���\��B����#A�Dլ�k*��xP���A�;9"�3O�����H��Y�F+��� �2=���	65T��'���WW KF����O�lU�3㓡��Ǽ��x�4��>�'�b���2l��R)�J�9�5�����8���	�AbL������u��ݎg�w����<�[{0s�T�Mg�l��YA�p<�|A�,�h#*�sۍ���M����χ�z�Y��0�h���Scc��w��cŉ����[j�4 Z��X��▙�uw{��w����y��|NP����@��Z��S\B0�>���������O�p`bj�	qR�צ��b�$�Хwk^J&�W�@����Ii.���>��V,ݟ�="�"OE��)�D��/��[����YJ;�E�H dw�h�3b�2K'�tF���@��d���K+��Q�nJ��<�؁��c�Ix���x̶��[M�QR.W�}%��Z,�?�4Z�&Ub]4{g� F��?]5�^o7K�5��?��rЋ�w������h����hy��ǒ��y��[%����$�A�E�o2�L4�-��_���<�il-Q4Okꃴ�@kB=��i����@�o�Z{���#�O�SO�;�Y��+�]Ċ�H>��������Rd`]^i�F8�x$T�Ĵ&'��DS��\}��O�x����N�>}�ر���_��Wdk�����0*mm�6+ͽ��������f]zo�omJ�se����?ǃV��@��F`����AP��k7<�%�s�l����������ϒ^��D�c'O@�Ài��<}�Z�������o�O_��׾��_���q.�
���6����Ęi��H�K5������[�>���6f�=z�M�Ƙq&��ƶ,���fIT��7$���^:K�6xm2X��C��G�l�st9�TI{��(��	*�SL�*Z�F�u�=�,#'Ț���eߒ�vE|Uyg�C?y=���?�
���3����T1 ���{�0��ի�P(|�8?��Q�*����L�؈�O�S��iSJ�$m�ա��Y��C.���j�3��&̩O��bt��%�W2�D���z��G��*������ko�s-��A)�l4�t����M���%���gq_Dyb�he�S��Z�J\6�vcV�z<p�+]Bu�{u�����8��I�-]+.����%��-��F����w~��\z�ń�T��U^;j�6|�=�F8�a��O�4�����H�J���b�gffX�	���]\���""�'W����l`�]h�+��3%��T��Ӝb������f]2[!.(7;�!�1�d�^�� ���b�ʤn�o��G?���,:w�9cv]�� Yc��A�`xC�)�o6���Y
�v�R|8�5�a�A��*0<����Svb����� ��ˊ�haaartDb�u��v�+� �R�Hh����{U��;<��Mv�C�&ٶm�����&q�~z*�M�'6��.k�l���e'�^c]&����˛�*�����;w�|�?�r��S��n~��m�|I�X����V�Va����I^�v�k	|��(`�+A����T���������駏=����?��c�x��^��}����m�K���+�Xe�?�w	�OJ/)B���:���Ug�E��3�
|�ҭ (l�64��i��;���Ac###0�^y�o|�/��ݽ��x;��&ֆoD�$����J�3��g���v9X5�`��v�ك��������q2���S�Ώ��K������8��션/�ne ��7-�s0qZ��R���{���^���� ��]��խ�.?ՙ��W�hX�Ȅ��S[�忘���a�!;/�{����:MB#����I�:�	��Rm�F���Y�_.g''��~;V��U��7���b-�Ǌ"��e�����P�����{Y���������	�Ζ�²�J�=�^V~yj"��1*#79�<�C��lՇ���=~�����P����+�-ܜ���y|��j�a�	�B�Mu���߃45u$����LODg�i��{�V��(�f��8�ͪ�!�J�\��P>*%��uO��]��m?X���E�+����	'�ʡ��Xe4Q�#5�fS�+K��xΨ QJj�.�����~^B~ʾI�����:��G�X������N�8a{����۷jY�Ѫכ���P3$�A��0��RdQ���eQ�P[gz�z�P5I���Ƌ�� 9}�0��믿����+qF�FB���͢�hoUc��@��%Z���
F�9��\��If�BZA�B��Ɔ񴣰�19A.CJ#���*�0#U���ԭYOQ��L"�0��G�R��E�4�+�B��*0>Y"~%�>��y�U�F���(Sz�=lvɭ���^��n/y�M�� �-����2�!љT����G�M�):r���|
W��M�'F��7�� i&��FX����+TN[�ڛ[�X���Q���^*�~��Ǐ�7k/����ڲdL�y�UV�����W%�s"��jKϞxd��	%�3�������j��(s����_��?�'�ƾ���\�~mz�܁���-?~�ƍK+�M4�;�ã#�y��|ߺ5?5=�/s��$@�!��U`��Z%==9U���~��Y����k7�������¾rY�UT��;�
E��x����wO>vb�opmiyqaA����ۈ��vD҅	a�(H,@�4���k�8��N*!iC���4�X�e�9O�W9N�:�2T�j[�i�P��]��2ц���Z�&���M��;�"y���Oһ��gc؃TN���t�ݔ0����o���f9�V�y�.mZ��̵F9�u�[�|�bRVr�`���0T�x�Pp�pa�`c9vF�	l��R7������(TF+a+C�U�!�d`��'T��*;��S�\&�1i����ɣ�f !n���l�6�b_�uھ�b�?��333o��f[0����`&:th��G�Lv�0=��;�0@.q��\��CU.̛�HI���Ȏew��j��|��8�?�]v�m[hi첕yς��][����@�N�Ӽp�p��֪b����6�adT�6�b�C�8u�~��>�����_��r���t�;K#�,�����K	oC4vfd;�Z���-��/��(O���ڵk�X0���Sǡ���8M���G7��q�*T�����ʷf���b��ݭ�e��@�6W��j[�(}
r��q��b�7�3n�&��zu���F�7��љ�?���P�1��@]���XO�jG��+�,�繬�s���L�i�@mp���ۼ�0�d��)*'�@����QJ�0L2��2���ŲQi[*h�p?�����7��NC)�/7���-��o@r5�����i��oK�w�����G�c���h�l'���B����J��1���O~B/�������//-��D�f����{/���/}E)�����7i*�)���ǝO�<��$��P옎I�?bj����م�E__��?��3g���͟�)x֏���-Q��A7�v�=�ʕ+0�\����lg���A��"��ksU��Aw�~�u��^�e��ݴ��� S��ts��eY�vf�JьLW�K�y�4f>�,�s������#u�گ��__Ĩ�	��D�R�/�I���l����fs7/�{�j	� z/������J� k��No��>�i�*T�x��0�Y��J����{M����U�/�J��������L,W5y�X��a��r�A���ie�����(c\�X�s���7��Ϟ:��y����C����G�[�m� ۱k`.���痗WGG�˵�*��d�F���(���bh�X����,7��HI�^M/�_�K��8��Mq��Bx[1_�G9����64 �[�������W�����\_Z=r�����o��Vymkzd��Y(����,7���B�Ք,�H�m�O��zasig*��X�)V8����
*v���6�J鳩�1!�(�	
�j�>~j?�#$�l�Q�Y���Sus�c�v82�č�*Wӓ���\��o��}� � -��[}-w�U�0�(K���TT�/�!e�V�J�������?��e����m���n�7��{�j<�Vo�Q��Á���K+ꍐΟ�g���J��L�M̞�[���B��r�\�\��;T���|�Gl��a0Ph��q�R�C��΁�& LMM����h6Φ%��"��ѯ��zK!��͍m�.U��� ��Ay�	����� ���l#�M�|/��/�*��;X�V��7���	�f8!X� �a�4��>���E�l6�Wdl]�6�����d�mll�����ޣ�QP�2.���*�[S��0{�lDA&��JL�6�{f'ӥ�&Ϧ����^4���]dځ)�%&����0"`����
h�
XK˺%�aJO����i�V�J���dO�'�!�H�)�9���U�<�t��xӾ��e��,�l5�EE���F���n��`u���3���|饗n�YlT�������7*i/�PM|�`h�(����i��[\��o߾��	�Wml��T쟚��+\�v��p�R�?��so�s�9>9�d0�.��V��ĉ)�JsJ���7�;����F~��M���?�&��#�llm��T}Ƣ{%ڜ ��ޛ��^[^�}^|�ſ�O�imiEr$��f�g�a�����4R�v6S�����;�`������l
�A�J���Q��,��в��Q ��,B��)�
bpSO�<�5%6C�1qr��G�85�>,�&K�;�3;n{�n��q���i<꺨��>jH��;�Th�sjB��t\�\�'�ަ�����D[I��ά���+�NLC�S�N��e�J.�˯`�.--��������B�?�����F�'` >�ģݯt/a��m&И��o��f}$��Ⱦ��g���9�b_�k��No
�$�%"�_�*k(g����z�ĉ˗/�x�}�X���xSB��sm/����M#��ﻛ�v��.L���4>
i�����7��]��v=�A�]�Wv�[�,�ick�&V 5�� �H*�h��/�l��2/��Y,�t>�Z[?��u��n{�idn�V����
�4@�|pp��ˮ��L`���7�4���r��F�������-����!B`��[���-�(�����D� M��$�Uz�8f_2�F�y��{0js3�:���� x<���Pz���g6��T9�;�2�,�&���=mb�y=�գ4���c�d(�j:	���0�D����j"Q�B��?Y�aH�{��k�~��z��K��I�93���j�L�;c���l��ҷv�80��1w�I/���;2��5���ʔ�o}�[_�җ����/..B9�댏�@��C����~X#��|��1���ư�(~k�q@��`i�����SlK� ��"���嶶�@~�!�Ը�a�����g&eg�����-v23���Q<x��w��^��1$��t��K����s7_]Z�}��7���(y�R]��=:�m7��equ�.�k9|/-�:��H�L|��ʢu�.���%���Vm0��D�v�����z7�ddSf=I��㽼��ѹl>L���,zt�$u�*����4��-xD���H��	8�����,l|�~�|��*�+�`9+Sd�!'Sb^J�	I:Z �lcm�h�k����8�;�Y���o���r�&ƥ|6f���4��]�����I��x����?�Kb�,���jA�͗D�5[�#���fssk2��Ͽ���s++W߽�󽾨x���{������8(HVX�{��ç}5=��x>]��B�m$Z�#{��k��=�!00X%^-�i�$�cMw{�
�$�����G��0;y/�ߦ&Ab�줪�x7�L56�wRר�ZB�bk���35ha���"r�Å���Z5	��QqP0�t]��NuB$6�˴����j���C�nnn{b4K^?|I����@^}pp��$����A�\��|s�>�!�8�
$D�����W����^�2g�O�ƨ�Y|�X,~	B� �4arFi��bd��<��'�i�3�_܄�R"�A�쀢�atif�)e�rnn�i�����x1�Il�N�Tə�'9D.���4�/�"ĝ��m��֭U��/d���k%�Vl2��8)>����>�\1����."O�h����{=�%�������f� 7�q�i�I?	L��+�S��γ@��Yա�P�t�!a��H�SF�~b�(t��(5u�L,>�$�����F�o_~������G*�Ko��������P#�K�H���-7�W��\�U���VS��f����.���u�P�U,ت����6���$����	�Wã�/H����&�jv�_�ֱ�ك*�K/��onϞ���$~�W�WW���={js�ؑ���[7n�>y�ʕ+P� �
���7E�����觞~vdx�R"�Z��A!)����3M��T韴4@��,��'�b6�;V�c~A�2�_DC�m�ٖF"(؃�׌4H�4�Pq�z7W�t�!�����w���}@"f�P�s�^���.����V�p�t�����w��v��_������VW%+�]���z�6u�Ywl6�����D�_v9�ddD�V]��a��;v�瞃u�����IzzZ-if��O��.V-�ڳ�A
R�V���u��P��^m�$ߛ�V��mE��yBQN��D�.�/��/>y��s�6��W,d�|�T>�>��+h:m)�_{-ں�g�>n�17��8�J���^����^��ժ�[���t��X�6�rf�0�˺�6VWl�U^-l�P#`���)J�H��L���3퐼�$���#��O+�4��x��h�T��;|�{���gffp���X`l�Ye�h*=��K]�W���陬�#)�Pg�_"0�f�H��x
Q�9d*'��09�'d��a�`���k�acs�0�E����S��&
�Klw<��f�� �q�9��OW链%�K¹y�߰A��4O.������@KIL��Y�K.w�e��L��܊e��ގ<$AZb���I�:�;�m�S5�yeWvt�����{�A�8�e�W0:|��իW~��~�W��O|
�297�w���˾}���#(��CbI�`WYh[����7'/����-�y�������JJ��etI��������dt������F��v�Ν�/:t��������4A�k�b����ӧ?��O��]}
\S��ම�/}H��k�l_s�)�$�����ݎ�'o�.�9�������,�R���VeF��`�������Md�!��Ie�a��c�u<�Q)�Ij�Z�'�BL�hRO����T{��3H�2�l�w�&[�J�3&�Φ枕pNM)�!HN.�)s���z@D�+�<*�Ɖ����3��#'{��O���W_}��C+iTōZ��EI�� �e��4�G֜N���]쮩s�� K6��˼T�M�B�F/	\wP/��_�K�ܾ5=1����?�Ĺ���ׯ���p���U_� N;P��g�۾4\�������S�2E\󲞭�h��iA�i�-_ݖ�k�s?�el6�PZ`��2�*Ȟ=g@�^����ڼ����wq���G�jz����,��磐��O~���i�^�o�(wc�v<N�hy���aT ���3öx~�԰j�� ��+NW!@ڑ8,W�JE��:��f�!Q"�3m�Y��D�Ǉ��z��v�@+� �^��Ԩ�Ѥ�� q����u;��6Obh0������:�
��ȑ#�9$c���nl�N�¿~���:j�T�p"gΝ;��.�?�V�.�����5�X�2�_.��	[aN�lA+�	P�7̚�i�T��С����Y�!n�o^�؝Mv#���S�
z�w���QdR����,//mmm���'~p����%��$iy�����2[�G�� MJk��z�丒��Zz�ݟS�����f�w�G�Θ0�DZ&Cf Wj��0�����_�����'>y`����޺v�M�$(�J�(����ط5�[7A6���a�ʢ(����\�U�2���|Q ��lUs�L(�98�x�!S<�V���a>��*գcc�Jmss=���}�{im/43�,Z�Ϯ���YV�������/,,|��g����_|Z݋�����??X�?����޿sC��+Q Q;ZS���J��[�?Ĳz�y��P��nrb��s�M�yȉI�C�.�Ty��n@��s]j:��e���ui�2����+�M�T�
��^ז����	�w���h�;��J�n��)��a���=�1�,5���;��"�6�VlM/�y���Pˏ�0����ݻ�uA�y�'`���reqqqiyU���t=^�`�<=��5|ǩ���7�X�W�RY�KyeS}����W���;t�����ǰ�:av��{L��n_Z\dҌdU��<ȴ.W��q�;d���~�/��&�M�a�V��4�]�kg�we��w�]���a�����������}u����?%걽�嫭�կ~UQ[��l�����������`���d��cmD�$+G��>%��|�^�*&�x�������[V��`�����{,u3d�hj���g��gА�Ge��|���	#,[[U�w�4$�C\��l�D�{�v/`�z���Qŷ��g8p�������Oõk�Ѕ����҈���m��V���A�3��Ax��8 {�p�lEd�i���p�vd퓻hi�a�+g(���`�e:���"?�� �ݶ���no�o��6wd����mL�G���g�kB��^}U����̐�\A�7�o��u_��I��Rw�'�X�1
O2���+�L�jI��+@:��ט;(�K/}u5X��#0���g�ǥ�t��M�\�žLgϞ��k�}���|u�֭g�}�W~�W@�_��1��^ziiiism��H���0<��g�=X!�f뇁� �5�w��i���p�.����*^8��g2��y��@6���^��h��q9C�>���v����5�~��u��a�C���e��B�B+���P�i��79G_������f��?��� �"�YgBFH5��Y#t�,�V��+�O�Cb���-�	��+�լn|���g�>��{��^�8Qע\������`)a����v��,�:�'HS�x^ә3E�����k)�Z�I>�v��C���ك=`�~l��g9th����{�/m�oȎ�J�&ulh���%�Q��������`��u�x�u�q8)ش|6�M�(wz$i�*|�[��@�a2�l$a� �:�#�����]G�H4~���@N��ҊYU+ܮGL�N�&�gΜ��tx���OL~�s�پ���zH����Q�=vq�2�Os1�L��ٴ^ϤU�M IqB匀�)�oߦÀ1G�f��Aa��r�y`l `2��W�%N�US���(Wm�zI��iԖ
a�F���t,�Cf�+	$��`&�Ej���3���t�^�eq4����C��������Ҍ���V�E���g�x&s���
Ƿ^լ��Z;~���E��G<�	��!�^�ާ�uX��Ȭ4��\V�y`�n������u
��
4��e�w����L�u��:�Ĵ44#w�H_*L$]�ѐ�R�b����O�|sic�g���ڳg�V��;}jnv(g��m(=��(a�V��W��JW�-��w�V��i�*�L})l����H���߆��A�c�s8����Ð(��VV�7Z.'Mf�,��תh�	�1@,��H�����_�e���w�S���گ����w��˛[�Z=T,�͍M���'�j��*��86�(Q
�^��̺�^6k����;"[�6a(7T@x�d��׽�3&�������Y��~����-?�P��u�:GwR�{��^�}Nm5J�0kPHO�e���U��3[�s�=	Ch�<�Gj40� �n��Z��vK�$t��~IG��Ƈ��9X6��h���?�sgAЕ���Q�f���Q [g*vX/��.I`R��V������Ӿ��5bA������a�K���>|���իwo�1�l�}��֚y��n�=���Dz���˶��x�N:��!�3'�:A.u	s!<'v�g��.蒗v<+�?����o�!�[-"�0� �KtS��X�����-���i�����<���_���!�it>���~�]%2�=�g;�R�Ч���[�"&ɼbL�W����)�K}��ݻwy��hԒ�(��MqB@�a���w}�x%Y=��7ے���3�~�$�@y��8�Lt#4@���ǻ@�b��ӈ���hP�:�(�޽{� �����a���t㶫�r`��$��g��_x^��FE3q�ysZ��$ɴ#�N�v��H���r��݃���0��5��V���S�T���A��,�ܲ2�""n| D��0��{2M�	��V�E�d�T�����Ư�<�4�D�[��M@[����Œ4���,
}�$4�*�TS�r�> $�UBG,��a�������6�����z���K�L�)V0�,�dt�a0`��I����v%�����W^9}������}��Q����k���{��[��m��\3dĝhŨ�,��2��2ɕ-1vt��F6��B�Z&���\c�cyW�#v�}��K	��*j������DX4���+$&���lO��P���v֊v}�s:����o��o��OQ�N_<;Ҵ��b�IaH��8њ>�`S;R0|_���Џ�I��"�"?bѴ��N��	S��JXG!�T�:όEU�ʋaĭ83�q�Z���%��kF�N�KR�2d>���7ŵV�s����pX�+���7�+kCC�����,?���;�ܼ{�Uo�bq�=ٺ�����0�틅�f���H���X�u���),���Ni�U���D�@�$�7���g��Ԣ�k4M�V���A��[�z��G0ٶa�~�3�L���ͷ%���sk;��j�m�	Ӣ(�Ll�\�'�8y�\�Y	@:�>H�&��ˬ��G� n,OA����������izA0�V��HU�s��@]o/���������5�;�X	�e������@��z�	 ;����e���b��u�V��l��y�gH�ڗ� ��A�%��Z0I�Q�z,��c��u{|z*�� �7"����O>a��7�|sK��m�<A"���urC��#�SM'+U�H�+(	[���T��ˬd���bfe�sM�l!b�p���ScAe�S�h?��r��]�J5��hs_�Ҥ����@�����!IV�ßێL����UX�F]���^m��lw��b�d�<�Z�!?<�N 
���5Sv$U"N��Ys���4g�2X�
���o4�B�J��H}Z	^>j�n���a��3D���m���Z$�N�iT���A�,�޷m�j�a�S	���9�T|��W�5���C	���*h5b����%�UQ�꾀r�����X��q�DaTl[�*�rUPY���%��M{x��i�4�r�ԍ���cO1B%n��V�������Ͽw���}��K�"vb����#åm�u=6}`���޻�������l������%C�T�"� �(4�ø�Z�nnW��oܦ�Q���Չgw(��������=z���X�;=����V��Y�r��Q�Y����ߪ�r������cg�|�3��{F?s�ƍ��뿔4�zmvrbue	�C���Z�W��aY>��I3��HK;o6�<ZA/�^�6�	��W�PC�ȑ��?�:Z&v�e�)y��[�i�S��5Ռ)ZL��L&HM_�q��#��R8�<I��\�rCT�$�ıJ9U�Z�ؑ�oN�bz�3��]��b�oBc��ҍ��8	sq��Ήb��!]\E���(P�:��t'm�s쇫/wY��E����^g�yǻe�V?��%֓cg�x���^�կ*�S���E��� �c�~��Z��w�(Ϭ�A�]����f�ކ!>41v�̙��=����V��������j^��C�@A?��
�BK��po*TzQW�S��FK�	^N��*��)����k��bB�&�ָU�СC�;:999><���hԙ�-;V{ 3�l��>;'��H-�2Z�Q��QƠ8+���&YO�DA��g^wE'I�M���gu��	j:���/�h�C0;^��I<.����EҶ�]�|\t��q{7}����g.���>;==�����.�V���5ݝ�hv��=��$i'D���E%ƨ�O��9�H�r�CnǇ�?���&+�����c�f��z�$ˀ��������N|)�ǅK�t�d��6=�t&��C u5������ĩ[䐨��+:6��Y]a�f-�K����>]2(��g�:�.Sݑ�ӑ1m~G�'�1uc��/��ϜXV�+U�2�(�l��	�w��T��y;������لkq���T����޽+pꂭU���L���M�[:y��o��x�g"�@Xv�z�[c����Rf9ä�"��R�
둧����7�ܹS*�=z�ȑ#����I<B������$(����ǆp��m9��կ6�v��.\�p��u�A� ~L����՜�,����g�@��J֪Dkc�v��Deoص��&�������k~��!�Ã7N�g��7��g"O��r��,�����e����սZ��i�1c������&�_�n�J�I��#��x��G�-aU���2_^]-�m�Μ/A�<�jU!�,�V7ױ�t���T�Z\� |(-ݟ��|,����l�e�xl�����Ѭ�MaN�@����>/1iR���7;�vh,�PQ�� *F��K��׊�S� L���Zuk;��M	��������홝9q���Ę@X�w�o���K�_ob���j���3'{&�
��X+�J����дZ
9� i�q� ��o��zV����<�`���w�XZmI��ޱq�����x��$�v;��k;�hn1�(��Қv���{'qA�&��s�ΙL��Tme�]8�F�:u
���ի�0X�Q�����J�.�����\�!�گ��9�uL���:������P{���<�g��g0�^[��a{'X��#��'�㉵H�aJ����¬�/neݸ9�v��pV��p\SӾ��X�r�]o���KA3i�J�����t�(A��z�T�H��L����U�d��~��|�:DH	��k��h�vU��a.���@��1y�j�&�KS���9�J.��adS�ip�#i�"��Dʛ��
3m0�d�m�V�;6?��:q/ô�
�c��ֶLA�/����n߹�$CHp���m	A����:8�`���`��Z���˷nߔ�M���U�r��T+�B��F�DxJ��ߛ�D���V*�aakk����z�F\�����z뱣�V7*�y?	"������g
���F��N�MM���SPOV�˰?�_��ܼ{{�֭[4	�S�~R�*"0�^���IT-�������B�et�����B����a*�� cֱ��l�g��g��Y�ݥ���w��]�A������ƺv�q��1�,K���f��+8��/^E�m�I3͘Z�u.C'��X'�Pb؞/I���$���A��I�Dá���L�E�������g*s�j�QP�e{i	��ÃP)&F�t��9�=9��ږ�V�i{k��ږ-5ȘC��
0����
�$��Ab �7�z&N���(�����<�~�Y}��b�Ľ���������G¾Fv�qby��%�d��]5]1l߽w�d�rZ(dR�3�<��t��$�h� �ٺ�.��� CT��)V'��"�ݒ�=ӥ�t&�:���L���Ù�R�����;��À�����'�y�.ߧ&)2���;��F�U�<���dΪ ø1YwT��Il��Ή��{�?�7ԝX�m�'��Ƶ]��%�X����v���~g':w��(��L�4���J�G&;_��:���4�������<%L'��(��=$m����R����ϲ�����٤�ʮ�ߖ�(����u
f�X�+�>�0N���y.���!��	�r�ݮ��[��qV�+�i��}��9r�ڵk�w�`O>v�-�W�����,��8�j�cǎ�}��.4t�9���YY:6K��� ԋ����A���7�y睸��9sv4���U����Fap���b>��f���&/�=�!i�Z����"�6�|)V�(�p�|�kCV��&�~l{���e{ߺ��9ߑD��F�6֫ue�����]>��Gս�2�9s_���d�M�鮼E��"��b��Qc���?�ѵ�L'�3^�r�&�rmɠO��t�V]ᡶ��4��L��ز��MzC(3���k�Mp��-V �q����~Z�6a������z1���_,�׽8�5�7p����O=-X��Q�g��3�j����߼9�����"d
�j��N��H�~&�+��y�Ԕ�A����%h925>�6;;�+GGG�jc}usy�Z�FΕ�Mp��v��hl%��F3�"k�z���q�:��LW
��!z���1g�O��L�6�[0P磰i Yq��R5]�K�i�Ԕ�y���'
�X���XF/�9�a3�>������p�M�����m�N^91>����3.C�E�0Hs���ϙ����i��|��Ub��ɝ��Na�w�3v�j�8�ש���lѸӤ=��N�����ѫwz���e��dζ���K�W<�;Tߩp�7rJ�5m��>������_U�#���Q���ܷ��T�TQ흖�t�=|jKG����X&itR���t���-�w�,��QC/�Ʋy�2��j�"�}�"��%#i��.J.����-��֚�雔N�h�zZҙ�=nv�uX]����[M��FL��� �3�~���a�x��G[�dCq��>��_R�ۭ�f��I/�S����pgQ}�����Zu3<p�U��	�sA���z]����%��n.��?r����m<==(���I}���;cc~#�/��̜|�QՃ�ɓ'���1�jys�څې��o��1��|)h5�[���yylXU�D�
��jZ$�'�Q*�O�@��4u*�n�)=�/��/m�;�YR:�D�v��^�d���D�G�]�n���+w�O�ڻ��&�۬���OB����;�ı���+~yY����=����/�pUf�GYtW�������1�:uj�$;{���("F.rP�b��rP��A��(f5��ɂ�;ҟe��;�
6��PiH3f|�	�W��!\�D?��a?~b��lTm�&�g ��څPb[���^/1AUO��ؐtd���t~coY��2�}���������\_]ƿ�����H�hw)/�������?�ݨ��<�R0q�n<g�Q��-A��!�+I�]d�J�t�IV#fi��8���&��쾮�e2~�p��:fUT�C��YNC����d4ɲ,ω��v���]��V�2Y׽���g���nטT��킦�Ԟ;�Ȧ]�qoeϻ^(K�]K`�Lz*4�I�#��e5=p�~�w&YA���[x΃����(g0Y��9:��S�t�FZ ��͏ǋ�O��;v�k_�Z���oqAbw����/...߻�_�`z-I�k�W���B�0�@������fϮ�w<�9-ȭ�$7�h�=9&�(��w�^�rE��I
�y�`��*������F��O=��Ց������8��`*�O0xh�鶾�966��/<����k�Ou���O=z����ĄxJ'�#G�LMLBӚ�3�XYY��---al7�_�/��R��hj��%G~���<�gŊ�w�z�~;����� ����ۖg �L:�VU��P9�������ѹjw���*s��~�G�89d䌛���$�,�gT?S���e���!�{�q~a�}��.�69�^o_�B�����m������$$���&�('7Y�E��B� �B��*��Q���5O��ۛ��j6��b�h��(}�je�q<�����d���c)n�9�ck��9f��r������	l���6xAy{�ޭ���	l]���p�Q�ϱ鑑��h��P��+'>цxkq�W� �7֖�k�Y7[�����V��
ii	%��H��暵fNx��\ݧU����=���.�3`�(^�P4��׺2|��^��-ˎ>��N�>�h����Z�Z�:�4r$�}i>5��^�˷6�����x����8��������d���X�b$"y9P��qS����bE>H��_��~�r�����u����o{ugi����Ȼ?���e�<��5�c��Րz#�]��z���e�����vT7�̮s��]R������.�����վ��d�s�䨅;�}%�W��B�r-gz��>�A� Ȋ6,��lV���Ra�G}"��`��/�������7.^����wo޼	դ��Uo�W�vE^���t۳*�y��d��a�e������wM�S��ǚ� �DOj������j�?1�+�F��G�.�\�t��(^��=����W,���l���F���x4*E3c���X������Gݼq;V(Aii� ��\��BT�������K�?����z���컧N��M�<{�����}{��a&fg?K/����0څ�����/���ƆܭV���G ـ'DA3�^L�)Fa+
��U���:�"$�?��m@ꂊ,�F$d��Z�|j���YZw���M�a�Lt��'w0��#��x��mm�Ց�<WY��t��K:*�$�1`fg�iP�5���$R�qY�oّ��<gĎF�V��}X���N�֮�����պl�]N����m����-�4Y�.��L"���E��$^%�"+������� ��*����Bu��N>���d�� $�f=VC�BO"H]0�����)���`�yZ�/�h,J�N/�k�/�������ٱ�Q��ꍛ�.]jU���t���Ze���B�%�s-�����r)]��eR���LK�&�eW����Y�n2��z���ӕ����ϭx�~LJ HA����?s��y�/��]bvi�W#�bE����d5AX>h���Tt��<p*(�%H��T-������'݌3K��8�ꘝlٝ�U�^��ޤ��N�d�����]�f����%�zw����N���!�R�Bj�?w�3;HƬ����m�)�ւ�1�~����1�d�;���eu�ڼK3eN��:A�;��T����޿t�^�r������ɂe$��+[k7#��uׂb��Su�;��@�mU��Af�����VVt�ȁ�B��8�ϱ%GF�0��w��ٳ��ﴮ����'�����Rޮ�0,q�)Kf��@�����~�ܹs�+K�n833���CCC��w�s��ƍ�7o��/_�}�f]��6��m�V�W�����!i��������)�FCpdZ�]�n��S�
���iꩾt!]���a+pw��G]/��:���Z�l�;���=�2}�p�S�KE���~��ɉ͵�b��4�'�3��O>���#��v�+�<v�}�p��<I��$N�8�2�K�SZE����4)�D�ޏ,����@R74�L���JuM��J}ZW��\nbrrdT���� ������UW�Vr�� �:�H�P;@CJ��+��'�1j�C�R{��s�B��~3���>�j4�`�a������_�G�K[يk�v"�6i�6���ޛ�Hr�wc�G�}w�����rgH.�!��jO��l��,`@�>0��:����?��� �,�ܕv��Yΐ���9���̌�sDDFfVU�\\�S������|��s��OR{�n�j�z�y>:��z�������{wCqGY[�ΐc�vK�c�A>�H�'p	�eD�f��;�*��J�Ң����(� ɩ����!/��U��6$�M���ľ��~�$Fv����V�х�ξ��B��T�-&�6�;Ǡ��8����`}џL�ä+W�
q�D�-8?�&����]�=�kIm1�1�L�N�����g�ΦБ���X�H�s,�:�ڳ{l*վ����N�'y!�\��U�x�5�R6� zb-n"�S������]�v� �e �����3�S[�֣R����t�Jr,ݍ�2�Q�_�K=��Q`.�o������D��w���ܺ	��ڕ�?��[���Ձl��r�d1nS�;։4#�?S*y����b��-���x���!╈�"I=̲��ǚXf��Zq�m�w�ѡҠe�v��=Э5W5ڹ�p���>���RD�w�fT��Ji��B~�j�h���rv�Å6����n���N7!�)�%c�xz�'��߽�!��J�����v���[0��^���߼>?�+�E�'���Ņ�Ml�$�9K�"�.������� �|ؤ�وZ혬`;"��O8����Y�s4	u10H*7�U�-|9`Uj���6�m���l+��/�L�1�ݣ��,/��iPv^P������{���og41�w$�ǆ:��D���A�{�����(3������g�Fd�OXo������Ŕ[����,U���Rl��oÿ���Qj��a ����}�7�;����X'��َ�G<;�g>�,��#��U��6&"�5��8Y�ʩ#�q���U�հl�s��"�����T2�5Q�;� ��HXUs%"�n�j ����D^�������R��K�E�s��	�Rا@�k���J;�i����B5���-���YA��0,�~~ �<�\x$�CmϱWoJ%�xQU/��*�X[[�����=��!��s��N%Ez<#~h�]6is��$k�x�)�q/]���+�����e�������^}��n\���nm���ج��U�i�|�֒gH�KE[ p ��\�j�0�+�Z��hZX#p�ZP�-��g���`���@�Q9I��cY���`~}A��k�/,ݢ���ǀ�677�k��0J���b+�.�6�g�6���,K�5ai����0ן�'a�$[�����b�U2���9��'�6��3�&]�D��5�A���U�Vy���r0QU$^e{pSۭ�p�����$lv�d\��6Tk6�Bˮ�?�ZY���~f���J�xLĳ�F���V8͆�Њ&����%L�8��D��r���R�'��-�o��E�MC�f0ċ��L��rqi�C��{���;[���$�����\�3�h�zaY�l���M���V	7�:�"��~��>�z �`8B��M�����8��v��FUP�"N����'-����n'�w�RK���QF8��Qe�v@����(UV"�q�R;�ZU���6��{v�'���RG�J٩��K��wZb>���.�8w��֕����O�<��d�Z�MՎ�.W�䕒�Ȫ����Ña�Mȧ�F�����<�,��8��I�s�u<�z�O���V��W8����
wB�b\�v:5�����Ix|�0
��d�m����E��\�ߍ���[Ai�6A�5@B�J�ԉ�S�������_�޼��G���O?�;bb����(�������!��ý=8K])�L�y��:�ma(�C����JFy�����!�V�M�u�A��肐�@�X��sQ�a�������W�d��wo�+����Lׯ_�u��Îg=�Q���a�t�A,X��B�d�� �C���Q㚄=�`�@I�e�4���3�*H��b���1vMr�գ�>h�3P������8�(2\��L��4���ÎF����RK�ERS`����؄}�$�J�p](�]*U
� LV�g�W�d�y>� ��ǚ�����j�4�>^�)DÓ��/��
���դ,�Ú�%DQ��?��>�6��~��r情+��E�ΣkGe|&�����pj�R�T� fg��mfyy�CL^��8�}�4��9G�j@p���&*Ĕq	�...��6b�M�_�i[RV�*��Fȩ7+.f�5C[݀҂D����Ʊ���6Fc�i3.��٭��s��)4gz�T�h�@�4�f���fqoת����ː���f3��ֆZL��I�yc�i�>�IkW�I%Q�LR�ԩS������=]b�j̜U�rL��S��$��ج%Bw�(3�&�9�������}';�w}c����wp�p���᭏?z���?�r��ݻ��=��]X@�G;��Y������p6*Qfb�y�"�eD�%��l��r��+����!���<���bAM ����zI��������]h�K�l�ɣ�	�vY��[,���I�\H�s}8��� WSMV5�^�*�]��rc�8�dPOTF6($?�3<y��/�+����@�'o������U�0�Oj6�4���GR8�Y���3Qc|����i�*���/�ƋJ�t�J{��Y�
�6&W��
7�����9,��S���%�s��s!�qijދ���!�a2��hPAtF�R0�lt0�� �J�˫�k�NA}F�X�bok>7�pr8��T�� �/�[9sj7,m�������"C4Q����m�sۈ�v"@R4�hg��������V�T;%kT�D$b�aj�8q��mJD�%x�O<)�H)����[R�6���#F��TjF�tFC;ja�(�VF
����E��f���#���
�NӶ�`�E��1�u��W�^�9�F�(FG��%��8�I���~l���̼,��'_>�@Y$Nە���o��sss���Wm��}щ�`,�J�SC}�t���*d�����x�Q�xs�	���& ��T�׈��1��
�!�/b�TmˇUP��[�'_x�W�g�?��7n|��/0���n���l/5?��s�����uhhu�9fa��a�5ln��M�ߋZ.I3�zoD��o�s0&�RD�s��fQ�b�6*.�y��j.Zͧ�6�m��z�B'�B���,��R�Y>Dqi{.!�:�n��N+��
C����%#��
S
ێ�ӆ�o2<�ҷ+\}���o�
=�hY�.���s�/�NQDcZ=F�s<�-m,��T�z6���κV�70�j�pN�O�k}.��{�W��rJ6=r�P`b�C�8w��_���?K:��-
5$�*Vږ�v���O������Wkogeȇv /I�zeKߥ���92�O'Ţi�`՜N�'1��K'�z�܉8-�p����f����}��2���h4�S;�ss{�X��x	q�z�r�i����s���6�<�k�L�&�nP<�b�+p�"����[Y/G;�BQO\?�A��g���|s�>��Ѡ��#HLh� ��eZ�������k|�֔����j�
��t�����),��%����!���^!3�R��gb���O8	�=uҔ���>�u�Ȥ�����@b q�/��.��mSt;e�GX4BP��'���.�y��lg����n�z��?�����E�^O9udB1��P�jX.ȧ���ȃ�ŮC�ϭ2e4���iD%ۣ�X�Ǯ��d�{�6b���X�� ��f3I�s`���Ak!/[��ΐ��Q��0�Ǡ��x	�_�q��,W��P��F>�8ʱ���z���Y;C( ��m��G 9Χ���g��;���Ax���cϸ����N���QCқ�ʀ��᚟�ڕ��g�Њ3劘��
a�2�D�2��lЀi�p-�)��դаc>�EGI��tu�<#��)���n���I�x>�9��"��CSܻu�(rLB�y�S,�V�J��tᙓ���|gafΩMٻ{[[[��=��Ũ ٱ��}�ڵ������$�@ F�|p���[�[U�`Pj�! �y�v�8]y������t�1"�OHEѦ��e��r�������tyy�ԩ�;;{l�4�Q&�G.m�iM5G��*$FKV1�N���>��-c�b��s:�q��k]h�a{0�I�ĸ��WbL�J1��WHČ�m���某�qy	���Mϫ�3�ߟ4�Y��p�G�ye�Oa&�W�v$Ťr�ʹ���Z+3���ģ<#<��'��%�nR��F�`�'��創�`N z�N��v��巾�ۿ� �]}�+W����c� G��� �O�}TX<�b(��J��r�cz0E�&FAu6���e�1#����\bu��J	(��o���Mi�m'��c�|LO8&p�#��%
�J#Q�,�������2f�ch�����L_�Jr�~z��Xd��"�5�DPjت�y!U�feY����U�tL���\~�8��b��6�xt
p����'؍�`�#z�y������{W��/9J��I��k!�
��\igW�&>WJމ�_��t�}K:g�*J��@jҩ ����BQa�Vd�	y;`�}�Qp���0K� GMH�2@uw?��n�a2aͳ�Y���hi�����WW�Ξ?��>��Z+n�.�a=�O���puM����&�6eEPp�=�	��{|�ƽ�P�N�w��W`x�)�3N,�zA���ss��Oz'E�*�@VzQ��<88x��!|b�G>Q����V��y4���"��pXãԐG..��b����ԩS�K:�?��S��������PMD{m9�SA�/����	f���	RP�p��vP�)B5��0H
�G`c7agV�D��8n���Ν{�~��~K���έk߻w��͛7n���� ����/{ND#����$�?9\LQ�@�+zr��a ���@����Ɠ�
Id�ai�&�@99�٣���!�J|�k_<9�5)�.,���=�-��au�q��+g��@
�}�,寮䱫��^Z
��RbN�8�b���ϚBx�6����ٶ�l��vFVP���0�>���j�i1!I�pL�Ё�:�Ģ�[�mE�����:0�
��ۆ+�HL�9���0����)���H�*��@e�nS�ӆ���FK��#,릂V�MF���@1�����14F�b+��Z`��TYA�.�"I ���4mlK�t�P���FmB2Q���Z=eZ�h/f P#�����J����:-�,+D�+��=�r^�,��ڵ�w�-� ,��������^��0�8��$3)��d¤
�fE��L�cD�P�9Z�SB����ay��ő��
z�9�a��������)9���F�]�.B�ե�ճ/�_^Y��~���j���B[��E�N�~�&�������Z������\*�x��ʺ�nq,#-*�d��1.�ʙ�1&�văA����������F���g��Q�������9s�Ũ ~壘ї��b��lu{��Pp&��E6�E�!'A�(��Bg�V6P�Vu>����7F8"����%�ꋢ#֘ (92LQ�=|�-,P�Vb(:J�e������kx����OI !]�B�E锉9�Q�n�V�r��E'~�����=w~m��ߤ���L��w�����'�YX؏o�b�X^ ċ�x4�aP��j �vr@s _�%�	NaO$�tZ �v�6�7���N;I@iW�&�~��>Q�ddTKҖ�d�d,4�a� �	������wo�����ɀ�!Á���✤ĎTU ,�����ډu�|�SJb��d�5����WW��<b8��I�����m�>��p��{���v����;���q�q��!��[^Zx��A��� &���H�gi`���cE�+2�6����i��C�5��ǣ,SQ"pO`�x$bLŋ5�
��6����V�][�L��z�ȥ<wB��x
�_�V
��)J0�]X#����� T��ݠ��[�;�����|�"�/!�U�������&�Zs>.I�0��H�6�y��)�� ����!h#�xm�n����et��D��:�wF`����
�˟���x#��b\h���h���R�٘���@�݁��@�Z�_������L%؟�cK�q����2@v)R����b��w↩H]UA���1|z�j�ۑ^�+gd�/��L1jp;�����>������re���7΃�z�p�m
���C�Q�Ҟ"��-;kV�P�ﹱ��\7Z]�Q�3�r����!����bl�������3�#�O:g��|�턳F<=�g����9D�O��:��?,>���|p��/�_�~��'��gL���a�q���P	%}ta�y�N��Ji�e�p�� ��i�%� �Ǯ��դy/�O�[��R��F�Үa(zqq����msa
�a �Y����˴����r��0�pqq��ݻ�d�L����J��t�քʀ�����&���L)��o*��5��R��Ϝx��j�Ǌ*ZN�>�h�<�o@)6s(��0Nꥋ�-�2�}�c��K9������ے~��Ϯv���g�[�i����)�v5�m�͹AKw� ;U1P�Ӆ�^YZz��#l�۟��8s���O����@���4��
�fX
�R�p��2p-�ۛEݤ,F�Y������J879��.hT.�F�9B������C�oh���Ov������mo�l&�v�e3誂^3?8�̈JX&����21y!h�w�Q�3{�*#4���Ayw��'O:6���}ɨ���cd*�B0C����~,��¸ҧ[�)w����O~]1n�>9y32�U�G3�*uOe��������������@]�>��C��֭[X���a�����! �l�Y^9���v0�tJ�T�rr0���"M
����Km'i�y��O�=����1K2i�UǴ�ݵM�
��&:�2��Jg ��!Á��V5��A�[9��!���V���,-��8u���۷��?0��6\	���ۋ�d{��{��v�vA�ε����cP���� ���w��Z��j%m� �7z��-v�vI=����C��XV�j�2���U���َS�z�~F��HŞU<S
g�}�ur����|O�5ҽ�:��_W{F�C�*�a�C���|���v���&�����vr�gB��p%��/ce�z>`��vݱ��+�6r��+��\�t�N���/���6�ض�'��PPuJ<9�"q�8�� ��<�x�`�M��'*=���Z��f�9�ɊFӼ�<,�шǽh�U1��z�^�xqcccyyyuu���?�7�==h`p`KGb�;j<b�%x�f\d�X>�o<5!�|v�|�e�S�'^�_)��	(�v�\�R�g7��R�&7<��Ǩ�`������gg?��	����⳵�cl�ɟ�j��/�B��� �-$��c����8{v��y�sp������������{����O>lo�I@��9a��!v���f��:�4)4Ai[������A��&������Ay�4o��țMog�B��������;���=}�����v��Ū��S�lkk�8
�l����ZI6�'k�w-r8��p`��n�)d����t���G���øh�ڻ�����UA9 ����g#�����"/;p��W�wOܾ&N0��ßV9`ჩ�)�^�����[w�$U.q2|&��h&�Zh�L M�����8���y�k�s�ܜi�6ˆ4U#?�l%3JG.U�CO����]Y`O�$B�����؂}i�����3�V�C����X�pd�R)a���U)@�+����sQ�bfI�\P�;�b%P>��A�!fm&�Z֭N۷i������J���ϟ?s��ٳgA7=��#U���Rي%u����\Y��¿�y�K�x��!E�9�
ޑ�ݖP�y�9G���I9�C��%ޱu�tFN��x�vp� B������S��:X5����H�%!���U�d
��$�K�]mz>�D�
���0j#^��I�_��w���9��ZfG�8�Y�:��_��&�L�����<sK=��~��o�@���>}�ѕ+W�_�������[Z.���i��T�b�U� �`}�t!a�6Q��M�oZ��<�5 ��^˩Ņ�#��+��/Z����׮D�`��2A86�[h�0��i%���pqqyu���s�V�Vo�}���w�Ó�s�'���م��@��}�Wϟ?���?�=���5q	��Sd�3z����X."/�t�i]n�2��m,#�̴�ا6�B+Zs%pi�k����Kc5����c}_!��C��Ϛh�3���s�B$y�tيQxtU�C!��r�7��C���n��� �ڳ�[/�r�<^ �E�n]��l�j�A�����zJ
�5��&	`��j|�����z���Aq�)Z+Q�48�����]��F2�uQÃ�}��eDp�.vm{�R[\\#�<����= �{�Iը�6E�h��կ}���_}�G���7o޼v��c����b�Snl)m�b�n\�ې�����m���� ����g�o� �S�C>y����N�c���hF�\+1$e1cn] ���s��k����*���I��>mt8mQo�n{�3 8��ֳ��c�W�XAm��n7m�������-<��{�@�}p�W�^�y�:ඇ�k���{ �u^`*�K�Z����FXm��z��
WZ�J���uVR%\I��൱��~�4h����p#��z�ҥ��΋�H��]��q���N.&X����g�sk�'p&�i��RBO�S��Y�&�9�����y���J_��4)/�m����aJc��i;���n�쨑����Wd�R�������,Y3��pR�J+�,��ëxt�_� 1#���0��u߿��������\�g.�5Q�[�|�Q��P�K�H��k4�r�b��[`
$����d����#RDDs��[1K���0��P�� �%8ใ|4v���+��-�.�p柊_����
��8�^(; �5�������'N���+gΝ�ˁZ�YZY�s�΍[7oݺa74����{sİ���5l%#"�.W��HR>��Hj����lf�լ�y������g�ûX]]eǊ	悘ї�j�� X튠ބ�b�m�~66�M�#m���T�����{���y�':}��o�{V��=
%���:9��R���:Y�c������S`vj,��;�2N���W_~�mPF�V{o{��?�q��O��n�yp��H�6�ȥ�Ȅz�ʰ뉃WٲI|���bW���@c�������AAk壔�?X�[#w�A�L�;��������
s�jÿo��w۝N6̒v'/rP���A'iL�>¦?�����?�߹�iF=�$ǎ�*�����+x�B��E<�Xw)ƛ>1��:4�*/���5�U�`4��< L�w��ݝ��{�M@B���Y�Ĝ��)x��
,^F
YE0���Ԡg���/K��C(�cm���&�J�Y����ҕ!�k�LWm$~���j�<����Y�Wk~n�W��H�td[������Nr8{B3E����8��M�XM�8��E��������[�|t��ƬF�̟"бx��%�^w�3�K�����f*M`�'O�>CURc�:P�`l�������>��Mw�+j���K�zQ��|K�|���P���ЈE>+�Dx���z�t��}�����̺3���vXIˌa��?�d�S!�O�q*ɠ��2.��Fk��`aH��5K��#i�-A!(Q�� !����$R��(gq�ks�}���_��_K�]��w���kW13�����/~1:8��M���ީlĿ�	��Y�4/�5.����Bwanyy���j��]�֧O�nc
h�:����q�p����"����������S�/���J����²&$uZ�JQ�"�̸J�JRQ�m����+z�����5��IW�ۺ�+���5���6-F��+X�ZRf�3��6�b�_�q����|��,��	᎗S���w�sv��j�>���]�W�Se�F�WV4��"���P�JJ�w~q�!��į�&�s�d��LX
�$�F�hzn����ґ�Az Fz�pʑ��Ҙ��M���Fƌ���L$��BDVC��D�������5��@C�rۃ��֖��Z؞v�_�I�á�M�Ƙ���U�N��N��W_mu;;;;��.,,�ٮ~���~���|�?8 y �?D�~�u
V�:���"��p��(��i���^^�1&�F����A�o�2+�J�B�
El<Fΐ���)���c%�� 0�`p�7���/�-+�i�?V��xF_DjB+��װ��?8��/nżZ�O��t8�,��2l�8j��}B�4�*�ݩ��b,��Q+0�W��z4R��#e=��1Y���+hUnQB�ʕ���A�;�$Ʀ2�c�(V1�\*�	�Vǭ�}SdK{�NW�����_z��]T�m���j?�ɏ��֍�A6f�=]҆�;Tҡ*k��e)�GC�Qi���&�1u$A��B�����A�<�7%5���9���\�swc]�v���X����a�[Zx���'�U�(�&T~5�s1?��e�󌞉�����_�����?�i18��X�u��.��(�{*rAզ��(o9+_�-4Qf�0�GB���xv��S�7�yJ��`�P��W���B�+��.R�sL7����'U��lA� [�q9͚c�eQ��MxM��k;�P(��U�:o��l��ɏ~{��G�%�A}�H������t?�+ŠǼ���1KY������G�(p##s���_~�#���;�Ñ����k�Rp�͢lC9�� ;��⋬c�F[�'8�=��\�'�cx��M�r�'�3@{�|�ɭ[��}��۷o�<��vw��p�H�N���ޡ��tr=0�W6e9�>Mi=�Uu- ���7|D��]�
�v�[���F�⌾|��&6���s��.��b�e�K P�`2���b�FN�
�5�ξ@tL���1N��W�������_�5�Y>ڻw�S����{�}�� ѭ�e�[C����x���-��"k���Vpb�~8����7��a���8��{�Fݘ=*XՅ�)6<s����/c�	`"�Ͽ����g�ԇ���E+� ���(�I�{��{��xje	.����F^9�?4F8c�{z��,�2v���O^��4�c�AY��8J���<����!��;`����A��� ���l�U6͔�1D	��� rsd�����yw�dm���t�=\�֔o��]ڕ�PX������r���s��J���ؘ"4Z;%E�7<ߨ�x�Ȳ �
/ø�)e���q�e"�ŋuX+�
.�Kj�糖0R;��;�ԊϪ�� �:�QI��
��w�������PsQEub��>�j��h)� �g�{ai�;���0Z���C��A���yxx��'�hk{c&|��Qᣣ�KPQe?iu][E3yB�M�J.ۣ� Zc�=��6��ؙ���HS��(_���F_�퍦I+=yj���#t	���*f���K��1����3<qu��4�"�z���ec�J�3����<r�	�y��pD|o�����3��?�"����:I�/t%�L\3Q%�'�_�_���m��z� ��\}����_�z�Ν����Q�����"f+5�[9�&�����5D"��2�A���tZ(��to����Erimu}}}ni�^�����/^|��W^Y9yf4��[>�B4���&m���~�;������'��ùN�_X �ocu���=�"�����G�����P�N?}��Fy}����[<� O#���<3�ĕ]�Ļ��3i���gay�gf<{K�W�}�+�ד�:��G:x��/����c8h�Y��7�\�>�v�$lX����D5��n�v�>a����I]{tR��{6��~7��,���c�gsS��.�D�.����Ế��Z�sT���n�������~M��`RJ��!]��� �6.���A4l�`���p�|6���D�N�n���Y��v�xΥ8�
� ����F$�W*�mQ_�{�G��Z}��Sɲ?�)C_oD�ڦH;ND���ҜGO�<��A~�۲�Π�����m��F���N,8D�����!�Kw�1o��ɥ�p�nQ2�C����|F����KK/^����m1n޻w���������}�ѵ��):�[���&m4E�E�����}؈�1G�^����@n�9�4�Z�9??��[b�#���W_;}�6M[Ơ;�F��B�H��$���/�G���w�kS.��I;<���{+7�g�uj�G��Z����Y�Cm�<�/��KFϰ3�m7޿I{(6����� d�c��(�e�v{9XX �D9&��Q891pyr��rqe�څnm 5�Ү�����4|\��8�u��
�We�W�D��J&�V2�3�y�%�0|���D�������$S�����9N�pW�f{�R%��R�ec�L��kɚ{���B^������,�0���ט����P�aB�7�Ept��k��Y�Ҵ;=��^L`�J@�� �ǭN/�2��|�ԹO��|S���T�RNfQ���_]QD��#L:U�(��1a!���a�8�9�lxn�vǘ��s���X�����!Q���5̱qf~e�XS�8��d
k�r0h��O|��i�M�Q�S�+��\�����:�1VOO���\��%��u��I
�#��o�Kg{Kg`��~[��p���;w�|r��իW�\y��͛z4�.�E�!�\ ���<u��4��ٙ3g`���>����u:i{��݃lni!n�]~����+k(�st_J��g�yԇD�3[]\�w��+���7���ɥ��|�m�d�����Y*��U��r�L�J��|�=]�a�D�.�Nb����7H��ԵC�2��]%..6�6D<��\�dW�B?�	a}qrdх�!���	+���"����>JU2:�/�$�xB|v���;��]kC���J�)���&���C#��R�6c�,��-�Ea� {v �+J{�c�I��z��[(�ⱇ�}'�A�E5�
Ł{���6��ڢw9#�~����TGf/�� ]�ÍÔ����"��� ��Y�*<+��G�	��p��$'����"x�4n�K���bx'���
�X����gu���^k��^�g��6���!��r�!��T���y2����]m^Q�\1#�����`�G"劀
2AIi�y�wX���Hcl�(2�j-�<���z��W�+].��kW?���k׮V���������	�>}���n�{�ҥ��=�'(���c�$���]X9��;�̯��8�(/�$nGCF`"��p��--�p�-����� �7���B�W�dq�x�� @��z�@:k�	K�Gz#���zQ M~��da�b�h�-�$z�4��P����"�'Ϥ��G�:�H���&�m��~�y���g!]��Є�;�K���0Ƌ�c�=׿Ϗ���^��L8����Ҧ@kO@x�sZ))lG�8�]Q��$���5
gf)�nV�Lsf��1�8<�R��Y�O��w�1�(�f0q��>ԯI����{E�%�'��&0���P�$iIJMOZ�0�U�qW�N�x�M���sO��L�����K�
��K����_{<
�|�q��#m� ��:Ϯ�!cP�u�c�ʄe��-��3�J��[Č��*o���Տ�g�l䷚h�-l|Bp!>���K�Q`*<�
Ʃd^VK���WT��l�CYq�:Ʃ���7�qz��*�>�'���{3�|R�	��	����]E��)JG�#�"�(q�/�����o�ͼc�J���{��ݹsggg���;[[[X��R�k'F��6����>��~����dn1?<�1����n�=�D���őe�>�1e��%	8�_��o�����?��/, |�,�D�2�̯��:(CX�V}�Z����+��/��rJM��4n=�*&�T�E�9���Q6�ұ�Ϊ�~�'Y��OMX-�xsH��Y"��;�%���C.-���չ� ���S�jh���g���uZ7��U`�6�����x��#rV�I�����NNu��v]�5���>.��l��S�3Q��"����ռ��8�q����?����F�hwFxE����@0�Kz��3��{��q0��m	����̵�[#�6��j
�8�Reh���cA�&6�ˉ�ǷRWX�:�;�Gc#)�JS�����������e��lT�qL4E{�����c�,�
s��ߚLTy�3�������L��Fi�r�5��y �rS"Zi�y3Ǡ~M`����J6����$���QԞ�?��=w�S��n���� �Fc'�����e�sn��/�w1�L�����*��B�B4���B�&���G�ӏ~��w���1�Eg\������^��\�+h�c�
���L5�_B~�3���:4�v*ƕ>�.�:��`Ҧ���s��r��B��_�m��晦�u��6�r-�^�y�w<�	Y-%Z���Ȕsr�{�� �c�dɦ>C�+"�HF.ƀ��X[�?;�%:4�����C(��`o�bD$�.ޝ^�Y����QLX�8,(!��.����ʳҞ%}�E�}���ӑ��W�����\.�`���~�m~��'�Ag���A�c�׏�#����Q4vk�.a�<���I��c�͛7YS)Jd�p�]�G6�@�5F�h���U�YG ф��<�$��ߦ�
�!��͟2r)��N|-��;ˬ��X��ͮ�llp�fĻX����u׮����&� �k�K��Ղ�4'�s(uOA�@�ޜ����r��w<_��f�{�Z�[����p�F�����dY������P�*��B�+K��F���^X5���ǹ��;�<��G~;m��� �$J�,N*��X�͝8�&��b��ҙ"m�?�H+��1�*��o2�R�o����o�����g��\�װ5�H��bM��jgb�$BT��R�S��DEI�HD�U�HQ��Uf�B�a�
V��B�Y�K�|��f��p�Xr*�ˈ)>]N� b4
&$_��r�m��'a��e��T��,��	\$~�NQ�&�[�a�<��_���m��6� ��ٶ\��'r�����$��}�;?����~%-�]%V���.j(	/��ō�gBT�ϤG'[�?>�g���wkL����"n��k"��v]����c�~7i�%DՅ�R��9��!����d�����oN�z嚴UN��_$����У���.̭����@+��	{bsԞO���ʐ8� ���J�33z>)\l¯�N�B�P�ؓ<��K�c�ӝX�rZ���{番��sHM�/?�я��/�byi���y��ƣl:!+��.Q��E��D�Um$\��U�g3�Z�5�*�i+G�w� �So���jC�cU������Ʌ�#���"�H���5�Ҏ�Xr� w{ݹ���ӧO|�[����wDQX�_�-,*�nZla�~�'�
�EJq�-�<�ċXΦ�oН��O�� _�/O[���QE�q���vgwan�ϲ�����
��������X��/T wz�n�S�[s��7^>e��Q^�Y�8�Z�6Z����� �3�>Y*&O�:��n�B<2B��_U@�����he;uꔒ廛��IZ۩�!��V��8>O��i<;6;��I�KR����̚�$������e��8jk]���w~������1��K�;;;��'܀>fCLj]g%P�ˎ�/��B#T��͛��ֈ黝������E��T2����n>?er����[F�W�L��<-���N���/�/]n㳊u��,�6'��IͲ,y�$\h��7�|Sp�K�S�U���/f�>u`d�zͰ��5{R�~}\H͛�8 �vb?Ț-bm#�"�[*����Ju�23E�8H>C�R�o<��p8���k�w���W�$�-v���x?cp�@�*[&�aE��A�*5l��O��O�<�s�����'�w��sN��dp��@��kB�P�ɬ��Yڸ``�<>��@F��R"��e囃y:(cF_(�u���E��;����K��N���Wn�UI����=�nKX�@6�Z�$���:��9K�����ILL������ �u�)��Q��|�5�G���&�e�|�`��,wJ{��(��44����ݵ�����~��K_��M&����"�-���#�֜�V�{$��^9yy-~���c��{6=iS��Л��zÝǾo��h�q�dmŸ�嘃��'vrٞ����^��eY�e7�1ϸk$[�lp���C�Y�|�����`��uۜB.o��.��7�<T�߆ZzccTI��P֛F�YMѦ���cWUApK�g��@v:�V�����3�	����v���'�j�|	�i�LJ�')Z�Ə�'��<}ឤ
��V�v��~�;�v�ʕݝ���ui
�ou;F`��`�����j��s�3Tf��+ϒU1>f<�_Bҏ��`���B4v���u��%
(��~Ɗ3tFbjA��Q����Q��,�j��J�XK#P	��Q�-^�m �o���[o����5�F���qV%�4�����7�=��;�:�CM����շ�����6wh�O�Qp$`>| 6K(Ȗw<����8�H��/�}�=O�u��樚<Q�vR�#J/��z�Ƨ��U޵�Ĥ��$9�N�'�p�
k	�g9s��FȬ�5���3z�$ɢ �����r���)����/ܳ�(y�e%�]��/��4�"�߁1~�w�/��/[)vs�����l��n�]� 5����\'�*ׯ�B�*&m���K|�H��1����3{�KٴU?nt�9v�28�- �Wg���pB�+.1`TT`Ҧ�v�������]�p�W��w ��ڽ�O�
�(�^.\�ޤ�'�$0���x���ߐ���O9�»]�ug�Q��i͋L*�*'��1�	Q;!*5��Xz!���X��Հ܄C=����C8��!�KLuG�nab&V�͉st��'T����EqBI6c]�yEݹj�)8UY�H�(JaU{�@��*�*���<��9lQB:d�Q`��`��j�c�})��\/&X#�t�~Ǯ����kr��dt�:o���k�^~��kW�ϲ�ݡ6PE��h�R��I_v�a���
�A �~	�-����X���e�Y��z<a8(��N$���QqAL�R!�?�"�?cq_���F�����$nbmP ��!�����sss�W^��v姧�M-�)��K*a~<�q���V�D	j������4���}#�q�L����}�����T��'���g3jem׊j
G՞ؤ�J�گ<U�7���<#��)����nq,��Gc��Y�٨QZ�����3�������sC��i��[��,T!��]�$v�i��V�x0T�>�J�ԅ3	�|�������"0����������������2ԋ�Ki`9�(�T�T�d���Ew�����I@�[��yj_Ą!4�q橯�<v��Oi���T~���qu���y�L�����B���i�#����* ��<*Vڶc�����\M�V�e����M.��<3C,k��R�È)�P�8I;?|�[_{�U��y���]��(�'�rs�K�җ ��=�ʟ�A��hҟ��I���/U9������3��qO;�b��S�E���i�r̷#�{�=�!���խV;��8�����U�je�z��zi#uDhl�u��9���8K4�e��c�3�B���F�"Zre,�#
����̀C�x�� �_��:W,��';�/%UW�'�U�RZ�PGa
���c��V��IO�7��B�;ۺ.&X���#�K��Ѭ�Q�F��E���g�\���LFK��W ����<��������.-.����O?�ta����E����$��Lm�/��ݲ�cض����J�He9��)�`SR��`R4+v������l�5�3���Tz"q^D�f�����Q>a��pO�~_X.'�������|��_����.]3{�6�Y��3&��N�H�����-ώI��4�`*�w�%����N�e�y&G����9N,�13}bF��k��Dd.�Q�/������q���u��ɻwnq_���7B�qh?cL2�M#ܑ����{�3�5f��1���0ha�,������I{��gWNŞ]�hpU�*�.���،㺀�F{Z�?�Kx�����/^<����YV�3�V�p<�u�т��9��.�߿4�4���x�o̳��p����)��r�\G�I�9�z�$�M�j�}�hNj\oD�(����U��ˮV��bV�๦��:I��A9�p;�2{��u!�R����)�Dc�ax7��/4j�f�\�\[@m�=���^��?���bg{����2'o�3_5{t��+3V��,aɹ�F�����u{ѩ(�[gk���(ó���7C|6��&%+�����rc�#�_�g�M�>�D�܊����R,�FC�ѻ|��3g �8Ӛz񺲨\k�ug6�/U̫��&7��H�K<��Z���6��(����,^k�8��y#��lN(�pH-�ef�-C��Z�[*��g3D6��
�~�\���$��o����wA v:������c�t�T?�<�4�������c�a�nq=5>�6�>B5 �9�2�.��	�Vy�Q��P	�l�)%�o7FǪ�a�$I�����;����/-..r�7�(46���s5��~�#F?<���c�N>�3_MmYM������fn�O^	�]�l����1ɲ!�z!�Ϛ�����Q�,�È�Z��������%ŕ���̊�ܒ�({��v1z:�Az�k8
�0ӌ�ƒ��x���ܦ@NIA�Zr�u2�l��=�D�RB��������o���?��?����ϖO.p!.��_O�������Q�?@�����RY���DE��	��Xn��#�y�
��p��=�p˔���߉��5�$?iy�n#����'N�������ɖ�!�o.f�e'd?s��%�y:nuo�}v�V�!Ï�[ ����`��9&6R%�}l�i�w����/��g<u2��Ōf�(�9�;ְ�c*�!�|�͟��g��^�x2��>c���w��4	�neom�I�e��k@�����،��E�a3w1�z�*�*��q�8	.���n���!���0�6V<*��`�����_[;�֛o����2�6�e*/rƶZ�����k�{,�r���gm�_*�u�MW:G��
���s?�n����p���{�V���U���o��AT����<�ql�{x�/��ѣ�#V*�Zxm%�H����S��ٳdu=��ɪ��iu����dd|MA����kk�]~�ߨ��p���%v��,AR5�lµ�A���g���е�JEr٨O��My拁�/)�<_Z3K4�N�6�&���E�IY󃥋+h_�t�W_=�����k'd�&��gjۗ�*�y�Sy��C�S�O2e&Q���xL����U�*�۫�5f�\�&l�G�Xf%�g�$��R�T-/�����������h4⮏R�R}��8��yʙEC�O�r�>5��n�8�eX�PH�gHz�6\ⶐҏ8���Yѣ���2�ݷ��(���}!�����с�b�(şE&R�c�ć&���@I2#�Ѐ�;�n�e�Q������s�͝W^y���F�a����\�e�e�.\����������N�~�4)��ĘL�A��:��a�����sI��4!SF7Ox-Y���5��h.tVF�X��d��!��<����|��Q)�M�+����l*�����z1g�FԊ,��dw���X-D3�W�⛭߼�yF_Hj$x�^���a����U-T;��b�Ǌz�bƺ�(�l����"���_�|<%��
��S�¢8W���(�,7I*T4�rym]���"k}�f���Q��3�b�n�A?M��ƥ�կ�[�7�P+���4M���nD�5�� ,`�KalM@�{))�+잮I��H2����V|��}��.ް�0��Q�#?+�i��KG �#]lmdi�`��$�&�1�G�$I�e���q���<���H����l�K�gxC}�Y���TF����O?���ŋo���p8���QnŏV	bF_22>�̗��:2��J�X��Q�r���t�#�3y%(ǙǸ:�$���8�1}>���R�)������D T �\�p�ڵk^�E��gg9ʩ�һ�Ĭ�b�|	��1O�/!]vc3�+A�8v�EaB�Q��8�с����:����1�;��.��6�:�s]�irxx�N jy���s�-��onl�����3�;��<�8���#��*P>N����Ag�㐜8��X�D�vU`9-[�������($�8X9�1�C9�#��!vQ��Ou���˪�ь�K����8�կ^�ŕ��(�R���P�C�ݲ	�Xo�����X��lg��V�f�1d\�Vo9s�<ϗ�p�����cA)�� ��ki*E�>�GWe�ì#A���[�VT��?)z,�rV����9��o���ٳg[D��>�$3zΉV0fu����]�?t7i�f�״(C3�4��t:\�gF3�$ڣ��	Ŵ$2SmJ�LQ���t���fϴ�IUX�_�)'i�/��"��\f���T������fߗ��E�O k�ǫ�H紵W�E_��v�P��tH�(X��y�0=�&�{N�s��;�0(k�R�����Mv#>ǟe�����S�k��淕J�\�Z�"���*��M?��'.S�Z-�Ct1>OEV�WD�������Ƃ݄p5�lٚF0��`@
�����«(�s���3sͨF��{`�ǂ�E7�]���wc,׉����c���\���Up�d��<j3:�|"є�����o��?�#CŒ��d㮅��rGq͉��[�|踝C29����+�?�H�S"@z"C��ߠG8���o�nw�Mhy�aLi���՘�����mB����0�XL���Tq�����a�$��k/�����R�gQ�
W�C�P�Ոzn	����5���&O�RU�t�_�>������g�gV���U�͚ь���@�h�q�ɫ!��Y4�������8��A�˗/_�re��T�ke��.�=��M�����t_2��S�9dۓ7�ِ�n�E[<W9�.�C闌4���i�:�J��qp��v�=l�ܒ� 3s�]��"
Qd��E��F����_9w�<���Ĕ<�W����ۨ��!@{`��b�<\�1�C�-p�O|��R������c"L��Ҵ���*��-o3jR��B���1	^���)���/��֙�mOu���gGv�h�g��f�Ȅ�y��8�>1!���o\~����o�GMI��_�����t�]Q@�L�b`]��t>r��`-��1Zd��k�?�õ��
���H.�J�W*{$2�;3ը2?ĊS�=�m=�z�����~��̙�/v�=xi��3*���i�����_g����l������a�Ii>:������
܎l��m��Q��i����� M��u$��#,�"bYc�x��g�T���o�'�-Ufrw�'t�x1nl������&8c�����SyaZ��(纯�FF:�[��v����&;���I-�
*�Dk��J;��9��V߳,�����Gy��w�o�}��L�.9S�@N��V�8{~�T��b���C�������fesQD?����3�i]�N�,GMdu�9�xS�U�`��z�D�29I��Qe�&1�hqq�����h�0�犜�FӂӮ1oJR�%'u˪I�a:�~q�h���J8S�u���� ��i.i �V�E]e�ͨ$�(���Y���P��}������oݺ�կ�x��mEܕgC��V6쎐�%y�-W� #�	򀆞��6�*�0<h,@X��t�Ҿ G��\\Vv򠙌o8�piX x��&���+��T��2�~�?j�ϟ`�`7H�>|�����7�vN�>}���ac<�s6��TM��q���֘J�LO��B��U���>����$V>KN�8���R6�I�K剆��)䟧�(�����S�+h���2f���1�c��d�п�n �p���O��={���뫫�;[� *�q�d����U��汚�'�g�8Jۭ.UW:4�ץ"�s�I�F��땸��&������?lbZ�"���/J��%"JP�gI�e�Pəs�_���b�|���g�}F�F�O�∌��dUU�F��4�4�3�+Fz�3�&.8����	���6���h&m*Y[=�[�ڌd*�z=�g�e�j�(�#��l�e��L�UN�82�dh��$�ɘ!(�RPiwc&9Uf����G����c1�Q��ο�����...�Z��v�&(�#���{%IY[�̘)� �l�&�nM��eh_�<c���;c���>�U�_�`�&��ӓ;h+�g�3$n��!�D�V\�������/�t�ܹs�]T��3��'Ϸ�Q	�+��1�$�Í����q����F2��ט_м����t�ۻ�.z��BE3����S�������cص殉_]�?�y��:T�>K�l����1��an����j�_y啿�����?^[[����ypp z�X�RƓ]=�8"3�f���vc�6�FS�B��� m�\�͌9K}��V��CO-Y���@�kU����oͱS>�(r=s����zY��������oa-uՒ��
��e�̄s��y��tDv��EdV�����9]	��\Q]��;�*�T��.W�3M��h?I[j��<y*JZQ�f��fT#ǸQ�7�W\�4�\�������/�K��e�*'}1�I3�Fx3�`[��&H]�E��ٌ���#�Ų.E�V�s��7���juu��$���8�l<�<Ja��v4�huN�IKIeA���'pn
���Pu��� (�r�t��a��cդx��frS��9}Q�Z- j�����v���ˀ�)�U�SQK�V�����B��h8����4=��Մ3�7Y�vHE��t�4�%�����<�3|6�I����0��j5�wo�҄��.:v֌�Ӹ/hۋ�3��ٌ�KJ*��h;�����o�����;w�����!@%q�yφ���xښ�>\2¥�#�K|f�)5??����%���jg��t��Ƞ�E�r&��yӬ���u2S�c56{������ݹ���_~���e{9�9I��Ì��4e�!��QnJFW2
�]�p~�5O���N�^lh�0�x4ں�e�2�3[�pyy4��2J�87c�U	�;I�o���)X�Rr�Χ�;E-$�9�HH1vW^ap����xQo\1��(���,��*��ͩ���׿������F#�ָ3�S��ѓ�am֌�a�U��&�^N�XO�D��*�猺&�h��,�:ǿz�e��*ˏ���6<���A�ۅ�|������.]��I^�8�����"�Q��3UlF%�FܘpQ��R3�����n3��	%��D���X�=E�91fd�4�Hȋ?��Q�����]'�a?>C���Ƴ���<=�O�&�a����QI�DX�!�\�h �����g7n�hQ�3����g�,�yJ3-��"]}Z�齙���!��C�a�*Q�(NWN���ٺ{�f�����'p����`0�	�3t�����pX'STզ<�Ѡ�����*?�N�a$+,H��Ep��5�E��A�i-�x3����K_}{�wB�ֹI���{��V�����|Qm�p�2������zKi�b[�l8B�{md�d�Gvp[���zҪ�:�[�3�2�jgB���C���w��H28�<QRdE+nEq��s���ӛ7�pn��կ^�+�a��PJ����3j��i�@��y���W�O�*��bB����D%��4Irb7Q��a�>��c�p����1��,��Qc��D��[��A��aRi��)�+�bey]���.�h�x{F�U�]Yѭ_r�S�Q��v���wn�d�>����~��*r�p;��(�
�~F8;l�M�6�ʯ��kA�ָ� �T�Y2o6���.u"B�Z�,10��hĠ#2#ed��ӄ�	[��-��^ouu��իWϝ=���۷a������O�t8�k������i�S��A%.Wx�8����m��4M%���0y~~���u�"~f�g3j��(HjP_������� Ԑ�\�ES��8V�
�ĥ��NѮ�s�0����e"0��S@RA�(f�G�7�[v�a��^~&���a����YI�5����n߾͝`8x7�2�eT��闢��C�ǷWl>#�x�34��dl�����6��3ڌ�����9s��~�n=�0�f}���q�e�T*�ٸ�d��\�c4��ض��z�f$Hx���-ᒡ�f��ӧ��7�������4������&Nf���F�'/1�����p7׫ ��g�.�+�*���9 ��vw�E�֧Ϟpv��)Bf�Uѫ�ь�c|�Bn��`�GI����P�ѹ��_[�O�0����͜��Wi����Y��,�`�2���E�Lm�bd�Xs��(B���fpp�gzyi����5��b�.rV_cFUR�?��6Μ=yjc��@�<�z�9�?�;�\6���F5�]
s9�~�pI���n������
y[ٚ���+���f�ƌ��K��.]z�?�8J�o:�:�� ���GZ�X���MS��4"�C�ѧ
�<U�`��
��s��h9����鐾-���#��r�Ka�
S�/-��ꫠ���?����v���v�����x���������{�O3�0~��3��	�&�(m�V U����<yF�����Q��x#<�"fmFy��o�p�B��`sssqa6����$�%фk���Xά�L�Z������(�q���J��>Sw4�a�N�������.^���ƴa�0�d4k�3�&a�aҿA�}�W���v�T�� ����l��H+4�����S���n����Ǎ�5-(�,�����f��B�/���K/���vZ�(��$��?��X���C��Rex�c��q�q���	�w�NB;[��e�7�t�|��'?�	h]����-����]= *�[��0̀�hc�����K�h�F���3�a����`�ܹ������,��82TvZ��m�M����яt��0C����.�\��ۃ�â���$�	���Yb��F����KGٹl��F��������)N
PJR'�q���;�Ϟ[Y?�g�2Z�$/�4�f4�ȫ��!�ƙ3� ����(�s�6+49H��>B?�p��]EU�cf�7�F��5���Zl��̇�	�'�|���q�&��´{s����ݻ�v��֍�#r��r����o㈿jSډ˹@���x ,��(�{�9$�1�h�܏�}�X�;�����a���I���B���. ����GV�o߾�_q^E�mX^.{V��[�'���8Av�B�V�@_j����������//--�U,r#&��(�Zp O���X�������8���W�O�9�%~�&si�菦je3fd���\�jeu�Ib�+�NX�om�ԩS�k����ғQG�/�O�&3�瑌m��)�&�{�嗁�� H�c\ta9��q�%����B3���L1<�&r��%I�p~���gڎ��>���		X�(��@l�?����)�[��R���ʂ�`j�r&�%��@E�����Vb��c�i�T�7�>\�5�Slp�eqn�%?c+4��S�ux�*�����7�b\�`p��u�h�����He�Ma��!JC=��Ϝ�Nzw���| Vhu[hKP�?^]9���]��(-Ҵ�f|x���3��$
�Y�d���/�<}��������9�t�9<������I��41.��_ZN?�vf��1�J�P�Ley/m�{���'7Nch�Ū,�Fr��f��v���.����;��We$oܸq0<d�916��(��g֊�%��o�jv�apHKi�(bc-�v�6�����>Ć�4�������PE�m�4����	�ɋ����nd������)�A}P�j�,eoH���u"���z���a�}#�v� KC%ӄl�>歪l>օ��d�c3C*���깶C�[%|F�&�y	�g�=�l����x|{s��9�"��T��
d4MHAJ��צ���8��M��_�\�V�3U�c��c`G��}��L3�`L�O|�ZaA�����/5�8�!}�	SEx���ņ}c�؍�i��b=�ׯ����S�$��]���Y��ѵ��\~���
?�}6�s(M�0����bq?�Lì.�FՃ8f&5'BsKϼ��~�a��.�p��r6ˣ���ؒ�>`��)]��س·Z��J���I�+�tv/k����`t������x�B8�k��j���j��??�0S�B����²���h܉�g�X?T���&��h�hv�4<�t)%SL`��L�4a�� C&�4��� ��W��ѳ,    IEND�B`�PK
     uK\�����a  �a  /   images/9aa3d03b-0c22-4f62-98c6-f5f844a0dc7c.png�PNG

   IHDR   c   �   2@   	pHYs     ��  a9IDATx���w�\Ց>zc��鞜%��(�P� D"�`l��k�6�q����L\��$�d��H�3�yF���=����:�����޺��QO���ԩ��p��Z��r$�v,����i�_�2M����\&!Ɋ����iӬ����5�;Nt�>�1K�";re����qҿ���v����L��K���a����ޒM�7���L����[:��I%ҩ�#+���r�4��KIA��e��b۶")Xe�_��d��Ā��Vޔ%�Pٲ�e�&�%;���wu�WU��Ko�+��(ֿd�l��j�'\�q)����|���5�N���"��!MV$���ht/�(^�����
��p�_1%���H$ ����\U%�86�ߑs���@�#��NQUնLh.d)��`u`�e��E߲I��c���_�t�4l�0���@<�Lɚ����ID<xh�F��8�"l0֏1$�U5��P��αUőm��!�%��!9|g��#֖A����m�o|ͶIai�
\�ߪ�� I6M@��b}-��k�\ZݐM���|WOwG{����WVe�W�6c������\6�7|]U��i�L�eR���`|0���K��J�Р%�R�o�1�\O_w>�f���R^^..�������vu�����R�T�,��~�&AAo-GH�e�� =��~��"��l�����B��K�A�9^[W]����wu�?|,A�M��z(Z^**��sy5p�p���F��x��f3�߷c�@,f�MT�45Ea��A���5"�pl�-k��4�2���h�Ħ���=u�ı�'�F���z���P|Ҥf,��P����Ś7x���l�G҂a?]-�������_�SX'ȝ�Y,�,��:�y���c{����� ]5ms�D���HD����岎���%�J������4y҉���P_Uu��k�.�֫�g��J����d2J��i+�-)����;ؙ7|>����av��⎎S�'��6G�7bTuGW����"�Q�.+)-)	�|>
VD�:tu��}ኊj藢��-�l"9� ,�W*�:��V\T�ןh���@UH��Y����駇���\���G���a �ܞ�[��dmu�铭v��T�踝b>�<��z&i*�;Ijp(9��(��w��b3`#���!������	��y��xl@ .e���ds�%Y��	���(���eLq
(:�j�O�:=c����.�?�,,��2�D� ����O��.ހ���j�������0L�V_S�DG�e3:���[[:[[F��/
GR�4� =��bBL�	
��i*��*
,v(�Ǜ&��<��ٷs��Y�PQ4
]M�v__߁={�!�myiyey�`��d��%3ob�����Hq���Ϡ����y����X��b��,�@�u��!��v&��x�����~�*�3IX�*�Ƚ�lF�'UYs4�ș���(�DF؊�g�>I�B�����8��� ߜ�K�R�P�%�F*�Bݽ�`Rf� <���<T�a�F��:>�Ov�T*=0�����D(XT\\�ϡh�P<��ǡ��d:-I��G��nk���y�Ys��1�,����,)�e�zKkKζm흭�;2@2��O��aIl���;�C�ϴ �XT#kx=zCe�ı��Վe��Ū��D&�,` �W���cF6�F�4����M�'�B��}x�̅�ah�h�8R�H�	�I�h�b�`lU��Id�ʹ���2�<�=k���p8Z-���_|`7SًW���,��؍�����*+`�
{�<�ħ" "��Yd���;��:p0��R&4�ݫ�BAoކ��
�}^▒9�=f?��{�+����A���m%6����o�,`5�^E�x�n5��9r����R3�ټ��p(�����UUgrӔ���U�@0M�ze�6���)�0*xI&i�+Yqr����F���T0G��>�v�G�d���ءF����?�J&᫻zz�q9��z�D��锠Z�Dׇ��Kgҕ5�'Teo����_����\>[�����%uuw�61���
P�h4|:�kY$|����i�i�>_:���G����@ߺ��',k�HM�Z��g��pV]?"��xt�ıc���>��E�����,��]p[��e��P*����LȲ��?���94(c2~��ckV�9z��h89~�؜�g%�U�%��m��0 ~��.)�
9��)�C�y�liii���H�5�ط������e�w��:vx�����Z�ǳw�ޡD�¥�������� �0O�|� �d���X,���x���X8���sN&3 P�ȘTj��-p�dz���F�c�jՄ�L��>DzO�iY�\.�Nێ�h BqG#W�!ət�6�A2ơ���P-��l?�q�C��4�:r$X<q� �<84�X���&wu��C֦��4��Z|��Ɉ�<1��j�R�{��xƎ��N��:�+J��5M_US*Ϝ6£��;;*V\rі��BE�,�b�5j���'""��W:��z�Ғ(H9�O% #������*+*.���SǏ�9��p�e䍢P������fl����E5u�WϚ�� �,��"W ��.����m�Ǉ���(�<�.Z��*ߟ�悑PIq4��j�u�fή���%��x߀'��L$R���7��[��CE�J7��=6��f��k����������8���+g̜w�E�|����p�\49��4x�u�ɓǃ������҉�cdB���X�L:WUQ����j���y<���wnۼ~���p�
0=�o�8�0rܡ};;:{�C��c�H��&19"$�8����_����o;}���#F��<m:v>,608���~�V��ɚ�!Hlh�0��%�~���*++[�5����D*KM.	�*�F�Y
�ò��caG�h�ǡ�%�bDZU���H�T�b��W�z��ݻ+��v��
.{����`�'�:�Vת�*������eR�2�T
�v���z=���sA�jk&NnZ��GC�?s��E�T���s��}�=�D����E�@�|�ŎU�)ME���stl&�s���E@>ۆ?v4.��;�l��4q���Pr`�ǧ��&SɊ��T2����O�}<~�D�q(�9�.H
��N'�kEt�9}��g�G_rΜ@0X[۠{�����ʺ��ښ��?_��v����Xi����4B$[�e3��1��yD�����~�f#����>}j\c#�<�5�*�B��fm}Cl���䉻o��ޞ��Hq_o����C��O׵� ��L�:�!,<!�K��н�?�� �w���U��ʪ���%�/Suߎ��x�۫�Fb�������W�cIe
�)oB�E>�`�N!�	���D�����xk+�9��`L��rh�E�9��篭����?n������`0sfL)*
��	ӣ�ŲA�ϘDΤ�j	���[{���=m��^�_�%p�㭧�ΚY3b����T*�����C������U=�Hdsy�� k�5U�?|��sI��(�23Κ�R��u#�	��V__/�Vee���+
)C�����9~�Xey����755�K;q ,#>I��Z,~IqIey�~�]W�~��&�u��������A��m�	����|s��$/a��uK�@��TW[W/�9���Ɂ�>��$�_ӧ�uv��z������A5�>_o?��i[�dz�ƍW_{� T!
�!�	Aj�=�7q}�C��A��eb��P_7z̘����>w��٫�~�jZCp+��姷m�����E�Mjn?���s����xkkkF��Hf��.��k��ᶧM��m��PQ�&�F�ɦg�5��2b�3��M%�GX#-��\U^���#ۜGe�������'�a��M't��J��Ĭ\��v��qM�כH��m�^WW������L�t��_��:}���ӧO�� 
F�3�<s�J��j5���*�$κ�Ryi���DJƎ�Wu�9K_y����G�c���nF4DKJ:N��@�[�m۲宻�ܼqc(ڼi�?*����E��[<{+�}Ee��g��}���Н:u��.$*�#b�RM�\t�,[� �d�� ) ����̸Iö}�6�i>K2��LeS��t�ȏ�0�Ќ�v�C�������ig��A�tQb0^[��ĵө4���2&�F��(	��q�K�Pl�W`af&(�cA(S��|��Ο3:�+����!�Ё�mm���A_���#G����� ����9��{t/�T��@{�{�.:;�����I?�����+�y�Oo�]�l��?�v:1!]r�#\�	�d�M��R-@'KO%M�����І��P����A�'�Pۀ����v����%�����mްa̚#v����8Y>��"'������T�/�=�6�S�G��g͜w���?��Ѳ�R�2��ʤ��?Pв���fc�hĎp?�mBV`_��!)����>�yt0����ۭ-�`a�Gr����ӊ��$��8��o^�`�4��R
�l�H�3�5�A��x8�2��mh����C�����T�d£I�,).�]p�e�x���*Dn�I�e�	�:���f��i�R���xTZ,ʴQ���#���ΊW�F#��c���y.��$hI	P>���ϣy1Z@�ô���"2�Ȉ�Bt���c�P�����[����4�aB�`b(�q�%KU��P��͐�E Zk�W;j�ɖ��@��M+��E��>cΜ��Ύ�ֹ�TU�b]��k4O"�X�K��1kM��a%`�
�"M�f���y� TR���*Od��{v飼���s�t21�J"����Tח�V>z$��@L0�S'���|~�-i�\��(<�"C��"�aU�8eE�m�����_�Ջ!�D&��IT�0����g�u��H"#as�J�[���e�-ڸi[&g��:�8��4�����o����/_~��˯���?&3ɐ�NL��X�`��C@�*�(�E$5���A���������?�x�F�>n	y����n=�{��#G77O۲e��CG�,Z�d�ƍݽ}�����F<��xt���oۮ˂X1a$�+��\6���"j]��d���Z�,�b��ŗeQ�T�^u�T2	3�t�E�=�LEI4�cJ�@ 1���o �]v��/�O*��2eZwWwxl��ڲ]��/v�c1���PW�I��F��:� ��i�a� �����1�y^ܲ�1�ށ����S�-ZZVR
f���s�9�����EL(�ۤ
����0�rd�KIQԉ%�*�$�`�)�-�$��%aTh]�pܜ9�Xqj���Uo�6mzs�8���R��d:�ŋD�a�cƌ����U�\�p��}D�����L[��	�Z`�����Hܕ9'eـL�k䭁����Ͽm�����]��X]H*O�B����x|0��� h�a��Z�R�0ryC���Z�E��S,ZLٕ����ŋ��x�K��i�3J:�p�b}%�5>�|ہ�-����j=1�Q/w&S;zd:�����\
��̤��!	�B�~�@_}��Xo��(~|D��V���d����d5�)D�f��T��S��ʒHw�tX~�(L������?�y��HI鬙�S���v�2y�$r���E#��M&��re��:�;'�(<��\P�ay8�SH���:Ւ�w�ʖ��|��ka�P� ,�	�-�����UJ�LQ�JÒ��n?�;��  �u�3q��Qwޑ���Tb��M��\�'�ԅ�p�q�9g�CQq.?8��z)b����y���r�4:��b��Yn0�W��׮��]��*d��z5��RJI���<�07�-�䬜#��=�B"BM%���Y�ᖱ-DD���X�2m����T1Ee�q̬e�`N�p ��θ"U'��
�B &�qK��̘nC�Y.ɢr�:b�H���p�1��)"�H/[�e9Ć�d��h8���9"gK.��p켑ez������
�U1`��.ޓ��?d�t��/
�mz�h����MJ�+�$�0;c�Q�A1h��� z���6q��@E�- 4YD3Tb^�ͤm.���F�\'���L/����q�p!�`-b�6KN!3/���R�*��cആ���c���v%��"ꩼH�'ℽ@8�$��_a��k�3~4,2�3&G�ß��( L�Sy�ሐx��`@���!N�S��hx���'���ܱB�+b���D������WEj�&#R�.�E��kA4h���{�(�O��D,��I��z:I�j����!N�'���җc�q��7s���p8J�˰%Q�D�Ѣ�
JVc�� �gRb~��R�<Kl_�P���B�H��eK��Ď]�BV�i#�ɂ�`2�NI8G�u�6��AB����������Q!�aQ�c����5����*� ��
�!�W	
�xyە5� ]�*�0>��jr�Rt� �{�"�t&���C�Q���
�!��6�8�ţ0�$�A���(rH�&{m'PT¯�{:�ط�*�_z�b,��L%_|eUY���HX�*�$�ˈ�6�p����ܺ���Ļ��G|l���3$�Op�q�C�{��t*k�&������։�P���X^o@#�'��/��F�J+~��Ŧ����I�j�&�ø> �z����c=*�Gz�j+ G�B�BVDm�����(�&H\�2��?S��g�==W\}��o�2�ʛ]KMo
{ ���1�q��J �i^�-Qv�t ��Hi����h���ƙ��V��R��a2�H�σ�k��}C	�>D+�����PRI����@�u�A�`�.�p
$Cv}�"��$A�
~�	��A�@���T�W�g���o�ؽ#G�v�4I0�L���*@���sSk(������C�4@lDUE�����--���L�����PG��_�%¢&73�z�j�׻d���7�_~�7lܹs�����_��-7�����c6O���{~q��M�4u�˯����p�������<�\��.��X!�<'A��!Dj�P������&O�Y~4�!,`Yp�5qtf@]�����U�M�n�5V(*� ��3C$,�e�y����{��}{{�E�\t�׾v�ͷ~�۷L�0���P<`@w�w�y�>hm==44�޻k���dz��m�T�(T�����/��ŗ^z��^{���{q�y�{<�^x�7��͛o�q�ԩ���a�zF��\�߻���k�byV�������|_|�/>�����v)�H<����;v���#PqK�
��t���f
��r�+S�N�1c(;g� 1�]�}�b���/�����_|��9s�66�v
/�L#ȁ�T:4n��7׭[�L$^x�Ų���ѣ`�G��裏Ə�0�ireU傅!���"�#G�VUV�:ur=p������^?n\ue��~�͛njkkï�>gas�ԩS���?7�[���]oذ���_��W�>v����=�׿<MĂ��!Q?�g��왿`��	����g��@!�=����<Y�\��7�\�p!�Y8u������#�\t�%p�>��7�x��������K���R���(����+** ������-}�ɧ ���>(��{&Nlji99q�$ht*������[���_���?X���-�f�޹s�5�^s����_~��g����w��� Ə?8���>�䓷�v�7���D�Y�p�1c�<��������^���h4:m�TA���4ǎ������O/Z��ЙìL�,1O�!�VZ6éӦ��� �U
򱸫������v�E��b/�����FNa..��4�]��������������NuU��W^����׏�ō9��W����o~Ԙ4y2D��g�WVV@���c5�ճ��ܱ}GSӤ��&�����|}�ܹs~��_ Ȯ��*(�?~3�/ �����2���B�jj0�

BM!OB!x��N���ۗ�X>v���#i�&k�I#BF,�3��߇ 炁 P�P�/+������={6�(�&#e8EL7<8NY�������׿�1VVVO�4eԨQ�&O!
Jc!>?������_�h	�����̙�3i�	�c9o���o�!g��sO8g4������ϿC@P[�B�%���c�0�͛6oܴ�;�v���	E��!�'�����i]�]�U�@�SRd�$k��{3�	�X������M��oQ$cQ����@0�?��C�^{ʹ���1�x�K'���0@�5{����ԕa�g�u�A�k�~��ѣǌ����._�mT����4c�n������Ί���#����w�
��?��{� �o���u�*E �.8�|��x,��PED�3+T���4p���⃒(�G�z�E��� Xb>�k^{���s�6OoV��":F!Y�XR���
��z�9�s�u��QP�q�rY,����%���ŗ��{@���Q�p��T����`�����)|��BLJ�e�/C���� �uȏs��>OWOgiE��N�N1 �ฎ_⨕:�55
qƎ"j�36�T`	���D����2��pﰮ{����:t��{���]?�3g�׿�z|�)�cY,����:���Ob<�y��J���:��-D���Iܠ z� �	��<^"�J@���#��8� ���e��C��t$o�5"�$OĖ"3-�L�64h��A��ӈ��W�aCp]ʔ�7n<v�0Kz��͖i�x���ScqJ.���"M�f��O�v��Vr꫒�d2��Q-ͤ>�t:��yө>7�aæB�������S���H+�� �N�)[�i�I�0
�)�A���:S̓�|6�|���f����>�`��d��(1�<�"x_H�
.�eG�;B�ì5�HN�>MߍD��E�]��\��q��?�ǰ�KS�!FX@�I,4Gp�SD̈I~rߖ���>���y:#�5�F�|�b���&T�V�<ZZ���I-��D��sz2�.. ��x�W]}uoo/TZR�"cQdD�����d2��L􋋋Y�L���t[�)���SS?�H�����J�]v�0d3�.� �GY!�x,��?񳗋�G�Н�W�
pא2G]D}  \_Dy"<r |f�YN��>B��)��[�Ac�b�:n��) Ple�{SqU�P�$������J<>���S�X`��b\6ϡ@N���oٜ���ںe+���9j$����΃~ڌ��EP)0�kc�T
nέ��};�wC8�-��߸��aHU���������������x�h㗥j��{�UPB�AL�d�T���ͥD�7N�*ɹB��9R����zu]^�A%�J�0�i
yAC�u��߸�zꁳ���裏)I$�J�H}�-؜D�F`F1�xy4ů{�9���a��@+�n��ޔE���t$��K�w0p�'J8�{<��/��B_pE�#����s�� %R<���_�i?[�*�-�&M.����իrk�%��-k몿{{�+s?St�S^XpNdF��ߣ'����.u�$�j�O~ʥg8:�Ɠ���]��ݦ�U�=)�$s�Ld��{�x��W�ؼi�u_��ܹ� �"����۳j�ۈ�.�|�%@��|ʹ��*�N9hYy�ْ
����Օ�x����ևӼT��t�٧u#����R�߷���w�Ӧ�OR�)��хg�����o�T���mj�$�m��e��/�}�/��srG�I;vX�D���L���Ǎ
�7Zb����:�v4⺒�z�(�5����d���$��o��m���=Gþ���E�@(���޽������n:���-uۖ$W�,��S����*�UJ&3F�����Bqu�_����ڿd	�F�������ٕC0��PB��h���{��#Ÿ�/���<ඤ���)Y�<vwg���Kο(��y��	(4٣�M�`���%�
�a�>5�%�
�-Dӵ֖�;��a*�������w^�(hb�������~��~��%KCp�#�.��p��a+(����6�kF���P8,���e�pt���z{:V�S9�
�`����& �+Jp.T��X�$�o��7_�����L�0$-w�Xǟ)�d�ZQ�p6CrS4�,KÔZe�/��즃(5Dc�)�nE�P1W��SOuvv>��'.���l:S訡K���--'���_r�%L�,)
�R�{É��Wy�+l��T�M͘�>E����zc�,��7�$�ݨD����I '�h�B���e�+��ز�8�k/�&�?0nb��\�&�ʅ���a�+�B�����eE�٭�b�~�n���K�.J'ӂe�P��?����4O��ҫ#F�M�>C�[!�P"��n��)�PPQ�� I�I��x�v1��Z0.�XM�[�P{�]j�(���a�^���S~L�ۘԊ���Ln�V\�u}���ɓ���:{�'����.S@c+���ao3�v�,����+r� ENPe�Ň�]4�R��E�&D�@2��~uϯ����Y�f�U��f%���R�p��&e�O���160lQ8�!&N�%�U�xQ�t,Ӗt�Vن$9L��,W�x���L_/)'l��3���Ve�3l!�a4L��=��`�r��R钷�i/������Ӓ�����;88x�������U�l���^�#0Er+,nh]�P*�آ�@��6�=9��KR-�s��,2� Py��=�8�_S���F�$�AX3�jX"����C>��\�g6�B#��J�vB/&(lwBL�=�wį�z2�#�̕�DgϚ��;�~����,Ms\�B��>��C�O��}K�H�rV}���kr����\����&�sު��$J� ��n��14�O�<�"O�lHRz�Xiy.��x�@ ��>�͠yU��6(�w>X[���3f�J�VbP��i�"��N���F^�h��KӍ�d���P�sbm��������{�7o^����_����.�u/����^{�|��}�/�_y�UUUB�"���fh3-x=~��ha��3�J%S�lV3�M�4�����w�PL�xep����)S�W
(*V����w���H�����ȍ�.�J�����χT�Ѣ%�����C���e5�Hx�{rΌ��K_�(��l��
.L['N���C������w�9��{�}��&�!-++{�����>��cO=������yc:�v�.T|�$7�(8��$�/å�k�z=�
>�^^�[ArP.�s)0�@CYJ�������ؖĹsJD�Y3Ti�59M#�S�5��t��n�5R
k�FY�Q;��HXgښXgᕸ���?�k¢d!����P�꩙ŋϝ0a��V�޽Kq����pc��|���[�l��� �{�B�"�ʰ�H�Hos���1��~
��)o��L.���k3�6�S����Q�#<+Eƒ��cZk��"uN�x<�'0�,F���sSG0�8e�����)��ah�IҦ7�e|d�pP�ƽ"� �nX|�-P���C�\7����.��LS�ƨ2L)�<�ࢋ.���K�v��R`L��a1��|y�9g�l���q�p�Ħ�<WY�����k����1����ɓ'?t�}���+7�ÿ��o1��H��߿mܸqX �E��_��555�����~��w�}wڴiw�y'�����=��s˧L���_���'���K���OL�<I�BK@ؙ�<�'E����t�#mR=7��6�	� ���$dbۚ!����&%n�}RUB��g��P"�R�\�m�z{�O��v�G}��[oe2i�p���u�]�7o��<}��}���ӟ�t�ʕ?����pU8�?=��+_��O~�gϞg�y����dmhh�R_�[�l֬Y?�яn���t:���oc�3���a*���y�7jaC�D������N���(���,�g���D�`�]�T�0��P Dܿw?���)�a%V��L��rD4����k��J$y�����sKd̤����?�+�����ヹ\��G-�� A'Nl��L A#L����鵩�~ԴiSW�^M���ŀB�"|����ԩS?��]�� �?��믎�����q�<���Yy735찄ʓ45��ÿ��/��ϯ8LS�SLhz�Ǐ��_�����n�������ܳG��u�i̞3�+��B䩇�W��m3���<
e��߀ys~�v= ���&���� �v�ͷ7l�p�����ǎs��QH�[�띵lٲw׬�u�L���s��t�򕯼ھ}��_�u�V�h0�H�C��G�y��k*u][���/����$�|qR�N�xa���q���0�~TQ;زu�=�|��$��>H��yt�P���^�S����z�m��qP���B��xow���
�g��|tm�)����nfS����-6��y��y���{�{��ggϞ�~�������?�J������󫯾����{��ǌ��zb�]}���mm0=D�S�N}�G�̙*�c(��Ə�o��9��駟�bq����>/�Ǹ�A YQ0ݤ����aPM'��k ��f����:u����T0�ѳ�>��K/~o�Z������W\�o����VC����"���8ĳyǆ�%Pu�vOB=Қj:&b�W^y�v�k�׫��{c��.**��m�).3fL[[[eeeMM��� <WKKk}}���e�JJJ m�|��ѣG眆4w����x��{ZZZ��G������ӧO��oi"�Y�)���%J�p�R���۟�2e�1��:|B�g���9rT{{���߀?�,�~�y[{�Yg�7v̱�'��_���]wM������l!�"ʔ2wn�Nz�6LƉ�G���@2�`�D�zU�-�:	����\������M�6���.{ꩿUVV�z�-֯��k��3f��Hu���dX#G6���Ο�p�q���;~�ӟ�?CB0q�%���/ ���ʯ|�]t�?�II4*X�HT�-w����I�&hN?;n�qd`ɒ%��uO,��X�|9.�%B���P�뮻nٲ��o��34�X��g���wr`�&�Cs^TT7�)�5�s|�Ν;����$e�\>P�Nu�˯�����׸ԁ��(@��x�UWqi��[��e-����(��G�s�r�o|����-,Z&k���o��&��1�����7���W.��r�I���yS���h:�!�%26��E�>��Sy�������7�\%r]
��o����/z����娂���x���911���c�ur���x�>�̏?n�ر���J&C�&+�S͙7����ɓ'�&4��>ȑ�.6H'@%��a$���p!;P���1nx��a��,��GS�
�Jgg���m�&M�*M�>��s��X���N`䈑#D� �߄������q/��Md�33v̎�� �n���.ȜUu��C���:eҬ�3?Y��:v�聃g�h6���d9�GO��P�h������S��=qr��Ct��0G{\$��������/X�Ǐ/_~فC�@@�~����R�$��;x�õk���ǁ@:�T6��������ғ'[�}�w��1s�Y�/���{�w�-��w�}/�����^L�2��5����ys�І.EΤ�o����8�i��y��;��%=-������������?���[_���PrϾ�6'�pM�������Իkޝ3{��~��'�\�g��o�1���7������+~��_�}��?�(��(�����H�#���0P����:����J 0g��Y��M�ӟ��0~<���y��g������4b��Y>����'�L���P��Qc��#�<�v������խ[��yz����BW�~gR�d#������AƠ�5����O<�8Ȥ��455q�&�%��|�������>�h��`��s��	�:� x��Ooš�k����W�C��;�)�iںO��t�7��A��}PC����������K|���q9��f�{	l�b�僰�)�CC�_��o���Λ;���C�h:M	 0����Mw�t�7��h�	M�v�#6��������3g�j�����_��CУG����7o^wW�ѣG�Λ���I��d���]�e�S| ���e�6|�7~���Ʃ|��i�-xj&rMM��9���j;����2�>ZGa	�%����-���_�h�mX6�u�5_�?��?��%)WnS@����>Y��"��$�i8T����y@�/Y�����:~�8�o~��G{����+%��ox��M�8��_ �jk� F����e���0�Q�� �W��<��@D#Qn˖ͷ�z3�p����w^Muͺu����e���o�j1nYO��(I/2�:��1W��zRS0�
�^�hoA��P���>{�?����x?m/�TA��O#��t�.]��ss[���z
߽�<��3fL/�(��:ϥaދ��e2C	o0�.·,@�Ӛ��`�w�q��� �"nl�v���W]u�%�\B|_�&L�xf^��`�B�������y�1c�s�몮���l��/�3�&Li<�	�]w��#�Gyt���<��#
���Fp�p8\U]�����/ټqK��CF�#�'@�&��BP��cF�~��y��,�����ߘ2eʈ���q���9�ѡ�Lv�2�1������IQ���sߒ^�\F�~�������r���.���j�������t�W4�D��X\U7�g�hS�̿�ux�9qTA)0���~�a���V��҉8$��o��z����ax�����	�fSߢW{�B[&'�<��y��ýb
S�N�{��O��yD��\A���|������
��Ypގ������!p{������~"Ǐ}����.�5
CG0�1!�A��i�Y����o|,.�"d:ߐ�n�ӧO��r�`���/@��I"���o�1Ͱ��Bͩw�#��5�^C$٦�%��,��Dd��v�����B�+R���ᕇ�C�2�V����E<;n��B���w^H�K�*�� r@���r�z�����1N���=��];�}w�΢����Uo�h9q�7BX�z ���ALq�0�x�/@
�o�>Љ���/E���'B?�X�3+ZbdV������-�@\�>G�{O�7���f
��-_ JF�2��)\����;�Њ'���p��)��I��>䜑����ԭ15����S�Ԅ����"\E ����$�C'N�����0n�9Ĝ�hwE�2qb�ڵ�UT�a��ĉd���^���T&��Z�I�? *%��e��ě+�BZ]��2�R����\ �X��Є���OW�Z�x57� ���h��_6R��=S����wp]��E��.�v��\�8h��r2ٴ�WA�G���	���EpGG�� &�ɕ�aps����� �H��,--q��= 8ܯ��TT�(�gSpw��۱dwQ^yG��"��'I�` �I����U�W�7�c��D����Ïqq>VS�;|�Ț5���'w-��RJ��"j�A�BZU��I�QU�s��O��6�SQzh�fA�YYY	�Q�H��$/Z$�S��3
"@w��	,ǟuu��DQ�[�Ԉ?hc��@d�1��k���.�m>Z�@w<������!�C��J�tM�2u�9�K�e����۲�pDk����?|����:�\��A~�?!,�(
! ��/����p��T��tr�ٌ���2Jgt���Ӽ>�2A��U4ެ�=�T��y�K���M�d��)p�DR,�M��/����i���)���3OϜ9s���tBwg'��:	ӀG׸�V��S��5����Ӄٝ�lY�vvR�hjG������<��&�!�E
j��?����̙3��6N$�:�\�?3[O�f>�&��<�w�äf^�p� "
�rln>)v.��T��(w�)7�S���wK��K �mߢ���^R���p^��;u��SO?��C	� ���3�?�'�q�̳��A,�{�� �W^q�ǅg�CeIN�S�FM��y�ռ��w�V�z�3\/��>�u����.r�#�d[4�$2A�D�ߡF��.�;�m�v�������6	�����Ȕ�>�᧣��Q.�N4���ZD�^U.�#��\�Eg��>
lV8;�.L,d����~��;W������s�UWo߱mٲ�֮���D(�HZy������'0أ��Ν<y*��hW*��tC��u^U�2��p�9�ev��=�C쥔���\�B��(��������Z�9��dE���d~ރ�aA�o�Tr(�I��aYD�"Q?ɉ���^�/�v�y�R�c�<u���na߾�.ذa����=v��?��۶o��[ZN"ꬨ�8�sD�3���ݼi������p$Y��4����P���[�����;wcU&N'R�rF5t�)�m	⺆*zv-��������p{�	V�O�5�.�ִ�X't���W_������!:M��?�SBH!��wu�|� ȇ��;v�x����R5D����y˖MDYE`P����{�dkEEŉ'F�A���6��H�ϛ�e�d*!)N�$���lؠ?�w2�|&K���n��z՛o��C�K����B�Z<�E�����p���aM�$)�IȩC�E����]^��ύ7�˖�ry���4QŉC��D�0	R
�(O��VT�0�9`��Ǝ;�v�I&���=_���.Z�8
���kxaʁ�N?�HMT�*��;o�����M�@�Vǎ}�Ϗc1�I�ʤ���A��+_�ꣵQ��&��D��"�	bE���3O�~�$R���9@��@�}j�v7�P����,>c���l����\��EFE.��#W��N�F�O'a4�t�o���/X��u׏�~��ŋ�\p��&L�P���JJ�PO'�01��L6�U�L�������.G�;4�У�d*�_3�u~���y�%66�z�5�'O�C��_A.��	GDYt��\N5�mhe�U����Jj���,h�7P��J���R�{\(+|�i�=�A��2��pp؄��ܢ
	ʀ��Q��o�/;vlyYY��#���ђɓ�4M�� ill@�ɝ�y���;S�N��Z\���9������@<F��}L6�W����	�}���1LQJpú0���CK�ĺ~��CTHT)1�MZL���`������[o����	&(z�8Ԕ9��z�y�,��x	��ne�<���*�gAG.[�⣏>ڶm�J�}� H:��5�\[�nHT/�|��?��0z�y��q?M�r��J*� �)�#�ܹ�{�O��_����1a������~����y��B)�5�q�	:�!�]�vʔ)+V�`T�F=��#5�z�/b����=�z��'���5��b���ѣn.s����%�i�L��rU��Y���?��8���B�Ʉ>.��kjjn����8�&�^���+b�p �BW��ɒF�S�
EK��9I�ˇ_�d�ӧO������{���d2UUU��<}��FަN�x��K�!<ϡ�(y�yBR7�t�SO=�hCu����2�ncq~^/�6�]��DJKd�J�e�d۔Y(�o� ��i���J;X�:���]�����J�E%G��o����)	��
8�^�dY�PF���B���������e�~�NSQ��y��G������Raݨ L�3�N�#=�_����z�톆�"cAp��	0D�)��SD�D:�H���O~uU��H �#7¬UH���Y�99Bw� 2|z��� ��h;���|���n�'�P\p���DHY�8s����o��ִi��O���K/�hn.���瞻�_��������j����׿vvv^t�E�/�LJE?�H�2���&�wg��a:G��oh�;�B�,�G��ٜ`	|~k������B������:ڻb��e�z����u�� �y�Ĳ��T
�tO~�+�d-��+�RgWǡC�zz�a���A$3�[�֏�ɺummm�O\�λs������ewn�~�Y���B��Ҳ���.�pӦM�-�$�B.�Rn|P��qw��� G�ޚ��u��������{v@�[��n��4}z�m[%�U��91ͥ��ڴ����+���������Nx�
7b�3#�'a�$��Aͯ{u��EiI�/2+~�S���	P�cuM݂����G���0�;wn�Bϔ��U�W|��k�p�}�55��|�k��
���4aժ7�l��=��ӳf6��oݴ	����&V�΂���Y�(Q��yk�y+d@P��۷9t��ʗ_�o�l�2��U�.�ں�g��;��[ovϩ����5
�8�8� ���Ν�q���=yjK�����?���ϝ3��q4��Ľk".[��(��������E�( 2�œ�ĤItB_ ��>��i����/Ovu����wB��gWW������Θ>c��M}��>__\\�d�b ��	6'��$:��92��0Mص�u��3����T*��E�O�>u���T(�~����\ڣ鼅���Ff�BT�es�S�rVN��>�Ŋ{p��}�T8IK�qюC�V�ҩ?b�������s�54�7n�F�)90�Hq�z�L��5�`4�/}g�;E���]���p�_|1�F��'�����x����Q����o���n�#��: Ρ�#wm��-0��S����]tnYY�wlm8]��=��ٶ�3�L�`�a~�gd�/h� �j8OI;�@j���綉ІV�L!+/#�;�����p�n�O�#9P�s�]4e��H�$��|�p�t�(����.))Yz� ��=^���
�K���P�`0�����\~�U`��O��]�#�s�4��'	�Tbz�\�o�..�pk(+�{X�{)4$k��O�P��}�qj��R*� ������g�G��y�?hӯc��c��7э�l��p��v��y���/$(6��b�B�ȑ
�x��V;G��/��ɪ�/��H(���;y��Z���zr�%��(e�ʓ9�q/���cXGx`)9.؈5 ���G�q��Cy��xLD1�A��I�5Q�C�����T��8���E���>����(�
郈?LqQ"X�cK�J�B*T�菟��O������Z���*u�ȹ2ΏH$_	��WYJ鲍����(���>�2]9�6�6�s�"��� S����-�.-q� S'���q4�QdN�X�-:�T>�I/���M�4\fzt"�Aa �a��(�|7g�XA�Vr+�ˋ�E�N�L�=���L��Q����_��H��ؽ-�8�.
K��t$��ג-�Y%Y�؜%��� Ό���k�Qy��]؄/'�ݍ�pJz��,)� ����v��L�'���!R�Q����D�1t�!���+�ٵ��� �n�9� 7&������nd�*�Ie�}� Ms�k�O�G|�ƫ/;p:��qS��(]z���jI�Su�������pQE{�$�=���{�(��9��c2��y�XYo2vwA�_�MW� DE.��D�F�I���Ǌ+�Wy�e
�x�AS%F��2�8���x�E�nMё���}��Z�!��Y���3<�4<��{E���T���'��0P�-���\�ƛ�D֜���:?�A�g4r�ű��1t�.
��̒R��*B70���؎��1Z�l
\N3�v0�J�b�+�˜>}j{{G_o���[8�'�Z�M��V/�p��i�����=��a���-R�/a��y��;^3����D��D;v�ߴ��$
���梑�Hq��(\
�WUU�����vt�!lN%�3f�5�>|���/>�H�3��Q���U�/Y�.�%Цl��&@O��M6���w��i�޾Xi4$Y����<�Q�Dϧ���3foݾ���������՚Ol�5*���!Ϛ�LU?�d0��V��Ϙ�k/d�W�~��+�;�Q��$]�y��p�Ʀ3t�d��S�}�q����1�Ś�($USQB�4�	~����cG!��X�ҫ���ʹ=]�=�=/����=�tڀ�ؕ�%���%�}�th����H=����a�@2J��Z$Z�!W�zͫ{�#���J��zq�C������UZ��2`s��w�|�ʅ�l���,~"���Q��zdg*g�6�I�Q�13���S�$q��Gs���#�Dؠ�^�J,�E�!��Lo�j�H��޽zz�ZN�76�����j?��J8�~�;��h=�}�.x�P�W,b�E��GS�׾����2�&B)�@��򓶨����'���Ç�G�ȏ=<��*����|�a��v"��Sj��m�7L�d�)�R�}��k�C�O��=!
�pE���jjЯ���%QA�(�aQ��UIl�.,1�O�@lP�]q0�����y��]|��Iy�A��C��4B�z`~��E>����j`� � oņ���Q�n�n��%G�Ŋ;e�t���ɺ":9�¸����p8��!��l��k���������j���m����Q�=��p�2�)��`�������7�3�/�<��C����|}��fΝ{��%�����Gq=��Y:���z<�0�Sm�e�v:�9����L��ǎ�=�'N�������4���ď�������L�"���8�BfG�)
�$��Zd>K�7����g��������D�	;:{mJL����Hq����A�y�R}W\z�cO�S6ܳ�ă�����*o%�XV�����_�--����䅋��dr6��O����gŊeL�d�ݶ!��$Ȑ��,A���@"�֨���ӧy�����d*��j��4C>Z��e�_���p_n_���E�� &H�Ňݲ�g,�Y�� ~f�� Qe!�*N��<���h�줧�P�σ����K��8��ު�h.k��s�_�֚���)W��T�I�B��.yH���+���w�b��| ���}�E�[�W0������W�^^�X���3��E�h�������f�"'�:c�Ц����{�BE��$����G����hYI$ݺe���M�y�l�:oq_�ad��(�!o��
�����B�}�D���I��y���=a����,�L�u����Qե�T��i��m��[6_���|�k�ܙ3N�8���,��8�L����v�ܷy�N���w������(c������}�J�ȥ�Yri����Y��ۣ&M� ��_2OA m���2a;'������PUE��G���I��60���FJ��`.���-�6'�L�
�&�D"�$
ͻ�e����kLl�pW���^܄��5�O��ա��_�k��R�dy��iLC���y:���U{��Ү�9��
����3�E�mY��ر��1NBR�k���'��GR�~ /���x��"�"����$vb'Ĳd��6�hVi���8���O���a4�驾}�Y��}�����K��+�e�����'�$���>��8S���`}K�b.����HĄ`e��:����~n8����[?qbFQ�?�F(�|�l�W�U�,�J�S1�&�UsШ��k�WF*�HL�7�{z�ۨb���O%� ��G�*���/q��O�
G\0k!;Vϯ��n�:�X���s����v.����j�i�c�ޣ�Vn����o~�o����tr&�\�A8��}GH\o/���!CLv��F�L
(Ai�00���f�}��l���	�L�Y]ۺ���{���a ���h4�L�sY۴Q 7wlg�@ܑ�Q���{�H$�����)�4)g�#�/�o�;�'�R�w�x�����HX0�k�&U*���.�`]||�˫/��ٿߟ��y�G?��|��O>��U�g�jզ9�z��T��+<���9��)}E�~�+˩d��h����!���
����f��n5�d�0L�Ѱ�8G<���}��g��b�O,�Au��b��l�@���K���/Lؖ[ޫ\y�����N����x��J�biI��f��,���]ȠKѶyM",)q{j���^P�$�i�A�	�)�������]�tgΞ�Vjw�m��I��2!]J�
�б����b���VD�X���;`�����w�����z=`t<>��(  �;]2�K��wa��#�h�a�A��_+�1)�!jw{7>�9Y(���3g��.�z�O�&:�yn �275�v�t �*�D�9���O��'y� ��#�W�9X��.���9,$�h�V���.j�Ga�l|/���M����V ��Q�v,��5w]�M�#V�B�����˧p�����m��cu�1�M�&��5�p�B��`�Q�6��IDd�jj�ݔ}y���d!sge�����7n�y�ŭ+`�DMQzk�ō��bm��PH�rJ1X������+d��%�ѥ��+�@ו���^oa��,��V?91=9s�歛�^��Ͽx�p����[�t���Cr���N�������;�UXe��p�D���1Ǣ(��6�[>���ɨjJ�
��Q�;�n��_QU��n�?�s`\��D%
���?Z։�9^Tr�|�s@��^����4t�/W7�5�3	Yo<R) 6/#��#$&� !�O��A��yx��l.?���z,�Vr��3�ϟZ\z�o�Ĝ��u�7EL�Q�%/A(���,�� ���4�r�3��U�]8~�u\{`2��!��!�L V.��.�t�,D��eż B�B�>�t;�tr��5ƌX"^�܀,�ZkA�Ri�
ق=4yE�-�n~�Y�C�D�ՃP;�gJ-L`	V_
݄%T���=E�D���� 1�Tfo�Px��ٷ��+���z��\�V��{��f����0��(	�u5q��=H#�I�Ӱd.^�BtXD]��9�^�����x�J0�jА!�>��}IQ6U�#�P�H�}Ee^�un�'�W�5f�O����ݵuY��{ݶ�舟�vz��v�'b^Ϥu�3���(GE+Ks!�%c��m����:���[�Dw������F�z��o	U}y�Z���3KI�kԚ1E��j2v&F9�a�&��x�q�|n2�H!ZI�����H����j��'(���������U�+�]��L/�-&����F� �5�O.����܀�!�4ڦ�s�u���4Y��T]�AP�ː��8,0�:�=dM9,��h�s�u=�m�!��PyF�{��.��x���mG����M�Q���<А�nB��rs�CJÇ�?��䢱��_����V�ѐd��$Exd�m��;G �#�vL2`���U|�0�%>���h�S���xc��}d�&������_\����W�FM!��t<>��j�^���v�"����:Ls�ma�L�'Z-�@��R$�͑��$����-j�1���퀫Z<w�U��ZHd��݊Y����D�d�8$�(֕���#H�!����d2u��7���k���y-az��;^x���~�j�X,o�/>���`�Q����֖W�|"��kR�"\Nv�X1{�������D�ȪDC��(Hc��
�(�(r�	�L{������H�#�XCȂ���@��F��$TE�l��mC��"�Fxԉ��K�o�$�B��p^�$��:;;��@��6����>5��/��;�������ֽ/n�?Xk6�v��(<�W
��'
�����?���ֽ�DD��p�7C�a���RU"�����A�Cl����Q��k!̡�x&*�a���e-��x,�����A�X��5M�?�H�+��\X��X�ϳ���z46}b^�<�2��o�����6�m�_��v����ʿ�㟝��ܻ���׿�%��)2I�	����f�c�܂0;&�O��F�}湫/�1jF��'jI
#�K���wCQfM�YG� %-�����vg�d@.��y�d$ �!�9��t�������:v^���ġ$�mY&ܩ$#���/���U+;	����!c>�B%!l��{�&� <�����v�[*�J��ͮ:���Y�����#�bT<�b�^��Q/�k]f���k~�?}���G4����J�3`�J$C9;;���1�pQ���0��&��)��r,��c�}�$�sG:����5�e*�s�u��MxL`�����|2��r��(a��H�Q�ɽ�u�T5��x��"��f����tx��/>}��w�@̗�=���{�ffO�w�݃ڷ�?������J&�nJءG�U:��`�}�0�c�`��0��ĽV	�V=H�C�����~̞<55s̱z�I�0h�dU�/����;�    IEND�B`�PK
     uK\zn���1  �1  /   images/245bc533-66be-4bb3-b22a-43c007a581bd.png�PNG

   IHDR   �   �   ��q   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  1gIDATx���\e��w��I�ѝ����$� ��R|��3H��E���.׺�ug�q-�k��轎p]dFQA����{I��W#D:	4��鼺���{����_�>��9Uu�*I��N��Ω:����������J	�O��B���(S�B���������rȴ�y���x�#S�����8ۯ���Z���_X��)	BMa
Aht�[�����vݑF�$���i��jgN�eM��X[�;x\��3ns��1�u�C��)by����?B.x�j�~��o��y�i�N�(����{ �Y���_�_�p�,mZ(ӝ߽�s�x�����.�#O���7��:�dC��}��R[7͹�Z��M�+?�C;�&[cm���곗R=��'��g@���J�M��i�[~p�l��=���[�gr7<ߥA������c�çR�!��ލ�>|a�� @���K�\S��6:J�vC,�$��4�����vC������_�¼B.�dS��z׍f�}w<$�����ű���~h���eޣ���O=%���^�:��oA �N��F��e��ӻ岿�؜�s>p��A�s�=��Z���������B^q�j����B�&��!�����_1�@��=�h;�n�,4�Jq�U��o@ȥ+�5_��|f�i�Y�߇ �r߿<d�_��u�����nrHzw���WK����)��;[M7���S��Q���{����ǿmt���4��o-�K6��s�12���u������rl�) %����!�j*݇�7wQ}����t��S�����¯_�)�4V��Nb��)x�!�����/�5$�f����-|�P�:���`�������f�w��x�|���R����Ȳ�9�瘼�uG��7Δ�W�/+gIu]��z�O2�3d����B~���'�@�ذt����oX\%g�[#�WK]}��@Gۈ�t�ʡ}C����w!���<w�����L�]m>��lȥ2���;�mE�B�z���}�|��c�0I�������!��X����8㞲8��"Gc�q��>�z��?��Yu�P1]���d݆wI�+m���5���-u�N�V̒��gʚ��Ȏ{v��k˫��y�ÓWL�xņZ��u)"�Ѱ��l����)�oɫ��v�Q��B�HȣDrCI��s.�nH�<{w�?4A$���hu���\ ߈�!�7�����M���c0���y���>��� �j��#M�	��c�1���^�<!�U6ܸ��f���ߐ� ٮ_��;_�ͱ�¨���GC��ن4Q@�.��A^��4�P���յ�P�%
 ױ����/�M6���^}�L�{�/����2{mo�7O��lw4��ر���_��Ɠo���C.��'�R��J����101�@���ݑ3� ��Y�����7^|�D$��s�Q���'ܘ�EU�2�?�h�ac�!�Co������tH�X�!&�82�#���oH��3����̅\� ��o���6�{�X�8.w�������#�mPZ���t�#2��N8N{��K\w��o5����������w�A*\cǖ�P�����ǡ�'p|���<I���5�	C�t�8���شס�)��=�e�v:�#�WT���q	�'��u�F����9�Z$���j����>	H>0�˹�0d��Xq�.���hNlD�1ᆼ� �@[�&0C#B�����vz��7�Id�x�Q�k�K��M�:��a�Ց�^����ϑ��&�{��M�����o�F,�.0G6*�`�Zz2t��s��l���7�xt�;�������ups�4�Ә��3��kB+�u�96��C�M>$WyطΑ	r��u��b�'�B�4��ɮ���&��o�,���raf�<�I���hL�!��@�%��� R���k�Csq�\{���WbáA#j�I�al��h��y�Z�	��(	���P�/����?,�C���-��l��
찈07�S&��W<�N8ls�߫�5�<�y �6��\{��F��1n�����j��'��+���%��L'JﺏH��1i�>#k��?>'T⃖(�h��sM\G��|�7�0\�s�[ģ�������3����8F��}z3�J>Q�ƒ���h���2W�r,���`�'"��a�d��֒8���]|�hr&���	���ٶD1����ۓ&������U�K�"�ky�|�	o��]�i�CB 9�q���Zr"�6V��"ќ��p~ۜ#S��:�з��ŕ����-��P���Zr"֦��g"dڔO-�L]w�3��u��w=&�:��6� *CK>����#{�߾��������>��&z�Ģq2��{%b�(����"��X#��u�3�3?�l����7wm�y��H�	��o�"L�螁���dE,��`g��`�C.:���:8�h���y��3 7IH$�3E3&��1��灿_4"���ۑ�ڳ#�Eh�74.d
:�p�8����i���lp䂐�(��>�|����ȱ%�o&�uL��|�EHWaP�a��Co��=	cE�]|:C�L������"V�!�~u�͟��"$�����p*3hd��'3H��������;��IRSA*O���Aql�51sG�s��]*�o�D�\s&D&VxG���l��pn�ԍ�}t<V��5Z�Ae�a��vk���!�R�%�@wd���=tl�D#g�҈Qz��'j�}[�,��k:9�+��ɶ�<:�7&�a����,a��X�ƈ6�.�	�=�Ƀ"kZ�&
f�k����p`���K %�n� ��:˪�e���=���w�K��ܐ�$�L\kD"���p�!%��y�xhM>$3�c�/���r�t����,z�/>�m&E�������PN;c��U�Rږ���\V�8*�$o��i#����:LS @��v,s�b�����VA��f4TD�������
�v�9�]%[�+���L��?�r�g��%u	�%�04��	�#"pI��]<|-4�s�P�y����аZ):�No�!�lB�mx��T�k�6}n���2|T�K��Y�J�V�x� ��2�%'p�7�?�<8&|06���2�j| s5s�|�Y����:�4����?6d4��m�l0y�u�3�6�5=��	h����\K�΃"4���d��r����굃'�F�0,h|YC4N.�4y2h�'��.69c6 /i�
&�x���O՞n0��9ÝY�L��"�΀��LoN�La~SD��d��I1#;��u������40ѫ�M�&f�q��{/���ip�=��2}
·R�F�+c��M� ��i9��I,�����d����Z!�jM�Tf�i!Z\�8��հ8��TQ���/��6��%�h\��V�_Y�6h�|��Ѿ��"Qef֫s�+B+���2����ur'�"3�@*2T���ӳk:����B��n��	���X?m�}�Q�F5���J1��V�G�C��`��\�#�2B��0��J�&��<6��&dZV�0�TC�w�#��1�W�.�:�h�ת��+u�9�4�RI�	��LP�-� �׬�xn̻h��_21p���c�O��*�TI�''���:���'�X3?1K�,�����s�[��9��Ҿ����|w��8�^�r�"veiq�l�X��o���^fʈ�We� R�
�Aet�+�T�+8��('.�t@y���~�ZԴ@�.l4�t�.�'(�IE��T֦�y=WhS�KM�{��g��!+P���&���h���Z2]����i�t�VJ��1�}��W&La��;<x�`j_OGj8�q�y?1�=�w�3~����T�6͕����r�W~�:&_a�5�G��r� ����Ϟ�bO��Z�}�UZ��N��Jڡ;�P}yǥ���������O���߽��������%n�����g����J����ߙ�:9 R�IO�B0B+Ø�g�'�]b�^�5�A!bPǏ�cǎ���̜9S�8c�TT�ZdM,-.�cop���vHNh��g�g��[}�رc��2a�����Դ*��>��:.��5�|����c����-^`mm�9��vz�j�>}��k�ɢE����L0���;��f��.����v���f�3I�mmm�>�,	2(h5��} "A���nC&4\__�̞=G>,s��u�"˗/�}��ɜ9s���xZ0���0a���[JQk%��F�}h+�����2PM�f�$B����4$:z��!����466:GT��@F�77'j��~޼���5k�H��X�(��ģ��Z���^HN�����Vq�A��̍����$dZ�������Y0k�͍ÇS�{��F��á�8�+�E�g�tWb3�tۀ\n|�G���J��F���Kz���[�t��.��Z�x��l���ym���j�o�X>���7&BavK�XJ{H��p�����Jy�R?$�e�Ng���P�5k�O�
�l�J�v�r����
:6a2�_bU���$���䋏u�I>	���->�z�����;�V�*K�h�ʩ��9��5fc���P֎��E!W�T���3;湟OL'�2n�=[$z���č�%��/���̅A$�'w%ơx�3�D->qu!�b�r��	��a)�����ioo��EB2���.G��O�Z��H�b��D}�?�IlH���FIh�[1�9��%�{���M\X̣(@3�R�H��N�����r6#K��H���0��~�)�e^Є�������d�
R�:�I�v�����C�H�a�
i<s���?";^ٛ���9\����93uY�A{���Q=y������rG>�$�m"Â�(�T�斢	Da���͒�����Μ(~��	���~D�ޟ�Lq��@�L�.,�"&ri�$���7H"�E���_����'S_�R@���h�¯rW�v�ju}"�r��L��ԟ��M�����P� d�����v��Y��=��4��&�/��(�z~<�mMN{��l]����(��hP�lM�(���A����Iú�Iu����I�+er��rSV�P�����k�UK=��ll���.%���ɅF��ɻ?:+j�(�0�I�U~Ǟ�аn\�\�_��zθ,�4.�/��UH���,�g�Vh� ̘�y.ȹ+��E���G�(*�P�)��Cl����s����A�3?nR*�;�ӣ�\h�����Xh���A�������Қz��
� �(������,���Z�)[@$�2�E��Z�W�'��3t�Bzފ�:�1������Y�O:��G^H{_J����,�����ƹ0�Z�)N�������K��~:�����&��8��ħ�{Mz�t�/4�ZR�!���r�1#�>l��w��f ��l�^J���Bd��"��r"d".EڋW1{���1��N٢�D%b�8Ɖ���0�,$����ܹ��J	�f�w9�+QD�+��~S�n���d1�K�wz�$�o/�i])bQ����oe|)�z�#W`J�&�r��(���%9f��GF���ZC0�n��=�b�y*�D(E.�JQט�o�d���4��^�8�h�R3���t%����@������$�obv�S/��\�C�t�RC,R������N+Ɂg�M�}؈{��(7����X �p�!;(���' Q�ɍ�? ��dR똰3���x�+���� Y���" ��:@�N�u�,T^�O!&���K+�3�v;d^�[e��X�%Xb��!�!�i]��$�&�3݋�J&�-._�B��ӌXeFke;u���8�v �h߾��Ds�7Z�1c�ٓ\!�w�<��I�qZ�,^�P���������-4
�Y�3̞N۵k�C����.��+8vd�h��pZ�q:^)7Q��q�m�:CM"P��[[[��B���v�����f>!���s�� ��|���"����r�x�ղe��ޫbҪ���絿�8-�ڟJh �b��{��qCE����������6g{*��-� ��y��8���H��b8�qZK�S'��^p��;zN*�P��
Ǌ�=ΖXzd��*Yx��졁C���������˴YS��_됁��߽���LҦ��d����W^x�y=���J�x�0ұ��SĊ��%sW̕ާ{䜑�2l�[ot������[I��C��95u�v�٩}n��}���X�V�{��7��`O���\"��N^ݾ[����i��i|�=/m��yֆ��)bň�������+f+r"��us�P���R�̅3e梉T��)��U]W-n� k��\ԫ��[�c{ZC���M����c����߼���1V�g���sWΕK�xI��Pϐ1K;��a޳�#��Hj��7>8�෮����r�O�k���Zgʧ�B�ѣ#���D%�����ؽ�ڤ�fb,��p��
�����}��t/�)h��~���L��� �|Qy�<AF��dt���۾�-��]Cf���ฌ�3��1:�I�����B$b��bU�T<�;��0�QW]�*�e.��%9�'�H�z8��������dsj&��q}�T/m}I��?2��.���fDR�����F#;�pm�6�8�z\G��S��e�-J*�	���]d�����z�{<}&=�!|����0����� f[M"�}�D�8mu*��^���&s���4�}Nx����$,�v޽���CA�e�Ii�D4�jE�|�6�Aɉ�c�Y/��-��S���y�����Bs{��?����}pB��0�ut�ь=��IN��na~��a�9�	��L��I�oj&�	&~�TL<��>3�	�]��RhD"&eѺE��A�� ��2U4���^=C|+ds�m��B�@2jY��=�$����f���c��G��s�Wx�-��;�p��|�{�J44���� �:�A�A�ar��6�h�j�A��5:`&3��k���O�T=�u��&}�A�ygh����Rta���E���[9�hL��2����8���/�]?۞l��`<����dkT���mp��s|"&��I�t33�b,L@����ꅡ�1}�4��?!�ouj�2��k��p�/�ۋMvCA�w�����Pt��4Ґ��h����ٶ&d�ؖ���r�{�J�&x_���I�*������v��:F�B��ڮ�zͤ��F;<��A�VW]� �/*"k󓛍`���t��c{�����s!`G��ܚ����r�=CpM|"i�p��d��@}7bo�̰)��$l�J�^,��9��X�_w~�#,]����51��Փ�kvO���04�6l��y�)
�9�1�TԺj%F��趶�8
���O/�C���/�6>��d�;U�F��!c�(�k�	�G<f�����F󊿴�s?2��ꋷ�'s�n��Ak���W �0)��h@6mP4l�&��d���H拢��4Ȃ�0Aփ�if�v�!��Dwh�
�B���s��{��y�j&?�5o����u��R�M��w��͙/D"7�m���M*{�7x9�!��k(� ��ppF�<@.n�?y� %�����$F����Q���S�������G�LX���?�1�ߏ��@�Wh[������_�z�=�{y揯���G���XL���{B�|��~�}@(N�ȀFB.z���N�ag[���JɅ�^�uw�1�(<����0*��C�8�;�y;�'�r�KH�Zr���|�e�+��`���:�!=m������W�u�@�t��e��g���7(S�<h,2��Q�֠�ptg�F���h"Й/M�/5���3�t.�j��Wˈ�?�l���R1 a�B�J�
g�$�-?��w����8�f�P��#L��^�Z}�6e4�u�35f���' �\����a�b"�Қ����K�͸A��������x�"��2��Z!e���V��N�CSq�� ̻��)(e㔜��O��f;=�ө�?���$�l��C�G-8��dh�=V�c��Sr�7R�U^��?��4� ��T�� :@|�@s�4���y��%�(��N�
�v>1��'H��>�t2�Xh�9���|k�M���$Vr2B@L��k=���6�J���q��C�s�2�C��Wsr�
	��GӄHw\�� ~7o�2}�,C,Rbvl�r�y�hD�[-�gaPTb����v'S?��ֹ������p�����[1/5�A��F%��PM�g����������!�Gp9p�ǂXl�9�Rs�!�Z�&�WE���a��c�Ҽ"�@$�R�� '�hRS��L=C�䛾�)m�K��J��o_o��ũ=t�$3� �$u�^@r̐�#��' 
[��GS�9�Ϫq^�IӅ��x
S�a}�ɁBщe� F�$��E�PIŅ������������\�
H�CNh^u�U���9ZL��
�ž׏�eL4�?K��\hH�ד��X r��Yh&xB�BK��.�(J*M��9�
�o؜�nд�B�0�rҹ��\:��&���P�S���(	b������>GKEI��s�0s^�}�����u.d!|/p^3����gF��	���&|��h��%C�|�α
D���e&��X6�S�YEq '����%\y�o���ӽ>VjF���>�m�07�P�&J�i��ĩ��«O�Nma��S�X٢f��1lq�h���;��hmN�Vw���-��u��k�0�г��;϶��aKH�%]y-�1o����!�"C5��F9+�����-��)Lm���Ẁ��'�J۳��/�L�\�f)8�q�Դ&�V\�R�;��ꀴ�,ym�r�0�@g��~ȇ��O��?��޻5db��=�^G�f_���j��`��+�B��45K7oH�I7�hx8�`��	��_2��-��feZ�w͗ٮ���<��B�v��
jH-6��B�2���K�(5���4����M�3�}�_���%�h�ڙ���B�2�јawt��|��M��l�'}VjԦ��Q�wb\c��6}�X/��������޻����7�0�{�<Nh�U��O-Yr�������{�e���~c���@E^�ō�)��m��V�l�L��k�E���oq���mK��x�&N;�����&W͑�8�]_�i���by%�y�*�L�٤�,ǝ臦�I��
����{�\qჷl�\ �z����F����~����F�5 ��f*����h��5�����Aŧ!��#K�	�Ax�& �@HaƑ2>4��Ш���^{땩�cX�L,M;���P(��^@ hu�B-
��	J�Q�A��3��X6����h���>��|��lL%��w>Ik�rR�ך?�)��K�`k�0D�H�]���
&� bXAN9Q�t�?¼_�h��� ^��� �n��S�f"~�	a�L�%Y_�M�'�>����b&�4�0șX;J���3͋Ѡ�iR��~S��7��V���UTئo�z�����mA\λ�o��w��r��"�yu���6]*�oҢ��&�Ɉ����j�R��=y�il
�����7p�횦|��n/ȠS��sE&lb����٣��$�r�{��͙�z.mLM5�c�3�� F��ǁS�y/ű9"阹L&��B!gb�T���;N;=BʹPЈ��BQ����D]P����
�kE�J6ܦ��e
މ���E@bqS�Jan$�e|�8^�کCM�f=�=�]���H�;��QW"���h���u_l����=�E���<��$k;��P�kI��	)Z����� *C>Q�3��;��I�5

Y.�^گ���+�NZ+z�/v�� hoP{|���{�v]��W�yn��5+TX�w�<�y'��nșX$�#O��P�����"�:Ș��ޕ��p	r�1��yz��iTN�s����Z�����s(U���~�����W��;hQ	��6�t@6�N�}>{�{?h�3S3kQ���Q`�.f��H�S��
��y[q]�$�tV3���ty���_�+�I�b6��Cæ�y�K�rY�>�Ĳ���O;�l��J�j�_�祴�Վ�������1�ߖ�f/��1-[|+��&V29�@����Z:�\E��z=��Et�N7t͝8�p�Z�&z�	t�	*�3����<�Y�+����8�����؈�ZJW,u�œ�{�B]!5��∼�D�����MvպqB����M�$S�O=��9}��L��t��m�ld
EP��R��ų)j[UVj�:���{�BV��d�{��m�t�NC��C��f��2�)�e��ؤŐȷ�Sރߦ<dR�<5Yg��e9�j��<�۵�h}�t���}�,O;�k��-�/�Z�>���S	t<��������ʃ�1,dA#��=/���qݖG�6Lw4����C�늛ߟ����9˾
%S�ź�H��*���nC�t������s36gIS��=���`�������^�M����ly��ny.�j]�p�*�J�y3�jN��X�BI�U��i(|�1��N�p�4U�����?��'���`^�-���X��2v��oZ��O�)σ_|Xν��T%?H��o�^��N�SA��)@��R�)��!*%S��gQ0?� �a������	t4Ogj�U�zМ�eJ�1�
wd�`�!y�U��=V���Oʑ��Y/{�3��\]{x|$�86d Ò�r�˚p�&ű�j&@$�;�;�e��5>����Y���{�Y�	RV��9d�.�z<A�����Ƀ���X,��^�ֽ@�xw���
l/��f�W1��@]��7Tpr/��U�;%sr)[��~k��U�f%x�i*��i��h��a��l�O� �^�NR��%V���P�����Qj'�u=���9��]]�Y�v�k�K�'�L
d92���x��ƥn����#e�sl�\��6Rn���n�<���?��'S{ͮs4xy�u:���h
��>WGTזˊ����Yx�w��P���m@���/�������Za�<`b�#�A�g"im�̙$��8�6��@�l�O>�	�^�=����H,����]{{�b<�����iO�ؿbC��:�F���N�v'�c�p&!�;(ʱ�d4�}�r��{�=0�� O���ҕ�Yƍ5�;��RB�>�s�l�5���w.��A^�O^|�!
7��Ee�@,��6�&~3��u/��O�<da5G�D%�M�|���E���=��D�X�	<=����_t��^!�G�#U�����S�-Y�<M�g�"��O�!O&D�o��T�j�&���!n*=�J�l@G������C�:ܙqi=��*�bݟH��F�N�%�a;;�����<th�f�I���B�(��&r��c��Ch��^��L (���D,Ta&�k�Agk��7��RV�=_֜�H�\�_X�ԙ^�v�OFy�_2f4V��0Z1�ڛX� �](��	M,�Oo"��]'�@n�|Zu��1�;���
aÚ�R�m5���r��8~Z�*q|q�Ohb��S�CC#�y�[�]�P����n_ߠ4�}G�V,�������n�ɈB�3ԟy�aݘ!W���t4��X�Y��OhbL�������J�,[<S�g4x
����e����ɟw��y�'�oq#L�.�<��ʃ�τ٫�M`\�x���VT���'4��"ƪN�'��P�TVM����!�����?Cjj&�`y�t� V!�	C������<���Pv�}(��	E,��~h~�̮����7 �Óm�
	��f�;��I�|�J�p}Ƙ�=(� �[�%Kj��*����`C��s�U1�۪�
�^^E���*Nޚw�!Qq�H���^0O�%Bb@ٻ7�oyF֕G��|�8�1�����)W��bt:!gb͞5M����S3&��j�q���L��$�w\�P�E��	u4��~8sI�H%��<@�c\�cC���I}��~�������3�Ҭ���r���?
4�W����P�"N�x�n"��^;�z���C��99o���J'��g.��x;�L�0=?��O
&O۾��)�Ÿ?��S���b�c#�~�K��6�ؖ9O����y렧�`hhX�wa/��}���f���)yJ[���"��KP�lI��~�U�@�ŋd�O�	TxG[pJ��<'�<��E� ����^�Lz�G�ŝ�&��O��޳R���O��!�`J�Җ'�����zd�M��7�m�5���`qE���}m����wG�D��<�+O$b���J:�j�iQ�i8�/>}��<�+O�`	9Ϥ����l@�EX�aJ��C�y����*,����N�sr�Sy�������/�87F9	' =�d�lR_�Q��$N�S��)�����d�<�^�%�+�����TFuD��9��Qbmq���-�j���d2	�ڒ��N�@�v:L���`ޞ�)yJZ�-�sx�1���?�V`�xr��)y��<;��Ur�*I��2�)d:��QTi:���^�\�\���Nklw��!o���a/�^?    IEND�B`�PK
     uK\qyဲ=  �=  /   images/51c64262-e188-46ba-9658-f0d60e053320.png�PNG

   IHDR   d   z   I>��   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  =?IDATx��}	�\Wu�_��]]����־�ZmI�lc�8H!�5!�0�L��0L��̄a�� I�2,� 66`/K�l���Z[j��������ի��nu�$�/W��W��{�9����kǲ�`J���E�J�~�Y�����b���b�:.���ץ^6����~���N�7�S�؝6��24Rɴ�A�fw�'�&mM��f���}@g�!�V���J����9�iz��?�~4�ɠaq-�׶ 0��#��:#@��	��aɆV��p�q��eA��f��mM���L�0�;�M$�:�����8ѾE�e�Y��k��u�8���/�3��
9a����!��(�[�\�w���b��*��8�z
�M8��	tu�(��6����XJ�]x��wa�{c�\<vU>���HB�يs�:Q�^��:� ��"�"��*Ϸ�mƩ�.��u)J��W��X��]�;�~��O��-o�z�Y*�����L�ہ��2t���>#@��M���p�����=�u�V�����(�-C���H�V7aǛ7a��aw9��1pe�t�'��4W`�%�y��h���*qH�A'����1ER$��S=x�GGp����h�)�h�4�����T>B��)u	���6�w��~��X��{'N	��|���:��}��V�"R���x�<
� �WQ���?���*�=��_;�ӡ3��B?�޾�}��R�a�d�#r-#HZ�m1^��^e�D^$U����!a�����(��E&:,*�X2�9�ɬ�k�Y�"A�
�9Ȇ'�M��Z����CW	�f~K��hl���G6��Ǆe�+e��הi���[�֕����py�X�*�������֥:�I5C��N�=+r%��%u�
"�����p��h���mXdԹ����ZK���8,��֠�݅�p/��5߈0Mf��M��	w����hX�Dm�%�VV`8��K	t�M��B�DF3�B�؝V4�p�i�խN��l���X��)\=�C,��I?{�DH��(,	��/b���E��o���[�1?�Ϋ�t�Z�p>#�p�.�ԎǺ�{�_Y�_���O~�8�R�p��#��Җ�BCgE���H`ɲfEH�;W�
<�[['��E�ç2k.I!�I��W����2�l:�g+�2+�8�jW���p�ِ 0yM���Ȯhp`���X��-����Fd���vT7;�d�}�=x��0�;�J)3Q�$�B�3����^aQ�nJ���
�m��L^��o�9�3Y���#����c��6x��J+�]�G*�Ex<�Dt}�Gd�dD����{~��^�ٝ�#CM ϶�cQ���kDFv�w�	222�U�K��Q\�"��iҽi�����AM�/}}��kR
��[��]��FƝ�&:�}~�du�4.w��Ł�?
��+��}��UW-����U>k5����$��JE��k�@���ۄ�Y��|��ãi�]I��CW����Y�ZGl�QM'r�un3���D��u��~�'r�㔒��f��*��c�;�x�+�J)3!�� e�^>3�R8p҉� �AM�[�!$���.F�����4e1��,�s�2V��A�z�hVc&��6�(2��_�MgU�RV�^����0z�����,��*��e~:�XJ�O��[��a"ê�+(���/u�T��ۥ���E�<YP�����O�6��I%$��S�A���RwKHݑk��H%�c����W���d���2�� (�ֽ�K�xDm�*ɲC��ĬA����r@�j���+�b8�tz��.G��d�j.�#(�JƱn����)�����,u���SR�/K����G�J��/'�.&��YD̡^ޓ�Ly�ax:N\{Y�?J������eL�u,�����C*����5��l�_gH&�-F�,W����ٌI��j��#���YDo��v�,H�?��3�:�o��OGa�@+��@ȋR���h���w���z���y����q�1����M� /`��R��75���^&��@��,0<�'�mR���5��l���\��Z�7�J}B�a�h�`�n*�;��C�~H�[�6k�9>^�bׯ�U��٘
��V�njV�t
��6�T����y���[>���������)�K0(H�Ku��� �1:����VF
�#�H��!�X*�{�/���,sF)a�h-;�V�Z�dp|E���A3�`n��J�3���)h7��wj�&ڑMD���2I����fA���l
)�>a��Rk^��A���=E� �`���B8�N ���$cA���6g(�rci��8F�W�B8s�Amyȧ��d&�L�G0x�Rlp `!+#IQ)����sVn�߇X(�s�����Qf�̈�Yd�3�y�E��;�Ә�3zS�������)F%?������Zf�!�~/@�9���@�i�:�-�͌�p�sK��tY�E�"����U��d��屩�C^�����)�c����!�v��ɐ�XJ�&�d�.+ls,΍%�>����\P�7�*R��oI}�Ԥy�ZȘZ��Ξ�(�)���@����V�̧�0��t���bÄ]��CT��XQQ')rt�W����LA�Yj����m�^����Ѵ|��|�,{`�>~�9f��aL[l��5+Bh�.V�DT�)*�ԇpȘ�\�%8��@*��n��[�؉ۼ���Pa���F%4&KlN����9+�Y��H�S����+�R�A�b����p+Ʋx��T˷{̐r�R��m�S�49�~ݼ@��Ɏ�����;��OV�`�eSE�,�}\�m�������ף����tyH�{Aր=�3�F��V�z2���MM�+Rˤ����u-6�x����HM�B�,Z�����@/��&��`���f���h�qQX�t��yfD�ƚĚ�b`�=���-S(� ��/���V�zT��s$�8'Q	?y,T�K00đg���6� �qq�0�H�徻Ǡ�
�qX�M�&{fM�O�������[���,k�*Z�_ʵ�^]ȹgX,��B�I��u���R��hW|a*oRy������lj[�F��(<��TBk�N��=��"��۱�}�`Rީ�R�MG,�|\��KC�͕��)�D��LXf���N?�Ċ����N����ڷ���/�q�@tF?YQ���yD���y�c߄1{o2
}�߉� h��:,ǢT*`��[���J�帔��g"�SX{W)*WJv��n�%Kc�Y�`C��]��J�("X|�^�*U>��L����	;��R�Y���T�7�/�p��h�z�R!2p_�C�U�Ë��Z�Ď���J��w`�|R�o)���:�E�
\M��c_��J]��*1�hH&D v�EH�0p"��H��h^�1��B�[p�_�!�M�'5��LD-�1�3B�T��R=L��DGJ�}3[H�(B�o]��B#����9�*Ơ.��ۂ��޳	�2I�X](f(����鐙>*@���!��RokI�U�~H�k:A_��e�cb�T+��9{��4+{	ey�aAJJ����2�E�x-�
Pi�M���hF���y��s�FEɉ�
�:h&�~N�:�Y!0�_��	a%�x��e��n�
���)@�{�I��%-i�٣�QZt�t��S|�?��"&ȠZk+�	a�l���bJ��F[��xn1�b�8��1!!�|Gp���3BA���!���RrD (��Q�r�w�{�Pԓ/�'�k1� B��~^q�J��Oځ����Tf+3jY�b���O��2'�r3�a�.+�]jBfq1dds�r_Իd�ZD7��BɅ�s2ؖ�2B������V�6�x�qV�����撜�/�D�_�����M� l@�Cu)9�,��Q�����J ��Q�/����r;`�~Ex��
g�61�mv����h����>�&|����X�(���7�~4z�zl�ֈ ����\ 8�ڛU�h
R*`����������#�5�E��83��	�ь���
�K�!��	�V͑q�{K�� xX��%H���{�6���#rM�O�����,���\X��r�����A�/}Uf�*e�BH�@�?Y)%��Z(�ɮB���:{C�^�ţy��@k�/��D�ӆ�,¿M����̽)�jfw��{F��٣B`�n�����a�hBIdD3����aKZ�J�eR�˵�|�kVޗ���I�٬5��o٬�9{��"�����+t���ϨeE��#�ta��ٍt!_�ϯT�t�[��HwJ|t��$�
�R=N9�x�w߈}����|G��R�\�l�x(�H� "nE߳���c���	Gl��\���qA�/������˒x�jo٨��h\Yg��\�E;gV_P���&�D�$��K�Oq�K���~'�Qљ6:җ��&�#g\��L��{�xa�8`�jjk��8\.� ѩ��f3�����M��k�d�]#�1X�Ոp=6�ʊ*��6'�4S)N!�I4��HO
u�|FL����Ŷ
����=?&1�����Q)�a!/m��P(�˗/!���񠭭M�zUv��aM�%������y�өY�dM�-),��3��aw誀�-�jY�G�X��c0Ac�02����_n�,�EE�u�X���U{�,@�P�bh��pcc��aei+�#��r
"�)�&d�!��KJJ������F��,+G�������o��J}�[㆖��[�	r�t9���Ÿ����}a�T`�O��D��#�����H"RJ��t�乌R��a���ӌv�t��z�$��> S�� zbc8�;��E����,c�4�x��2%�� �N��u�PT�����-?�@�x��u
�X,*3�z]Wt	r�0��D��DNU����R��nGcc��,����n�x�e�TB��c�.����#��5��d�w�H���1�)���B�7�conD�f3.|F��K�,Q`s֛ g���ѿ��x��vO��W6�"n$u�LgYK.�`׬�K��a �M��W`�0=�#e���"� �;���d<���1��p�_Lj ��H����U�*#HD)����X��� �1��ftlT�d�jG�mo)3|I���d]�R?�)�B�d����ԏ�t��x��=a�R�íT{#]jS�K���ߧ�^�R
�J&S��(�kkk���L�̚uB��,�fB��a��n���p�M��B�)���vU���0���6���6�b1�]c�5Yh����M���=��Q����E����Vb��v��`��SbhhMMn�̥ٳ"�����v&�5��<�5w���� xEAτfs��ԧaX��"͒Ȩ�ag�s6Ÿ�y����@R��_"v��!�3���"� �zg-��(�l[�U���޵|�}¢����-�����R���iTr�W��V�+1�W���`
���S:-��3WiI��-x�!��X�Z�:�P�
8e�)��hʨ-��rKUR��Ftچ�,�cՔ-�A-ԠȞ�nݺ\?�¤"dݚEhj�D�~����V�4�4�1�W�#8�rc}��7�4��r�H���\�f1W���%E��̠����d����Tn4��y�%#/_���=��glܷ�U�ڞ��2!�B����te�PQ#@e�y�e��n �#d\�n�i1�cR,y�.�a��fv�\r�ߒ[*L��vU[f��8\�&����`��2FBڔ6y���{(�Ĉ�˂��09WI?���3*���^�w�#�A���nf��%�����1���q�hM�]h[��uL�g�u��ls=7���]I�ұz����a����C������*�GF�M�1�Q�5��y�<��'
yY�_���]��g���h_T�ѱ0.t��=4"MU�f�y�C"�!�y;�c�� �1͸88"rŦK��uv]��NL�d<�d�����f}$��ԺKE�-E���L�f+�.�*dg�c�߽M"�k�tcA�@.-��Kddd������
�%�UUU7�U2�,H?ɉUM[d�DĖD0�%e�`]'���*j��-F��Z#��mԹ<��܊�k�l4�؅9� ]����-�p�b.p�~��n�h\Ѫ�*C\.���\��H�.�Ѵ���͉�IQ"���2	$��I>'�3�`
����I	̩���6j�̇k�����R�AH�ӭN��3�����>��M�%ש���p��2Cڍq��S3�A4&�o�&��B˸�ќ�5��hn�!9F�é�6Fg"����k%+r������˺�R��)DH����-YdS��+u�� d�xsA���Ţ6����=j��w���.!r��Z�x�"(f�L�Lee�/>BnX�m�$�g�h{,���t�հG�O���Ϫ������.�&�u�T�e`��@���.�S}\�I�P)���I���q/n;�5:�6f�.�N�ܴ��9�l�����Y:�%F�դ,flI ����y+D�0R6����FkNG77O3����T.�eɱ.�d7|n둭l@"�B���T�u�u��lB)���n�~�i��_h��Aa]l(]����X7����uFҁe�p���%��㴼]��RЀ�6��bj`�"�9[��9��ݐ~�S�RĦE}V�f�e��\�_�ط��{���Mi�_x��V� 0�1ku�er˗����{%4Bu�
���]�D�����XW�G��)5~G��Mչq���T�A��gwY�j�g��t��<�k��حX������d�zl�g-N?u����[R:�+=�ǲ���F̽�v�{*�2f�k��3Yݮ���i&V�vXu+�t6O��ƌ�@��mY̗����2:�,3��+5%Rx�?>-j[�f��(�x�l��\��F�5+��^�\�6�Gz�ZQ��cժ%p������.F��$�K��A�����t�Ȑ8v<�[߸'�s{���%�T�˂B�8<,ڹ5+jtfFG���ۅ@O@f��޸�H=�{&�j�Ѐ���DE{��N�w�9h1)F;Ge����-������{�O���H��9���{d���%0v��M[����������!���e�YKFWLQh�^	"J 8��D��q�����o%�I_�wu��!k�N����]g�u�ܙU}c��*��p3��a$�\�̒�������X��g�]��=�������z #G���~W�
3y�wނ��.�s���o*�T*��9��3e�?�G�7����>4oi66+���v��c�����ގ�g:��Ǟ��F��j<��j[O~�I�3L<M/uX#4c85��x�٫�v�kDX���aP�'����8�ĥ\椡TL���X��c���n�H��{p��4מ�(f��kf���h�ق��D��n���c�6b��n��woċ��Eab�V�͹I�7k�l��%��.HM�핸�O�ƕ׮��?�~Hikߺ��\�׾�|逰�������k���������­�s��r/����*�ٜsKR3�Q7�HO,0�R"�1`ړŘ��
(}�bp�����]��})yRT_�֪��jǪ�A��Bj$�h86���3#��B�[�9|~���}��t�=�(�^\c:�u��zN3|n8�0^�����?Ͼ.ﻌ'�I\=pё�ʥP�c��x �׾���7o�� w�m�������9�-s-�H������i͐7bӟ��0F'(�gn�y�9SV�ݼ�}�QAFJy�K4.Rή?ޅm����_?�#��q�G���(<ƺ��CYSz_�U�t���%�F��7�ws!��ji�"I�ڌE,��5w�64tf}����`_do�Y������*݇�q䟏`ۇ�a�۩�8����-�k�f��J�.,w�N�΅���D4PC��I�ֹ�p��
%V�Ĳ�\"�O�����EafDf��%�cʢ�lz�n:�V8#B0��?�"6��&4omF��::
�W��+89`��$�{���Lk�5�����k
i��D8����Ƙ0��}]���Ͱ��u#�#�
�[��S�VZ���-�$D�+)��3�� *�])�����%q2�>������q�6.Ċr��>%���A�&èn���3�kjYd	]�v���T�W`�}K���6��V�ܥQ���^�ss�[?�-�Z0��2H�:��C8���(�/ŝ�w|������eQ;����MƱ��E*�I�saY�VZ��,z����j����\�QP�}��#�<���*�y��whXW�G>��W6 N�俞����K4�]o^��~�v���/��s v�<C��[~�4mn��/T�>�1����z�<p���1
��S�.�9>L9���mN��:[����v�2ʧ��c�لU��noE��\x�V=�
��[��ϞU������Z��a6ͅ�OՊ*����s�ENE
w�0�-H��\��LC����Bb���me�ܧdE%�%���F�(����,���UY�Iڷ�"<Eh,<k����]��J��G�q�hJ�VY�ȓc�
t=��n	�Ԍ%���~�d�P���r���#R�wA&{�;nѶ:~�O��޼J�ܪ\\�[�VU$}����~]=�?�ޱ�eΆ�L2���6��F.�*�5ن.��a�br��H&�+�Q�K�f�f'���^2��eը����W^��>�4V�^���cX��둈&���������Q��2D� �c�#+q�����d-T[��AÂ����_��W,�@(ϽtC��^�5}Jܡ�R�`��˱�%z-!�����;T�ܢ��B$�R��W^����5Ɗ�\�Ĥ$*	|?s�����'��Nג�1c���Ԭ<{���	z��b�ʘ��/��=��{�u�^��/���q��Ǖu�-v�B�K��ꪉ�	���P�m?�W�/-�h?z%�����
eE���Ue�3dQ?��OT3�H��j|�w���>�Zi՛���|�JM�ӕ3#�r�A��5o]3������ut����˝G
׽3Ja?R��*=�u��H�P�E<��QDJҺ�W�Nu�(�����aQ�E��M���T����H\M�����˽�7��XGX��0�R]I�Sw���r�����CC:�M6h�m�k\e���sL�"%Ҡ�����	i��I!�I�[D��g�ml��<�S{�c��������f��^�K�A�fxC�/��q��Q�\[g����6���\��ܞV�6&5.wx`�U��V}����v�\����g�9;�u�W._���U�G�*��!�����(S�6�?�6���2�U��7�0V���)]�3��熻�m��O�HMA~19�T�����b��.��wQ?=	�8e�Ex�[Xh�����.��洬R�-���)�����b�k���s8�߃x2	oʁF�_'Yo6�P�u2pyHU��G�̵�D�nL)��f̶����.�LQ�l�������D0��}gy��uz�̖�5O�`u��a"E��;�駻���K���'�b��0l�I�����BO`D��4�	/��rCb�����FUM��`�.���B'B���DFsna}�d�A]�N�R=�T�%��т�F�J�m�ծF.���PD�c�����E�Ϝ0�eǰ�B�58���([Z��߼�[�Zt����Ջ��$��<~EGc�X��E��l�	����s�L�Hdt'ǕW/qTO�uz���6�xh�a|�{��X?N=u
�G{|B[*�Rg�_]���������H��@o ��X>p6��,K��g��ytb�K����u��^*��h��ߪ.������Y= gj(�&�es	s�fBdԉe��W���x&�i�Sw��,e����t7�>���8k�e��j������R�eRF��}x�CO���TkͪԮ�U���ȌDU���p���;�k_����.}�Vwz�b�F�m��Ƒ���iIZV4�ii]�|ȩ���96��Q�i�S�Y�Sv�#[b�oӻ7��=�ݣF)Q�V�y�:/�d�F&)����x��H���
R�鶷{�j��b��{юE\���#�E���������u�6b���j�Ӓ'eKt��IVcQ���>���X��J����:UX0<�`F��6d1�<��T�:'�ҁ4��p�2�R�W�󉳘�A��&�lUs6�a3څW/�F��?�eэ�	��؛-ԧ�i��I0R㒙D���&���_F�!���7��{�w�)��/;�`����R��|䕌�����jփ�Vo_��A��F#�Ƨ����;0�3:c
���䢂�*󱚋>o��n-��#=��us���h�}Ƞ�k�֌{>y/�B�t�t�>���}Xv�R��Q�lF͜�/З5u�N��j�53##�,�n�gּe�f�"�	dU�Z�@cRә��W󘾸�u�ה�nIƇx��p��Ӱ���aM��|��K�nn�Ȁv4��x���¢$��W��U\x�¼m��S��u��� u�Oݨx.� +k)C��梀��S��~�H����~u?Zw-��v��+[���a,RO4÷��n�2'���M4��@xRX�/�H^Ւ*�VIF�O3?؍���wfx΅�1\���~�AE�l�/���3�� ~���w!�ٹ[�]�%�[�o��,Q��ރ�/��s�ח�k��x��On�[�U��F�(�afȕ�W�*��H�R�̤��Rӈ$�c�ؼ��l�0��R8)��@���L��B6P�'�"�I�~� ���8�,_�E[Z�t{�h��mK�`��\n/_"m&�ɋ0Zwۇo�����OjN��^����K����yh��ԙT�%梐���f�ν��h������(���,R�;N(�IK��o�*��\�ATiM�Z��uye��c�G�����E��H�-R楲p��߳Y�ۂ}A<�gϫ���̾0����r3X���s}75���6ESX�^��BŠqC�����b����!�o��Խ�����_��i��T�6w?���y#�k�r;���<���
������~��ެA�t3����r�����әG�A�Z��\b�|�"�҈�<RY�귬F�����Q5ɲ�x�%��'wi�̙�Q�HJ�V�0���>~������q��}�x�6������t�"HiDs��&�w��4y�o�:k;sֲZ�����=��?�;;��vM�֜Pd�
�v�r��[AFղ*m���9`��k��,�
Iu��E{�~�k����^ɇR�3��g~��e�;7�qc#:�9/�p��ʱ��5��7����l�����¿�}�~<���q�'�5�x]B]Ób�E�����5f��Ր/�<X5�`*�R�ke��t���_:�nM[epIf!��;{-�D�e��̔��d5�Ed\�}	k߾�*p1{q^�s\�-��Ο��sx�GGP��HH+<��cp/)�ÿ}�ڪq��e��שe�w?��ǯ	lMZ K�W�J�7p�������l��ܥ�k-=(V�|@�:�;S�2�3:F3��4��ۙ�2�¬�Cm�ދ�y퍔Ì�t*���]�[Y�u���($m����a�
�b�|��{/����ZJ���$���-H��2LZv���vrY�/|��Φe�	g�w��ie]2����ܨ.v���5���K^���5(ѲԵ$+��hX\�ӃJ{%�+��fƳ�3o �2'�(_U��?�}���/9�1�0tvh^j��e���n$i��nd��-KnŖ�1;���a$c�LnX���x�i�*u�l�S����B�8�z+x��n3VKi�z$,���r�9!�����?���ÚX�R��B������邠��2�]����,a�$S���]��`.�����Ren2Sd�����~� �����#9|�sD٩ɞ���
�h(>ksgYbP�%8b�y�
Y�u�L�w���@���:WhQŦ�**= 4�Ư���o�b�u&g�>o��X&3��B�u��-��:ևo軸�EV��7�@��n�Ö���<�H�^�2�l�;7b�#�4s��K5F1xj��H1�a�I46�	�w����X�
c�i�����?�X)e����:��ny�-�B�(�v~t��C�T�S׏m�*{,GIu|�]8��<}�u�m�Q���^��A������q��ܵ��=x��j�5uzZ�̫��1���N�T�0_`QQ���uG+N~�$^�뗕Ps!�����}�>�t���բJ�t�S{�̠L$�SI r��������CrZ⃟�m���b�L`�.,�]3�5�[��/~����cl0��Yhj����jX��U��<�� -����^��Z�-lxl����������,c��kba�T�ItXFǍ%nd3Ժe��|
�^�F4�Ҁ���_3�	��͍����?^�3r� ]�T�磔�}�M�>)T����`��v�liƹg����{
������> ơ�z�If^;��=��c�x�C��|���l�6F�n�XS}&�^Li���L�i;{>��X�0�?Ԯ���9�����py[���*p�]=t���T�a�a�}�y��GuQg}[��%B3��e;\��뵋�g���+���u�i4����iS\~�
F��L3rn��bָS��9m,��HY'b�����uo[�j$jW<���[��jr�<�����l.��=�>�hR=�="k���O'��ƧZ�}�ʺ��FB���0<�m-h����:��.�u�tW�M��S=��c�����t�s/��v�qY�9�4�t$ֳ 4/˝G
_�>+:���EkZW�
���x�k�q��⫟f-�����$�,�g�f0r��]��n���"��j!Z��5�����5)n���t��^�ҍm�����v�t����t��B��߭�11�+�:_�T ��U������˩a=���ϱ-�cu`(Bgr��<R8P����6�;���Hd�7�B�2��|� E�ȣ��|�X���#�Gt�:��]B��������~?󈮽\�����ϱ�y�6,�Ԇ��
:O^�!\L�ϣ��.��t��x�п9�sn�Љ��21�̎��
�|�RC�K���p�kA󞥝PO���s���K��Q����;(�se�J��"��a�F��3�Z!s����v��swg~/���ϗ���װg��FVW��IM�>���=�c?��TR�u>�a��y��^t�B A̚F�m��i+\2�X�;�t4�#�Ld��#5��'��p��lB�Lv��&��%�P$��{�Q��O����?.��:]��]p����=�C�q�{Fڌ��3�؍��z���%_|Nw�X���of*����vS�4�v/�{�U[�x�����e�p�L9��@erg��L�0�#eO�V��r���XCQ�i�z4cH��([�|=uS��x"���KsGӁT�d\����+B��L d�a��2���pD�px�f��u}	�˽룩��$�c�����GB}2���o?�TC���Yw��_U�B�'�P�sتK���pւ�u���9{��00&G_M��oO�a�K7�а�	�g�U��n����vPEQ��'�4PN�7����H�%�M���Mm���L�#ӆ�����G���,�	��0��!gk8��k�r���
�'P �Ƃ�;=�)Y��Eqz�Y�y4����83�}jTS���^����FEU�ඇ�Ѷޭԑ����ؖl��m���ǰ�� B#	d<��v�e"cƄ���Rq��[�Mj���X�Sۿ04�O��G�{�X��W3�,J+���pټ����<UJ�Ő���d������'\S�੠��n+�m�&C�Q8WM�[����p�;�Q�ĩ��������g��~��c���Y�C�q��S:���ܱ�Ǝ;��Ϥ�˃�z��Zꨁ�:��\.���ڱ���h\�W�/}}]C#p�k�[�XW��r9>������S��X/~�!�}I��Տ:��<�<a'O�Er��
+��ǳo{�_;M	onr��΄ѝS��[8�����i�%i?6�O��L�pe��Q1�[���η�㧂���8�]U:��>��j�d�g>��5�x83i���<�[��ͫdf�;��fu�� N��C Ci�+��b��z��	8��E�[~��_��zBN��%����l�ϭ�������]��U;3([�56�_@�+���υHGu��U����~g�h�-~817�/��}�;��Фӿ���ܱ,���cc�`������;A/�Ճ��xB6��n������3{#HD�8�䫣B��ټda�{���x$�a �c$���z���N��]!���FQݚƶv����~�t�>jj��UP�4���3��[7���K�,^Y�H�/�ر�RP��6+���>yq�"1�N�'O(���,�Y�|=�s���~�)�0.j��Tu��2~�y�T,�*β,�v=��۱���q\�2��bE��d� *&��1�AWw �ZBhj�G�J'U�v��1��HU�Ks���,j�!��V�e��]�<��9e�`����+'��n]Vc#�]�����J��:�{�g8��w�5o�S �q����<�Ƽ��Ȟ�D��XC�B�/�������PKUiF�4���˹���Rfb��ڽ��?���ؓ��b�]�7>f��
�,��x���n͟!����n:�����&>O+�������C�N����ܣ���y�0�H:IG�u�_�.��R7>�m����NУ����pe�~�$Obt<�o�3��t�t��Χ�����=��,$�Đ-�!S����@璱��CM.��,��L\e1f�Bۧ0����1�\�LR����?+B��%f�V��U%�����zE���b�Y}��̇�+�P�����.����R�4���m2<�3�K�����Dς5c�϶=~�Tl�ln�,s�nt��"��x�;���	,Z���{ik�Sa�� �l��qVTU��xQM^գ�0ԙ�hO2����l_���7����q�ۿ&�� ��}5`L�e��fx�^tv���n;��W���2�b_���&{�N�������'B�:����z:�?c�]%yl��K�k���US�Fc����=�'���L��_�_�}"$���<�頲��wx�5�J�'tl�:��*|䙠:'g=��Ok��%�§�{Ǜ)x�?P��]%��7�\a*��\�'v���!��|��l�����/J}x�NIi$��g�h\�B�b'�������4z�%�s.��F�'�u!�/۟T!t}\�*�K�vJ�ӂ尐\d����7,��<w֗�e�,�R�ԲNJ�M�_�q6z�bd?|��thva[@F�/���ƾ_��R���`��    IEND�B`�PK
     uK\��92\ 2\ /   images/7fb2f62e-2fb5-47b1-9980-8ec272392bae.png�PNG

   IHDR   �  �   b�y   	pHYs     ��  ��IDATx���ُ%�y'v�X�{Vf���f�I6I�6j`I"4ek`�2X�l�������c0�����`H͈"E�l���ڲ�\*3��9��72���	4nߺyo�Y�����s�J9e���TB)��p�)�}�3��	��ZI�7N(�,}?B��%|����~x��f��O�����ͥ�R4N�P!�҆����	��/�;�Q:�z�}�����!L�Y�������=Z��
��st�|\)p����E����"\�2k�V���I�_�%��(�@�͠2�w.>,0-8wD�b<��)�[Bj��1�~ï<�kx ����c�WvS�S6�i�aM�]hO�]x�xi-l��ց��}�<�ϗֶ���X�Z_p�_��e���=�B)<�?�	�Uj�u�>��(��J��	R��5P-=F�-���y^nr��5ͫ&'^ MW�O)%.�us����Y� sI~��=��_5�t��o�-N���"
�z��9=Q|��YX���z�_���č�&����m��,��Pp�Dd=7����������%z~���[Ȯ0QC���W𝑣0t��<6�oY����%(+������u0���W���p_��$O`��q�j;z:�\�ȸJ�5��%Nn�S^-שּׁ��j�p��#�VL�[�W��A	���U������#�6N����60~�2����"��R��\�)�<��[��c<�P��\�(�s_�@�2#EZG�R'l/�	3�$Z�9����,KJW�,z^p��iŗ~�r��(HN:�CRz�c��8$���� ���fSQ���܅�-�!<z�O�0�tC�&.�/��V��vYKK�L^��IVt00Sk� n4	��c^il�3�+Ȉ\�B�(������I�����磲�@K���(�p�D�(,�u�*�¡�e�1$�t	��_I��lq��<I�yq�J�6��ҫ������x:�á��}�s>�o�7m]]�2}L�U��@E��)޵"W[�?A�w��]���j7���������M���|]��.r��A^�P{0ZG����Ě�p��- ���+/`�[��/T�Ox����q3}#��R���Iw���}IB�
7��,�pi,j��F�
�!�5�d���%����ȁH�����`�F#5��R�^�p+�������s#?��EΡ9�(��j
��<	�c}����.P�W�"|JQ��R_��>�XhL9�W8���:��������L"����$ p���@4�
MiR����@�4l+�^a��cxz��[__w���p����gZ�P ��`�}�~��m��JZ�ʨ/T���������t�R�� �"�E9Ȭ^�I��ተ����)>oY.��'��1<���uI}$��P)LM�(�`EA&c�n\^��|ɉ��^
�8�Һ���хV��yʋ��L�F����i�Z3_хB��Tn���	߁�I�̶��n�kI".=\;Ct�����dyJ�\j	�9K�F?���������: �������V���ղA#�a�Ke�-�&ն�
w��|�n��Z�E�O?�>�D�9�<�W�*$"r3�$^"��*|Ңo�C�Q�Y�հ@�a3O����!R< 京X,v���П<*<E�TC|�ym����t�CK�\,�`�8~�L��_#V���Nk/ �F�5額]������'�`_����*6>|!�.�e�"O��wI�ţ+Z�U%�(P��$�X��e��\A��\��-^�*uӚUC"��sC��!��mC�LjHv�N �ob��q�mN|��\��}V$��O���ۖ�,F�z����x#�L@��x�V�VH�y�7j.�CK���U�Q�vW��e������:O�{��l���sTb��q�jׂ�nH�I��dLZG���;_&����{�ĭ	�7��Hp.q���H'�;d��_� Dn����p�,.ې<\� F�Ol>�3}+u�|,[8^��-K�6`��f����_C�],P.�Cx�X �`��^��g΂2�����d29�x�i�$;��
�WN��e�
�NY
�0�TEZ�Lv8b$x����Rm�1�h�!s׸��<O���?��0a��Z��[�0�-�+`�s��(� ; ˢ(v�\.��ȤI@�7����YH��Ȋc�͍���K!E�����R�Ks�,-������񫝣,\�X@ {���H'���Y��3�w�ច�b0���l9;/Q��R3���$�F�ǒE v�z¢m�>�m����o�)��!��~:���}��6׎�K\�b	�π��i�Tˎ������R^1aCy����L/J6�0����ʆ�����K%#�� ?+FxܚAy�]v�~?�ǈ��(�eIґ�`���oI��D��$k	w�9�4?7Պ�:yd�τq�1mdҾ�5�EGJ�Zɑ���:4���C�׃׃�'���y���9p�z��uk�����d��ʢ��i�� mCcn�7H�Z[���;ٿ��ðL�ǉ=6g�QN���]yI �y��ݧ�b~2��!��ST3� ��<OOf!����$Sd����������fg����ng�
T�����ɉT����<6������ɳg�������A���~��Ķ��$��)+u��U�[�|� O@��n���L������&�����=O`�E貮G�m�XL,��</��I����'66�U�P����U�K�wu����'���R�z�7M���R~q&�0���B�Ǐ�H%!���L��y|v��l��[[�[��|6{~���Nt;Z�suI#����򡲕]%X\ �j�lF@zV-�6�JѨ,��O�����W/#���k�=m�m�7;ϟ?O��ը�赒Q/�v����s�E,;~r�4�}����;C"\��T^�{�`6�=<y
����5ž��L=}��7F�Q�����4��T"G;�T��Щ�>W��q�/�z�^��侠�W�j}_���ک�b����x����f�ޓ�(���X��@�G^mka-la< �GR
�g��X�O�
]$/�x%��J7������qY�m~~~z�BsЕ�L�"��˨�o���y�R�_�v���!�^����I35�ڃ֎�7�����ĥW��
P,�����W���ϓ
t�^g�Ɇ��$;�=B��PZ��O�v�Q��}�? ���	�KO��+ ?�'N�,q�^)T6ސ���W�-o�.k��h�j���`���Y���Cߢ��w�Y?GT�ʾ�Ue�MԚ�0��q:��k��$�,�{t��n�x ka�8Z�%�p	-� ��@������k�[��J���nj����Jw��d4�c�J fM�1j�%/t <�k��S�B�s�M�ۖ�ۜ�SՖ	��x�t�Ђ� ۋܺ�!!��]���e��2+���t��Q,}@��(���+�t��<�qo��6;��LV�<;[v��f&�,\�W�#δ��%�b�z�>�SX����r�e6Y��] �	#�b������V�)>�{��9���X�{�q�>y�XL�,��ò�,����j�f7_�S).�tB���(j�fo�b}���*���K)����{m���[�/LO_ݼzzz:99'T��$��j�;�������5�f���ڟ\�%d���^B����dOH��*�@��9�G��Υ�mF��Շ��˟�������g�\\�K��4z�� ���s�f����{5� �a�a���@�NNNA��7�5QآA�핬Wo�X#Q�Er|�����O�%Xϑy���h���z������bh�ҊW[!ז��u	��W\mꯠ�l��詌"�Iזh���ցԞc�VV� �t�2������j��]]�7��,�r	�ѩ��"�&yEV���E�n��^��r v"z���L�E��WnX��d1��4�-X��P�����emPlS|�T:H$��b�U39�!0�*D�+�;�f�F�K���b�<`S�Px�59��?x�d��/l�gi��-O�������GA�����y� �:�M����GZ����)D�8��v�##%�t��� G/A
dvg�1�ã��d	�?,}dב�ݵ�{��0>���@���Ҵ>4f�艑��]�Ţ���c5e�CP��Z��i;�ڗțW��U�^-�s֜D�U<��Ÿ�VY1HzF��GQ�����UT�d���HD' c�6�l���=}~�P��i�#�7B�8���cb%�Vb��x�%_�8��D�J�Y��\c���]Ԧz3qF)<b^5��L�^{K(ϩ�hfsiv�����8qAM�K]�z�����Ǐg�c�e��>�R�� `����b�"�gUm���V���*�J�"��2#p7gr{��A�u�N*q�	����E�q������}��U�]��~��bg�h�X��N����_�Qw�����]pU��� Ok�z*32�*G;9����e,|����ٚ��Ⱦ�lO��Fcm��M��O�q�<�܇��n#�:+F��j����� ^�Δ������]��Җ���I��S���˲�����R���چ|ZR
�a�ɮ Ic2R�9nX���QP�%����E"�]���6���G,�L����)�F_��(���Ȍ�߻q��EQ����s��nG;��@���2I3��5A����%���ʱ\'�6(0�gaQ�K��4[L�;�ۓ����ՎƸ�+�%���lZz+�}�`��@���y.����n3�V~dT�!���-GTh1�{*ے��$�O�u�'l��}��2U��u�vH�j��?�Iϵ�6��Eo�� 0�&����%�omm-�$M�� `�9 `�\b���/��+_�ݗ
�WIqN��cA���޽{(�O:Y�x-	��D����~�LQtS��=�Gm�Pbl|��`D�䈃͂ +V�'*�~s���U��J��3��N�$`̓�#��6n��Ĉ;->H�+1f�`dz^Y��Z	�ls�**��!^�Ӂ��"<��ĘB�0pd���<|�t�^�\���hĴ�C�|�f��Fg������%�-�.V���;�֭��/yx�0=��"�eyna� �aM#�x�OaJfm8 �\.�~m�)��)P�u�j�\[�
�]�%|�r���[�x�F_���N�U�N{�&A��"���F�(?ZF�[���	RC� ��ӳ,�*o||v�yY��;��q)J���]aY�qY�@[kS����7�+���������K;���m1��<L�HL��3�G�*�I�A�I��Ol�4k���°@C����� ��ho{�]	�:��̐m��o�<�e��e��lY��Btdg��vg�|^�qf�=9|��.}v�tԁ��Ɂ
�H/���A�Ӛ�f����,�����*~NQL�cg���W��<j�MZ��;u��i��d,��r�ʨTdf���L)g�C܌`v��{{{�O[㺽�����rІ�!Ht��߿��X�.��f$W�a�3^���P�+8��R��Q
�:��o�����kg%Rg'��;b	�E���@�O�X�`>*%��:��p$�1�ۍ�w���E�	&��,G=�,���u�z�z�h�!g�E)+HU��	}L78~~#,G|RR~���!m�C��-�c�|�k�o�F��?�R�����E�2���D����!����ݻwa߁�� ৩�%�
�I�ڻ�rm���GH�.)W�7Y�a���r	�k�ϊZ܋���N[EvD�U�=� ǸX�`�)J�Қ�,��c�~���-������c���4���Iz���!rf����u/�;���֌/з�&�[�X"�ߍ�2���E��1�~?�y�B�gs�M�%6�O���AK4gXL�|M�����R��4YN&v2�f�Ȣ�)��B��'kk><��ֵ�����+j	=��"�A�ϛ�Sf�Mt #/�.KD1��G���a~|>9��}����(�L�b��VE���^���@�ʬ$�hUi�aNV��
h`��	t����<;?���~��W����<�bpm�����<88 ��=���]x炽od`i~��B�
���/Z>��#�iit�MI�@L�(鬺eIH�V�Tկ8��휊��ƃ�1�օQ����[(P�<x� �]9J�0G��K�f�8��6	3��7�UD���s��W�o�r��*܆N�0%�����6(�H�zA���$�F��[$ִ�
J���z���/��W���n�������I8� d�:�爵Șv"
oN��89��F�t���h$�b�ppI� ��۷o� 슳d���X_��]�Z��?��������O�=z��}�Ir4e�>}��A`n޼	 U���@�h��*��<�����.��*�Z��L��\+�ν`�]���Uv(0��ΈP���۩�@����QF���)���<3�]B�͐�,��xs�z0Oڗ�U��|���K=͔0�\�-��;���4{���?|���r>��no��Rg��(N��x:N��4�����qN
z�� 8-��{��..X�1cɺ羁���*�4�MJ�����/��%��!����������SWd)��n����x>}VΧ�+|䓣l��'��wF���Iq~>��c��s�`�]��s��Y>�x�W�1�����89��Y����0��J�EZLOO����X�18iaT�2R��(*�}����U�I�oRP*�()�RTB�&��"�,s�ա�6�W��%�/��{L쥩
dtm�W��D�wP,��G)���UD�.�D���
9]������||i�� �Lu� ��4�ڀ�����Y�3 '�����[ϒ�g����=���n�<�;�l6X%W�/g V��!��>�]L����uх�iD��c�9@6M���yNE!��0�?��7�0�u��
-�8�U��C��߭���\Vu}h���$9I+V� ���q���<e�}�j	ں|�~V��w�W-7��*W.��O����u�\m��W��5��K�����(k��23�gE�ɯ<!t_ hS2ĺ��$0�p�D�R/j2��-��J��\��ySl߇��G�h���i�c��{}����+��d��t���b|tH�p���\�o�2�d�1��9����!���}�;���GG�'�G@�xћ�!m� ���;w�[�i�!?Rׇ�*A^6�v�'�+(���()@���ޚ��M'��&'���f&)�v�bV<���Ngm/^+�[�'��0��N�aʐtB�3ñF��/@e�~#��\D*��]��O��3d��{���z��ƕm�\e���4%���Ԃ*Z�44emJz�����3!uΛ`�V:YR<�4��*Y΢Ըfc�T�bIڃ/��*D���o�J�S�ǫ��U�
���<l�r1��T}�������Qu������:���^�'��Z��'c����֭[�<��'g>�FI��������S��q|�ٛ�or��l0�9'�b�&�8)��l��5	7��cB�M�2��	gGK@ϓc���J�̢~Hz9� �����)h�K>��̲k׮�<@6�=1�������X� -�N��]__���p&g�sn�$|̑���)�c�~G����ؒt��]x?~�Sx���#�����K�F'�](�h��@���JN��pu���i�l�7\�½�w����,�W6O��z "ժ�����+�h.ϕnm�V���O����F���`!��P�"۟!G����8���e&-OwW��o��d��6�_{�6s��F�?5?o�}��X�����{�ko|���g�Y�#NNO�6̀��"���5o�3�����w��^o���0�0ϻ2lF��i�Ɩ�<J�t�õ�v����~w6��w����O`��s��Q������PP~��(`��a��_�'��kU9Ɨn��@����7d_?K�I��#-' �<���B,�Iw���c����s���Q`�������2�9>J�H�y|��>X���/z�_�`m�-jC�]��;'�U���<r���!����:&mi}�*b��5h�{�q�w�e8�K6�Ć.�W�L�cuO��\ ��yUYV^�Gy��ۦ.]���������ʠ�z��vt��3��e��JJ�����)�Pd��Զb��\�$������oCf���6�u��Q5.J��7o���kc�`���6�=9(}����)�Ih�Y�"#i	eq������`!��0�7nd� 4<���?|�]�,����;��3�pz#�����lgA���x`����~������`0����o~���2膰�=�{���۷^�1�y���~�|��Δ� ���y�<?�7��h�B}����?9>>��w>?���o�
�Q���F���1����eli�i��p�l����p�ᅔφr/�Z�U�m�U�\��ɷEډd���E�t�b���<*�����lH�JK�-BZ��w�{J���\?.��b~8���c=�Y��MpUW$x0�"s�==x�ٱ�~�z�6��X���o����/\2��M�J�H��Et:����1̑b��h��!;��X�e�@�^�-�U�,[�ESD���p05�����>����}y2���W��a� os��?>>;�����+h�d�6p+�c.�||B$KBAE��a(Jq�������Q"�������G?�я��⍍;w޸������Z.��|2~�dmO꣋�O�%p�@TI�|�%-�H��u=/�r[_|�M�V��[���kkkŭ���8���,\�b���Z�>�u�iI��w^�[U$�Xz8���I�vS����K*m��u�l��aY�F���op��5�i�|�#i+W�gKy��T��a<�ԒTV�;`�F�sк?:��E����Kh^�.hXS� R�^~e�1�ϭ�y�Q�i�����@���W�kRX�X�RY,��Vo�կ~���, e�U�]2�_���K�D�0�b�����60h ��Kt� tZ������
�L���v u���b!#�~����������۠%�2�	�.�vZ��������'K���*���%�2��[�K	e{�9J�4Ka���;�z��O������9�G=�9���^��ے�iHGަ�Ko.�f~#.Ti�W�Vnz�d���z�u��*�RU�V[ �K��8���y�o�Fhϒ����h�SP��F��5H�o����j�V�c�T�O�U�����D��+�'3l.s[����dǋi>���Z�����w���������t���~p~/����b=u)�I4m����% ��ӟ~}��ۧ��l�q������AQdo����+ׇ����~�3�y������0Y��)�s�g�X�����9a{�p5y��ý��P��?���(������g�@���X_-��.�����J����nlOÖj_Ol��1��q��7_?==������B\h��@~�y��ņ�/�G�pv{Kڪ�N���N"�i(E�(j�<ʆd�j$:P�Ԭ�Z����7�2)ǅr+��44��-V�� �-�3�V]�|�ʹ��ר�\��)l�T����Y����$�m�U��F^�~�~h�/E�%l�r����cz�����>�?�ح��Ç@ �@(>����R 2ưTƱ<���W�L��+�F���fg�ʕ+�����=���βw�}���c�-�� )�^�Z������M!Y�=�{OS��cC��|�K���h��~��ܵ~�=k���� Dy����Q���S<�m�]���)8��U�Q$�],k1}����G�-����9��Ǒ�w��O�G�ȓ �R�0*�>+���h�l/�G.�H�ь��*Ͼ�ܯ���eڹ�Z՚]���.ǀ։�7��c��Mv�!Sh娴Eeed�>[���?\�%"/��zIF����m�A��P�W��i��N���E?vE��E�-+��=�.d"��;�iM�I F�[��ܝ�>��F?~��Ɂ��8��t'ܾ����wvВ^�+�L��(K�-����C��ͽ"�:��}�ڳ�{0��̳��d��=-�>�&xw��������u�<_]�Iz0xA1�*<N�5~e��5��䍍�۟���+o�|'��kõ�t��`����H�����������~�S����\�SJ I��Qz�%��|df5qa�/'r��;������?�Y���mo�f���w�ڧ���Cq�ܞb�\枅����a��G��zz��SeS�Q U�K�Ùz���V�#�h~�xآ~U�nw�	�{b&:Qk�M�����$����?LU+K�U%��K�5�2�j�F�xL.�dt��u�;��%[7U�Y�m5�]��b��ɱ�+����M��W��]����e�v��1� ք����$�&ΰ8�3�����)��M�H��!�H}閰�V���d�'�&�T.� 2�㑔�e�<��u6�nY)d��i]l<��~��Q?z�7xHX�����[��L� ?8x��1b�$S�+�׈��2�t�=��� w�	��̞?G9}|s�۹�g�à. x�|�����(p���eVM�DmI�KV���ٮ�N���߶��/Wߴ�l\�9 /^�R˩3��8_L���r۾n/|�g��y)]��X�n:^ qfW�O�L�Ƌ����� �D���#D��7�z�P���؋T2n)5!"��IZKr\��\r�C�D��;���jH*�pä�O�0nߔ����<��9ڶ�������Vro�0���f|��L"qF��"���fL8A�w�g$���	&�D�sml,�����<;���q#12DQ�G*^�����8�
�f�� 
R��P�����3��&ܢ��e��Cu�g�dz��ã�q7����G�)p�O��zz�_�޿y�Y�{�c�z�I7�̹KLv-kq�踞!��$Ĥ��Qq2?|4�������|nGۣ�p{:I7�k��^�;� ?8:�D ��/AÎ�!�r��π
�}GYbU�*��P��a�ʭA��2L3��x���5�$�=�+��"�
��tL�gE��ӍO=��������%�����e
Z�j��b���'ʹ��p�^.%�#���� ��� ��:�9��˯(Ms�|��x�U��bΘ�g���p�n�r4�����jh����hɉ�/����Cv2k������6�6��a�Z���>{������6����r�6[~�']E.*$tP������+�ruF@�������!w|,��V��s[��V���)9�GmAE���b�[��B��~��]J)��Aw4�H�l��v�8�sss��]�Ó���޺����>��A���C��Qv��H�B�J&_�A�h��\�<,��&�d�ݰl@J.��~^X�U�HB���8#��$q�"�!���%u�b�CY�<����7+#��(F+�$��=�
2C�Î�QW�qH��,94]�حw���'ʮ^�!�¦6@��:S H8�'��.A|G���c���0'�kf������6���$%��J1������lauGG2�,����xr~�z������zX�����V�9NU}�OY�U%�o�@/+�"��)n�qq��#�c�F��A����q6�e,SZd7��G	X�[�V=�D� �&$腖���؝�3 �����|,b1>?���X�}�J�����
_���دƖ�X!+^=C���H[#k߉A_��^�~{��;��$S�e���9>�B_�I�IW-���`g�[@�>�6^�!��,`(҂;�(�!eDe�3��l����5ʻ�"�����8���
�PJ�O���$��F�Q>=�<��ƨ����^d�t�b�B��}5��?{t�i�[�{D l�#���t���H�9X�!֤@OJ�@(��Ė��{��M=r⬲��)�E��S��W�"����b9f�[,:�LЇ �
���U�qWeԈFҸ��6�������g0�;�Z/F/C6���"���U�ϝ�qv���2�x�y1�3	�@9|r�<��\_m�D��!R��E��F��[c��R9VS@�ơ_�������I2_M�����h�cu��H�:���Wx�߶���fک���q����hy3���D��f"��bUJN9�*�j �kήi���j,�+S�����9I�W��X�dM��"���ƥ���8V>\l��e���6� ��[O�﫫���A}�����Y��7�\$�͞�4/����~sM�ԙ���Pd��t8���$(ץ���h`0�6�q���M�����AjҤD���X�%���y;� �`�E��I%T Ϯ��}��!�.�o��}{z6�!�9|.�w0F�ɪ^��@�^a���dz�P�mA}7a]��L��MY�"rZ�,�M��F{{o� &|�8j��㏒,7v���z���s'�r��A	z�� }�����*hʠ����q�A�bs6ým�^�'`"���'����>}:�S����<	�2vˎ,|;�99"e�J�[q�ft%�)M���B����Q�����=�v�,t��QX$J�U���0���q�f��^P�����L��g�����B��A�r0 q�7u����'���5�b�`�\�-$�$��G��bR�'�ˎUϢZ���dOv���Q��=����5z���%�z�R�{/D�)tB�v�
]�2jp�,w�'oM�	[O&vh��mc��{���]lֲ�-�k׮��	�9]�R�J<�"Җd�"7D��ɓ'�Y�{qX3G|OЍ}J��?�裱�P^Z��}ѯegb��q�6`;dF���k�n�;��t��[[[7oބ�;�\�lu�u!�0q�ѪgPu6�%K1��	}\�+��\ē�y`WV˨EMNI�]Qwpo�9���zL�UO�-%;c�c��!��D���w�rۉG@=�6�	�#(-z�"��Ү�tI%��z�s�Yl�t;E��Ʀ��b�|�}]'�����3 �����^9�@Oh@ ��A���(���] ��^�_�X��u�twׯbs[��8N)>X��oy�����ϱ��,�a��9Z��Գ������l�+�(�����x��f�efOO��1�Fܿ�u����,��?Q��|�Oታ�W��C�J�_P�PH�m���w1L��|��#�Q=�%������|^����TG#}��#��Э�d�	+܌B�Y����!������d9~��E`�^����N��`l�Q%r�`�H���@�p�qɹ@d� z��P�T�\>:?S���`3�SX�PeV-��q�IX�����/m`�4�!�Eުi�0�t��w'�X�Qb5�f��F�Ѵ��+y��7�7:<U�1vaΓ9��������~���3�tO��΀�]q����$iK�Mؽ9�>Y�X��Q[�H�i���,)W$�U_M��s��wn�.ȼ�ݭ��큿�=��'����9��ߺ؛,'��/
��tJ��W�0;��6�ê\6&���Pr��R��}���P�~���p�c�����]a,��hZ��&��29%D�P�6�����\���&���,U��V~o�ʽYRX�G���+�|K�o$`��q��讃�5C�(�B}c�"A D�ϝ�^����P�>Lx�<(HPy!X�b�7)�{���]��=�p+�[OC4Q��AhW��B���`cc���ȝ��?�� ��@�e��{���7D9_��#)��jcj��:M�S%/��/1��Xa�0�,9� U>`�(mBG�hL��4��Y�T�h��P__���/G��k�7��F�ٱ�#P_5�tڗ�l#��!U�ۍW7G��򓳟,��E���3s��}摙塡V��Re�Z����"x��;�ц��i/�brt���Jdu�el���AvÍ�7DP-h3�x��R�J�����n��(Փ!��������P*�V��ĺ9��7Q��'t	����!��_�#�J�j�J^rE�T��C0Γ����
����f@�c`���|7�;E�y�+Ư d0�O���Di�*ڨ�ᨔ!{Z#�~��p�Q�� ��:j07s,_ȱ��9��H�`LQ~A�����QDB/m���dcR�Ec�dZ\��>S�~ow��6~g�Ƶ�k7F[�k�q�4�vq�����SVdq�������Vrp����?9�)�����2UK��.!�|ȯb��(� XX�J� ��2X��Ƕ��j�'�YIY�~=q����9�	�}��Q����oUݿ�j�N5���Ԡ�`&���4H��I+���,`�xI?i{p�A�np�@�Ir$����Ԫ:���ְʘ\\������؋�@43����kAy�VS�,�2(d\�g�2ZPD`1����:�Vj\���H�2}�9v��1�9�9������I%ʜ�d#�Gf�OZc%��Pa�d��ޒ���e'���FG��^\�%�vK`�b~Z�!�K1��+]��Ή��OҝƟ�����0r>�*��7y��	��G��j�x��������_���om�]��sH�M�n�)�}�a~�Χ࿍��>��$ؾ�G;4�HU�=���r�Uo�GB�4\���کL�M4㬣�^��d�䑡c�r���W�/������ʛ�ۛ�M������!"�R�F����')��+�(B�1z}s��I(��J���<���^��z�����)z����+W��������Ük��U���g�th�#���;�B_c��� ӣ$7���}s=�s��S��h���u���*	�Ly�9��s�>>EQ�C# �3kxw�Sd�&��P�
���Q���~8w�dר��'��A�*���yr>W|ڱ��T��G=����"b��C��tFHߤ3-�L���������"(�=���/�1�x�E6���Z���&�I~��޸�Ʈ7�S�5t����h�a��}��ԕ����?�~m�������a�1#)�q�V�`��ޒ3���A���.fQ����]�wEp�%lއ��6��]�{��UP@�=hra����>�s�v�����*�6f}}��ݻ���:��3��ĕ��D����^�9�@.S� !�(�b�N��A�j� ��H:�/G)>�!N%���W�<�ڭx5�1��ϋ%fES����I�8a$���c�M�P���5�6�Y(|�,����L�� �KC�ӱS()E�\�l ���:;�d��Mh��E=�6�6�+�'�P�C�uO��|3#ǘ�8��c��y����}b]38F�#
�i4򩂥{��>u�S�h`�:W�	=R����4Ru"��a6Y��W������{��Ȋ�����OE��o��޸IX4�N.l��L4|P�$
M�2
U�-`��2 eqCmn��w7^[�+��*$�Z,����*�O�|~㥋KE��J!��Q!om���N�2)�=����pc�vt̏t�4�Z*7eVbG�|�<CG�2���O��T��M �A9�Q��}��!���8�z���o�?3��N}�D[~f1��i}1u%��#|���i�Gf���y�W�;�o��!�����%�d�S����b�+RQ�H�����(RP�WԱ���>ANgѷ#��3��oM��Cs���)NxNoV ��ɴ��M��Ǳ-B>��#�p��� 9R����77����d�*/������n�s�����e-y!,�!��v5�����yk��'e�߂@Sys��+����=���?}��j'�7��,w�og�Aw�9���&/�W�����R��а���w�߷߮�b�X�'Xo�M<�\:>��r�Ⱥ���neepx�bb��QO�o�w�Ǐ�O�<�C#w�-��	�E�,V�@,���R�-y��T7ꊳ�����Cd`xlS"�p>�����!|��4&��=y�@�wD�"���G65nu:'�S��䨪^��	��e,Xo8)���Qn`@2��J�f9���|�f:o|5���Zp�f�19:� �$ꐑ���z�TW&�F�h��sIIi*�B@4--�g�d �S��L+ꅽ;w�ܼqs�����p��hE�j�����/ج'�x2��B�Fk�o����l���#��چV+\c�4ٚ��l�Uy)ê,�+���J����鍛��[��a��x����I>����8����ִ�S˝'�wGV�8��D��S�7�����YG&�� �&H:�{B�=Ġ�?՝����G�WL��N� ���E�d rƣ�[��hXЩ�OlB�� dh��H�e���C;l�L�,_쒮;�Ǉ�ґ֎�|]J�134^5g�r7N���70"X����nC��.��8<�)7[:#� �yn��, ��"%���dD�H�|�k�=2ɘ�JQ��/aU|/�1r�H��h���,p�ع�M�I �q%-��P"
��鬜���vrz�-�У`��s������{s�
nzbC� u*kV��e�D���t��0��C�|v�&S׆W�k*�-��@N�8�&+ݒgM��}���wA>_�_��+������-kk�M���G�,��F��U+[:�^�~Y��!qt����q䁥fdE�d+~�ʍ�>��D�U#%a�-Hq&��Η9lg���$H��\:_ j��U�O�s��cB�^���=EVrZ�^��K%�ů0v�z̱!ؾ,g�ed獳�|>g���Ka�}�|W��'P
�ȉ]�-y�a�^��\X<�ڒ%�ݭdU�M�#;�Cv�Zɖ'���Y���t�����Ä�������)y����eUt@��UA���!��;�8�!��l 2�M�B�P�HK��/.�T��(Q9��,�9�k(�o�QD�@
�r��>��g�o1�k�G��B���$8� �,�n֒H ��a����S�b�]�2.f��-����{m��Vo�"��=�-�:��}�-W�+����+psO���C�S�H����GGǓd:���c�et趷k����%��e&�����B�X���f`����x<�2��^A�᩾�g���O� �`ٗ��в�#��pi�R� �K����O�i>�b����Bo�C��qfG�1�r�͍��������1G׀�o��Pޗ���� z
�Ͳ�(zT�d<]�x��ؠ��:�����d2YL&���1'�{u�P����<�f�{��Wg���"���
)U�K�G�L���!Rڑ��_��y��G���7����đ,��w0�.N�N�z.� rmF�}�BJ�D�B.��v<�F��0���6�����+kvġt�d~��L$*���ū�^t
������s��4�^��W������c��e��{�\�����@��u��4)g�i/�3�����8	-j�2Òot{�F�yҾd�� �+��/��Ad�#�vw�Q�Fϰ���K
��ڱ������a�c���l�����c�E�����ɒ��N�瘉�{;;;�0@U���|���h���C��ggg~��c��01�=b0�����7�׀���x:����`��JG~�����?>�Wс�=?z�������S�`)���> 0��1h0�KqR�ԙ���`ˇ4݈��N�����>x�`/a��f���S�����]n����	�w%�V6lqV�O~��()��0l\h8,^���q��\��#�˾��w�~�}8�)'��a�/
���ȱ.W�m)��V+�ӷX8����Q��>�RS3��$���&L���� ��+F���h���3`I�OI<_=3iY�C���%	���iZqk�,��O&3�Y� Jݹ}��ի�a���7ۜ����n��YfŢ �>�t�����jXx�)��ܷ?�}��Ϧ�l�������m�z��6�]�ȇ����릓>8x��_�қ�`Y`��`!��
�� 2`,�i~�����ݰ���3���C1)F��1��c�#���G�>_�r8=7o޴~�3���ED�0�xt\8����7,H�h/�6{o�?)�����[�lt��7 ���V#J
q*�Vsw�s�g�t�kx,e��w�B���g�Q�d�t��_��]����?�i������H�>��*�=tE~p}����>�:1h��ʹ�N��m�n��1nMbs٨��5j~�0o��{%�.��Jn�R�%��nb����m��lA�!� ��/�˿�[�u��k�2%Oa��������O�#��1Jn.�C�|�9���׍�b5bh�<��o?����ɟ�ɧ��a�g���g�ɻ��o�����{��~����|D�1��La�J��8����k�9�-�C��'ǧ��o]}��_��?��/g��q�L����w��o�xO����M���E/
U� �<u%9LF�4VC?;�ߦFY_z�s�� �a}⭵�������=
������ͯ������������6���;���(1�,B���2y�/�\�U��ʒ�`.�P� *2�H�h�H�Su3\q1�E�b��&�t�	�^�mh*�*���c��a�җ�����JJ�}
��zG��������{�>:ѳ#n���K�K�=zA�Q۪o������n j� 2 �(4@�?�����w��/��'��F���w[��B�Zt�K��e	d��PN�5�]>}<�������O��������T�nI�7��|�֭�k��ַ��w��<�����.|��q��^��G��T\e����s���"ܚ���g���O����������3Y1/�(�v�;W�����������m}����޽붻���3c�d�/:������hx.ҿ�v@�����g_�򗾌�n3�;���������O�����ʿ�ޏ?߽��|[߹���w=�f���b�E2�U�e��Rf��5/+`2G��ܾ:�Y�_E Rv ��L�Z�0<�)�w����?M�1e���o8s���-�` ��B�P03N������h�x�~��(z�cD��O#��,(*�&h�p�Tgm"C[Ѡ@֒��O�_G����Q fx�/|��_tP4��#����g�g���e����.�n6(@�9���9r��?�� T��{?{������o�6c��.�����=CXq ;���������9&^�+�0B ��
Ҏ����A���ߟ�N ��������������N���� � �|��_���1��n���ml������.�$�m�d?�l��o�o��\o��4�ѹ��~������?���W@G��w����?X���W~���̡V ���C	��S�������\�J��LUV���X{�Z�����T��jl��@�r�� /Q^����L�Bt@�zES�_�ju���0MޕE!ffX�̀pB�<)LP&��q�4��N8�MǓ���|/����]���I�\��.Y�������ï}�k�>�����H%������ɹ�U��6�z���=88�����?��ݽ=���^g����C2l!jcnܼ�?������~T�T΍�^w�E���@�ɯ:��zAߏB�N�ήo�}����;�����)�����
?���O�������Gǲ��f�*�@��
l=�������n�m��o���u����r1���~�������k�i��Q1/&��ٺz`��J�eꩂ��Zt��>S~�z:�,��S6��[��˪u�[�rN���(>a{�C<��>�(m�l�,4�ȶ�>!U�o��KI^-�ÿ6L�(vc�S��U�3"��|�$�>qʞ���[�)��&	H�{���������vJA�f��K���� �M:Gi
��?Ƴ-�3��O�b~0�=��lr)������o|�kkk`rZ�`�w��y��ڊO���_�¿�߂�''��L�(��O��cD���6H��|��o����t���������JT�"����~�� ��������<���'Y
�f����A���?�ϼ��[���ؖ�X�4� ��	�R�7~�7�f���?��?��#<1�pM|�)k�BkH��vՔ�;�~U�J�~�͕q���u=uW��O"�V���=ϟ氋^�kU%�Sw���G�RЇ��!K���4n�'���<,�+!��M���p��y��vϰ�1�Ł���.�6�e�x.˃�-�x:������]�z=��@�2�>�X�h����E��8���~���ӿ˱%2���L�9C{e^���Б�'���k��ַ�{û��v�J<�������v�xZ�8Z�:����������@�v���M�N[`vq?�*+{���{��უ��Ͼ�9`/�`�;��jƞb3�@�&^��ō�k7��<x �l�SX1��t5U��k�0w����l�o}�3�xݞ���5@��@��]��p
�8�����o|�{�I���K=NG]��ga�yQ��K���G��<F,�0Xeۛ/�	��`���^1@�E�֖�ܔ:����$%u����b��T��Ds��x�P����^�>,�Z0a:}]qB3�V�/;5]�e�?�D����Y����u���������U��3�r̸�F�<�'9�qxҤ�Mz|�qyQ�X)�_��\䕳��.�-T/a��6���,I��x�L�N��ApQD�h� �yj�l���(2J��`��/��£b�J��*֌+d�KǠs5Ld�␔��h�x�Xj͉ڢ�Ӷ����U�pg6?��9�J���X�u���x ��`���b�/ժ�_��5�J��;� h���"��ځ\����+¬ւR	ec_x��Ib
P�%g��w��S��ԯpYW�2H�[W`.�2��M��s�'�T[���;��6)c��R/'���ρ��2��Y�v�N�m��`>�	���n� ���Txa�^d]W�$3����`�aS.�9PXK�4�;q�aptǪA^��2��Y�s�.,X,��� ��"�<�f`
]����g�~���_�m�<TXZ���M��a_-�b�A�V,f*��S�"+�pKn����Ac�@�4Ϧ��}�h`���<��7�>E+��>Ix������nWge��Hbs�L����;��1�o�\�ba������5�j��A�_��F�
��U��Hwn��03�8�"st�bʷLs�M�S��˥�!/�N��7j�mB<�p���N-ݩ&����L�_�� yD<�ӁONN�;G����c�Y�i�g
�If	��;���&:K|�U�4�������x���A��rV�ƫQ5!0���oS�����Y
R[���t�V�)� �Z��y�t+vK��0,��)��l,��t������[7E�w�('z~L�Aڦ��������p�Y��)�R�$F��yE}�p{U͉Z�a�� �c��~1�M90r̃Xo��$��'[f�n���z~������|�/�a{E�gI�7Qg�&��r�nf��8��η֮&��|,�s]p&.�����ٔ�!����H珞M�,�]���bч$+�KZ���	����)��<O����ë7�+-;@V�K�J�m�*�����>u�D�	�Ц���YVb�K�t�/�^x�����?{��΂5�iF}�L���@G�{Fd��������y����@�.e����j6V�M~%
��3o'�C����������$�q&/�Ȼ�ꮾ� q��5��(�]ΘI�����m��vVfk2[I#I��k$��}wWw�UyG�������� h�5
YY��/��~}~��w_�>�yW�(QV�ДN|�/3Ե:q��t<pA��9x�rEY=U���TY����ԤH�����A?�J�k<�Y%��+�]��}�t��Vv�����Iu�u %���\�M=o��{ 3_=������PչH���(pAB�(`pn`%O�*���]5�u��DY	��q��E��h���y!���-"�Ri���"��)�Y��+q�
mk�$S���{��Z�-�㹖+Lز��Ȁ�2*���M?�~$*󢚝����f���>{���������)C:2]���&����}������-i�Υ7^-�Wҷ�����~�_�����Q��g�0����|�s`�hE����7���^`Y�r-e�i�P�!!��ܻw�7ͦ�r)�c��%��@����٧�~s��b��+�
�9�8a��:�ܽ{���C��RsF�����x��կ~E�L��|��NZ�@�ˊo�	�7A��mv���c|N��D��x֢��][��
%�뮤9�9��<�������,�*���q���������Š�9�e���jQ*�>Oa�������NIȀF��P��$���4!$V�XL���1�@��|���]�q��?�q�����l8n�X�B�b���'�w�=*���b���A��!'�J�F޸��\�$�t.n��;������?��_�%�.���[EgPk�O>�.�������>�]�3�^i��r
*�j�WB��ы�������[W���8y���W�~�?�����H1 nAw��_�������������A�Yz֌̛c+O�w�cX�d�.���[����ѯ������J��<	&�ౝ�8����}v���'gg���O�|ZL���\J�mlU��w����ɃgO�.�De"�,6����I'hs�:E4�'������*#��'�ǴTL=���;k�/�t\�:{y˚y�������k�)}#�s�w����E>�����ϭ\`&
���Zb��i!a�FJPH�'���@�<���GB�?��oa(�X�
�'������{R��{��Ǵ�"��?.� (���x�\�t�ʕ+�hW��'� �����UH%��m� B:�o���kA|zu�4b�>.yF�G>e�n��ߎ�x���ƃ��o��ι��w�g8� 7�OO�������?}��EƱ:1Y������3����.\�@[���?��?"���'G��Eė��>�裿�����MW=�Ȅu�m�+k��E�Z�9I�^��9<�����1;��GuM�l� b/U)9K��t���;"m\u��8+أ"���Z]ǯ1�^�he���v��iU��0C��{W֍ӕ[�Z6�[<����<�w��{ŏn�����B���U��a2��V޷g����ӏ?����i\f�X�;����r֠�!y�m���ݱ׮��G�8%[�y�ۘΎ�����{����ѕ�[��j8�x��~��fStXMx
�մTS��T�(b9E;�V��Ou^��m}k�����~3�'�|�g�g���T����'�|��_�����bt Үk�l�u��e�*�0��.q/�}�&�?�ǝ �磋�7�G�?{r����������6�`h/������������/$'��ȉ�^�:��UNC%��Wd��0:N��՞�������������������~���N��<2toC�~�����r��Yk�yҜ���YG�y6ѹ��]9|�&|�Jm� �E�
��t\M/5�=�dmK5���HM�طNa�1>O1~��3�Vk>ɉ�8��ʢ���6�����Q��;�g��5cq��c�j�&RUQ��(a�x%#�Y~~�%�3�
h�F#R!�hZ��A�nb-� �l38u���@+���6��*f�w9�4ˠ	�*�?�s��B���R��d��)S� # �L����b��>zqLڴ�[��t揞=���W`��B?�oe�vȓ�w1n�,�g�<��÷�zk⾠��{z��l��e�v��$�z���#� &��\[kk<;S���c//2-;DP��˗/�Cڟ��O���~�&�3���OO��G1����5�;o_��d_�7���<e��ս|�������~w�_��_�y�[�o�N-C��t6�#O���Ђ�lΈ�;V$A`\��V�Z�ڹ�F�B��ɓQx��Zm�V](U9���4���a�s	�4�'�.�b���	�D��B���z^�e�r]�-���o��Y��:��-��3/���|M����I�OSǬ�.m�ʋ\���rt����+=^J���G��vW�T���p>�|������0,�l���[x@=�֚b�c��V�`TD�b�;����~ߝ9��lX���DgFk�i���}�ʲ��|�����:~���FH6/�0C��kr�B����*�5�h�ך��֣�{{���^:<b��~6���#�<��م�ZY�/bB�0�LHV��^F�Ɍ�KB|V�Y1qA�����J;l����>|�1 ��q9$���e�\ml��띕��cM��Q�Ǔ0x�m��g�%�WQ=e=*F��.]
������&g�?���=�zE�$f��S��N��s�}{�(M���N�S<��/��C3!��@��RS�O�ʘ�*)�_=��7�x��!'>(T��©(��9W���>a�P��V�j1���iQ�E	&�a:~6:>LG'j�V�D��*a��j�09Z	�%�Oå[���W��+���2�]��I��i���ch��U
�A._����L��բ� 7N�rN�SR'�=����^���D	�R"�ٶ$�IVE!GN��hF��W�f2f�֒��B;��e���>O�� \u>=��>�3��9v���ׯ70�ނ��x�L�Ȕ�l�E�z�8�U8j���ú�Jc�,���S����45s>���I��6&	��gz[�N��4�q��Ю��"����E�ف�kk���w����9��q�޶V�Q�inoo{����ʒ�Q�AO%��q�|$K��S.ԟ|��yAW�n�wg����뜲��昧P��Q�!G��aϝ:���M:Ϫ�A�/�%&(��W�c���%�t+����)�M�B'����Û}�b��6� �E(�n�T����*.5�I��2����%}������|��������D�z�V��n�k�h��%DC;���PH;��[�B��^�]�g���{��OHRb��̥�H��;Q�`�����""�!��[:��M��i]T�a�������>���?���5�C���\��V^��$UwڏIs&|Ұ�shֆń��pf������xֽ�A�OG�x�V������,k�j�ĆN#�C��Pe1R0Q�}ͅ����X(�^�y�䥒:*��lL�m�w㢺��I\:�~�6������n!�54�n�V'�V�Q���r�яV¿"D
 �N�4�b�N�v1>9?�C���5g=��M�zV��=�7�9��&"RN�=�����ݣ��%{��}�sz��[*�HϖY
���U�t��s�����b�8B\Bŀ��'�IZW�\iE�8�"�����f�ů���SB�4wx[����ϟ�}��������/��Z"c��FW!����Aݜׅ�+'�d�j�y�ЫWX�F�?�Bp�y,n+�+�[�s� ���Q�� V VS2�PF�,z��*�@3}���U9���  �d�󀎘�����rE��E�؄��$�.O�N��u��zoccCu�p&�g�BC`��SѼ.ꥌ���.�R8�k6��mh}�
"�لmќHʹ`��"t�gcLS��H���veDN�E�wΟ��gO�'Y�;Cܗ��k��@�,E�f�Ek��a!((@"�d��h��Ug6<���ٹ�m���E`ǲ���4|v%{�u�l�3�bt!ח�U��T��܁U�v�I/&�=z6N��9�΅+ݕ�(��X�8ö�>�F��3������ g���ylƧ�b��R�Y������MlY�9:B�a6�BYxE����+�lRr8Ey*&WI�~SD\� ��)��&8-u�(�ɜ� �c��5��v�t-�g�K͵���e.y:m�vu;D�3��bڍ6ISpy���V��)]�v�(?hc���4v��s�	;nN!
�q��c�f�09�.��w�hm�$)��Q>��إ�t�$�k��
�3���<f�z��*��\��;`/9�ro6�d��%�$�PepZμ�{XCY�����Щ�x��n���}n���P@��U�� ��6F���:�n�F`�)���r��':�;�ˆ��=�U�a�����<�z���1:���N� &VB?�>���_�{�P>	�y�}0�&p\ȏA|�7�ޫ��_.�:Fz鸛�<��e�)[��cK	�� Դ>�][����)�5��d��95�a	�'!i�e�0��7{��#J�,8t��yz�e��6dQ-#q�@	�o�y���� !ԘCJ��	O�.3���~�:a*ּ�8h!�[�Y��"�Z}���խz��֎�(���
��ɘTc�4��4(�R��}k��J�!d�h�B;�17����$߄�%��
�GW�(q����e�H�Oh?���"C��b���R
�o(�]13���阩��"�D�@�lz����Q�E+ox
�L�S�|FZ��aA�8���|)�Y(N��$�A�'w�4��>p�w�Y��i��S�l2:��)S�D�=�u�C�'?������t�g�T����,?����^h�ϲ!:׉��������4+Kʱ���@�v��҇�گr�Iʈ./�4,߯�٣�?ݻ�ۤ�ݽ@g�j�h��\K �-+��Gzt��Y���)��}}V�E�$W��4-���-&��쯠�Ҧ$����'�L�]�bdL��(K�5�*���2�!�z$n����A�H���4T�+��q��`'���寭oa#��HP��Yaɉ����W�.��[m��9Q����̖�0s��h�g�v:)�eO0.<��"��ϕ�(�ὡk�e�Q�K�i��(�NI�O�[kg�bdV�\	m�K�}��@) �E�X�o_tS�gnCU>>�.����V�	W�`��禶ѡ�X3��t��T�gL�
J��z*��� ~V��F�wVo�}�_�,�9{,P_[��L2��pF����O??}HZo�<-�ű��m3�����h�(�˓�b�DsW�HР ,���2u*^:_�[l�W�cXC�&�K��	o��xh?�L�V�d�����E�E2���$��)�u�:%I͛��S�/./v�22�S��О�裏HO��Vȫ˺ɠ�Bt#l3m�J���6<���8\S�)!���Q#5����!;���P��L�k�z��X��:�F�5�$��B�FFF�t
�w6��Ld��q#\�lԊ���Y�3`G �dTSO@_�oa��tIg"��2L�����U�Z�@��V󉒾��R�Ok���*�{��8,߁́�z����s�Ǚ�h�W�y��|/|��ж �?�wv����lt��H�0Ũ�INQO4;������+L`͕�$%��5з�L$���yt%qR��⳯�({�m�m����Y�͙R�$�?�*};#�<q �!4�������M�f�([tx��I��#�$�>�	����L���/p�wA�\��.*�l�8TC�s3j�Z�n|����t���Fvq�&�P5��Py���A���T)����ȇ@�)BD�r�O�0�d	�`g�i4�i�<M�vS��X��5b��$��~�C�9{�Y�5Izl��1Kw$��)n���\�H����LաG�ŀ�el}^���}�=(�}t�f�}�l7�#��=�uj��/<�2�2,���b�7�����З#L���\#�X�]E��T�*�"G\z�P�Y���mfM�1V�6&?ԉ��-{�g���a4�6��X�?G�G�s}�Od�"��1�Rr��t�1��O�,\Ħ殷�y��X��s��v��/�����y�5�zJ���r)she��R̸N��[��6͆k��=ͼ�\�z>H��� <Z�h���fid�.�.1<A�q���$��;����$&��H�]D�'�]G� {�#���>�ئ+.Jɇ��x�f�Yh�)$]G_86�ܢ1��c\�8E�;����p6l��\��{kkk�Ɛt���D6�0i��h!�r&�8��3�*f<U�� 3��"ߐ'�A���x6X�e�<��-�%�v�%�4)Z+��g��^�0/c��%u�����f�YhL�#�;Vb�(��)W�Ly�eb��yD��'^j��Z�괉Z���Z�:?/%�u��ܾf�X���7-E}"c8������3֪��3��Xy^��<���U�R\�>�?B�%��1�\z)0�R��YEe�1��U��0{ܚ9���GN3(���A��.-�����c	>4�5%3���U��8�T�M�A�d�e�,gP��94_4%%Eb��.�s+�H��*mcݲyi�f����%+Lx�3XdMv8�Zv��C2)���툄������Mxi��<�����UXRW��1��5��kcP�ɋ/��k)u��h�W69�N��RA��W�`�Ι�İ���+�qE���}l�e�h����u��}��*��ùz�:B�®P�����p+�96{QA6��6�-�l�
�o���?�*��P��r99G��ĕ8���t	�Fw�A��Y�6����X�	�@�c�a���R����w��p���|W�p��:T]T�{�9o�Ԍ���t���t�K�u��~vC@��"f(��������[l�j��Y\F�w��H�4}r3�Ǽ6t��lC�tU�\uȓ�C�I?�(�+�Ǵtwk��_��)6[�oDt&.\�}����O��\������8� _֎
�:�lS0;.az����������!��_�Zkk;A�v�\yև�y�� �x�%��ԫ�����x=�<$������]�<�:sn��}��2l��V�>fb���<!�b��wf�Җ�S���=>�sE>�m�f���F��X�5'�kT��^�yhh�V�@�^[x�En�er�$�E�/�Qa0�#�V���BO;aYXXP�ۉ&�f��Eh;�w	)baZ,�x���'��M:�6�4kwe��˭V+h��3'�e�&�����k�ۈ�ƨz=�M��]��,/���l�pn&9R��)V���%#��a����%�N8��������F��-�3:���d���l֘h'˝	���]�>���o�g@e�O2Y� �9�
[ș�S��U��s���G�$��C�h�T�H�W��cg��N+,�GI���)T��	8;�rv-li�:��[��$܆�X?��'ӂk���-P:��a���sY(yw�21|]��^�F�i�tu~-� �0�3a/qQBk�ùp3�U.�N
�X;�KxW�ܼ\����VE>�z����\�tQ�̑��*֐;h�y�I2�fN�$��.A�#�5��\��9�6z�{�{,�-�?��>��8�2����w�zZy���C���0Ox���z�r�A9=!h톴���yx��1��0��g%�*�&A�6�vL�A��2a�OO�<9>=�w�2������e��q)֋�s�I	������T*4��z��	8"���t���)p�gx�^C��őN���&�ýx~�)��d�ڶ�Z�� �:�2]q�\A���H����%���ٙd��]�7]����K�lW��zl�0�W��rrEs�z�!Ɉw"=�;ai}Kr9�v`�Y�j����բ���.���lǵ�u��?�j����V19x���' �@���d�1�ă^D1-�q�J#��/<#�pn�́m��JHq�qF��i�h��4����`�Ԟ)��Vn���__|ao��~�>%��Y�����q��a����I;G�m�A8�<ѕ�wւ����SQ����&���\f� ���1d=s�Y~�h��m$��w����l�`j����Y����ӕ�
Á�J�7U�vC����S���1�:@�oq2�8&G����w��V%���<��/�_A�ζ�?���M�N}����ub�i���'�`��+콰	6�N�h=<��n帖k�hj%��
��(����0�w�b=�]�W��P��E^�J(^��:�y��x>#�����\k��&�b��8��Y�s�P��+QmRV؁�I��r�T󨡚O�񬗚�j�,���Gz���f^n�lbo�S��4�\�o\rY/�~�\�9U�ZS֚�ѽQ���E���pw
��TǺ�WlYk�������Z�q��[o��v��78��._�Lg謷H&����������7�W�^�w�t�/��kn��u���r9�,XN�;B.pX����������N�9<��ƍo\�E�NXX$�]��ɳ��S�A,��)b����s�yHaJu�Z|��.��8�Ԅ ��ߚ���:B��Y���G?��	�0�:/���	�z��P�%�o�93cI�/ΒDN�Rc��#��*L�t�|�<d�20V�B(���R��B>E�c{-89�e���W�-��{��&��Ϫ�V�fg�Bg;��_�7
�E
�W�x���h4G!d�����ti��@lD�u�r�v�������^`�g3R�<9��Y��JS(�ʲ@�/�;�(lG�u�1N�<yvpH�2���ۍ�x���'�';A��M���^�Oig�|ZR� �ޞ��Y�����`���v�u~��NU�j�r��&L�%j�Y�Q�:�^Tӭ������z��g����
&֌�^o=������=��OF�r�C{`��ĳG�`�"�}G���ǹS�^h��B�QB�q�ʷl���ȿÄ���d�0Uq�����.�V��5T2E�j�T�5��)��Fe��G���f���5TL��L:�M�����"�zP�ӹ`ϫg�%�p���G��ݙ2��9�j��S�ne����� jOU���w`p��EZk���~���%�u����a�~E��2f]��|�@�9���u������幗.]b�.cq�k������ ���u���W���~�E�<9W�2l�|fj�C���=秅$�x؅a�)�l�f:f�S�Ugi&�I�����"r�tHC�F��~�	�]��9p���ÇH�J�P�08��Qm�0Lrf�@QBwņ���<Z���q��4b�ړ[\�)y�{.��������4@;.�O������q퀞��E-�b�Լ�~���e��`���9���������J��X$ҭ9�!��4�~���]��G�U������t���|���qR�Qm�B�8k(2��5�I0jS�h�Y�I�Й�q�[�v�_Q�KD��j���z���� L�kZ�l�����"-��βx�����:�K���p�e�v�N�^���=x�|Ԅc�Pw��欿3�s0�lۃ��+�Q��"�=j8�`Xo�3c�����V�U^I��ļ���^�g��||H�}�5�ӭ4IE�h
\э��m��$ǳ��ˬ ,B�f�ݼ��Q{k\��|c�*I�h<��;��M�:!����9�6��tE��/ ��f�*����'x��4/�ܝأ��t����9; I�;�NZ&`>�;���,�e�� Z���S:s�e���`	:v3�h�B�+A��������,���Xh.a����~K~ʪ�-Q���ܜ%�6H��Y�1�R�O�%u!�J��o�y����p9!¡\�,��)�{؜)��}�G�W���@K�w�AK��7��[�hD���9a��c����;�c���80bË:>>&-u��ţ��^�G��'}��Ǐ�+��l�s� #DZ�E�IE>����V������*����x��������?���X��/^�G~is��Γ��n_][[����&�V|t�X
�7��FL�s�/��=a����Or�U1���~ Ѥ39=<���\�$oHpv]�@�� r���^�#������?����5[[[/���GON��UO�c��s���e����˲�HW-�6K=�R�Wa���1�<�d+��i-eL����+|��\zX/�7��T�=V+�-3�T�8陗55�;@��d	�~��	�u!�U�yN>���X���pᴙXU��(�rxl/&J*[8#��BK��j;%���0(�IN��7�Vo�$=E�3����^�z�R{վ��{4��]�Z�ӏ?Ѿ]��Y)��+��ݙ�sGe>�U�)�>��������t�Q�^���EњlA��4��3�bϋ�����]�wGv:C�x0؏�r���	��Q2#�x��u�������U���wm�Q�&������+o_Q���"�����Ƴdk�v�V�R���f�[�v���}0BG���G�5u�%��S����o�y�֭0��k��|�wּ�e�╭k���?��ڴu��d�!���76vP¬�LN��~ ��s:�yF�%U�U�tU� �%t!�U�
��3�Ru3%��<�F� ��6u�Eq���g���V�|���s�e�u��~U��y�p�?n�{���.����5#!�_��g2�8����\9WH�Q�j�j+������C��\���!�s�m+9��K�|0���'�;�Hs������Y�'��
�u���p];��(��0�f� �)+���Qa��ͩ�s8�u��d��.��0"�HO|=��u��
��x�'.:�h�ҧ��B{mccc����g�g���X�ڤs���FQXQ�X9&�>s�R�,=�7z��ʢ��������{��ٝ;w�r��?C�U�Da��ZX�W,M�Y`Ʌ��ْ�#�����,>t,�+�.s�\��$�rQ���zi����e����u�*s�sh3�)P�!�.��@�1�W�vg���z�/�
��>�'�Ѕq�YA>��=�{����c7�cSҿ.�<�/ST@7��U���@��K���90ie�QZ������Nc5��o�^"�tw�ģ�"�v��z�i�+��i�t�޾�V�d�][�$�
�)[��X�s���F�<���M��麟�n�b'���je��k}tt� �� 0i�%��u���ߟ��@u�)�7�/^m��������֭h-q��)S�i��Nq<n�f�w�ݮR��~��sU��$?:�b��\#ϧ{�?��"��[Q��f�M&�q���<�p<gg��z(�o�[�]'i�:a��� ��װ�O����ы�;�������������P�&�����+�[�:�]�L��N{s��D�h��%�o����ѼZ+�zYR)��6ZT��xZ����E�C�c�.ĩ%�u��g$��0;�3�xX<�I����?ej��P�0?7�HZ��":�"?�KLr��j�������ܤ7$��q���n�𚎨��7.�����%�'�uI2e������o�׿CH�jz2,��jRNONN�T���N�a�{�%!�D�>3�Ŋ�	�)�0���\;������ܯKn ��]��e�?E<�#'AQ�M'��W�WO�����Z�������u�i�*�@��q����ۏ��\��.��w���v�����o����O?� ��!ctpbF����ҖEz�ڍ�t��'����H��|��?ǢY�{�G2���߻w��4�\i����/��b��k�L�Y������;��U��o爻'W�w�:�>�e�.��?@@5�H&R�e�,���)�_ܼ���E�Zr;������{�c�����@���^�9�gft��NV���m�������U;p{׮]k4|�Ɵ��ݏ�ě%M��F���ڞ�ʍ.�Wv�m)J�ܮlD�K�����YZ�3W�'k������ó�����6�8+_�t��y��wɧ�|����pg�
g�����+�"������%�85`=rRf���Z�u����J���wrX���!#�����@ǃw��ݺ���&�io���sK��v��Ν��.aTl^Q�F�O^���r��Ӫ��T�\���x��4ol^6�,�!Ӥ�J�����Ƌ���]�	a�"$N�)-�y{c���P}��'�tH|�]�N�n��9�;�Q໎r/l5�t�Dʍφ}�>�����7=�z��ەq&U��:���a�Wgn�V[g��*��07:���h���s??�B!0J/ ���Hj�>k)�nF��J���Ǻ�
��t&՘�]q�-�9�k%�hα�Y$�l���N�]�/�_Y���Д
�fRɴ�W�{����y��v�w��J���+&.�w��V��s��v��2�r��E�j�?47��b�y��D
f�K@oqZ��/JƔ�v��?x�`6��
>ŌK$�r���M�|�fN�+�VJ���P�$� �,�~�\��>��s1��!a�J��(��y�
7V��V�h�t�� j������γǏߺz�4��n���y����&�u�b	���[�ė��΅�f���y�=���~w�ƍ���tt��'R������#J,�C�Y��޲��7�x�B\�B}�4(�������!�R)���*&�� T�^���Uͩ�˒��v�ka{������\'��<�/�Q���$�k|��y~uY|_���[¾-M��&��e�.l+Vt�������kH�Κp�T���g�������n�u6���N�Z{n�y��b��D��aiѿfn���J�62��DÆ�}$���Q��P���Y�[��I���� o������������@ϠE�]�0��2�ꬎ������f�,Xx�������hְy�L�8���ҭ��q�U����J�����������$9s����dwtJ�vprD'{��g�<�:�*kl�4�W��n��a��۳�t:n^�i���6:�p4L㬅���A�Bk5(�  )�In��4}$��L6.���{�����9O�|������~�뭭�|<�ȁ�3��dB@���v����b�\���4MtU�Ӹ�����<��y��&Ǫ�I�2�F��05'Zi�]���R�L&5I��x{�Ͱer��|i�H%��Z��˫�X�_��	��0̑�
R�,�a@`\xQ����p�y��\W�ׅ9�/�d� Rc�L��I-ԓ*m�� U�E
����_>B�"GK�3"4�S���˾H]6]�EL�Y�"Y�yt�|������d���B����1a6w���F��E����6{�s���>(��D�����>���.'/�q�)UT��7�A���0�������$��>}J�	����)-��/?B�� �{��U5����U�[��)�dVI�I2���'�i�666D��:�&����ޢu �@Zp{{�����z��f�l�5$!O�$T-�$���8l��0��|s�E��f*�-u9z&^���/<��|˜�m)�M�R,}LQ����s�|�5�Z����Wg�7Ś��,��eA�^��hǐ�P��C��%��ȫ�r���nXT�`:>������ۦ#L0C�S�����hu�3����=/
��k���a�\;3ځ�C��,��]������)/�ΦJI�����o!�݃����������q�ѱ� <�r�B*2>$�mX��Ml�e�;B#���*����=&���y����ѧ/��6D{�H�{)G���U:���o���PA�f��s�;�d����OH��av���^���..nn��b�h�aM_��Y������u�IZ4��L�۹�GE�&���2!������)Y$r��^D�(���nؽ��O��ˋ߼N&�����n>�~ա3��*p�_c�C���� s��G�wc�g�lҲ��֨*��6�^t�&�h����&�D��픐B��o<*Ѹ
,?2!H:q���a�4�UF)Q�g�3��Y�����/5�{�pe��U�?s��'q�+�d^n\z�*�^ ~��U64�Lf�hec��j���L�0��w�}�~��H'�͛��Y%#h���Xp^�b����c���LY�sf
%��c&��np͉
�W�'¬5�tO:������5W-�����{�<A�C]6�q��3�|��U���{��7����W<�<��ZFy�D{�M��^$����֕+W���h�3	$���L�e�u���Rw�\��6����Og���/޻/,p+}OHhQ���9��������v��|�2ir�~���O��B7!����;;~�۝�,���٬�8���o��`qf����a�z��n�[r=�ˮ�ȷ�*k��$��|���dF�<I��TK�2��Y�@_�K@coq��\��z%鯳t���؏ �x�1��E].6Sc��k��J�����$Mǁ}�J���c;�~<�}�{��㏐m鹶z-�4y6���O�(�s����}��������0-���^�7+-���̞�r2�M�'dfn� ���l@�C'M��o��V;��Ĳ	YO�jݴ��͕"-�f�k6��-R��>v�,B�ۑw����JW�#�e�t��m���g)ڊl�L.�F�!�d����u�N�p+�NC��]��zwx����K~��ŋ�j�m��ƛ$jU�ӄ�>&��l�y��N��O�*]68�&{��Qb%�v���'��89�������t�k����n�r����LV������w���u�l���[�q�?x���s���FT&3����A����[����_|���yJg�����ȭ�7��VO,��;�
��^i��J��֪����>�Z�%1%`�XB������oڶQ�����;$;��c��.jߌ��fu/�ei`�KuS�O:C�X��1���Zu�꼶�=�|� Zl��f�C;��w���&Ɵ?dH��g���D������Nz�h����.ifQ�]�5�X��K�l�\L]R^��Z�yF��v?�{�-���h�ݵ��~{ԩ~��_i���,|y�z���ÏE`aщ��i��/�@�pD���7ަ���yr: ]�d���)���o��%K�`<<�;�ʳ�cP�7��`0�XEԌ�I��$�$��d�h=�����ރJk�?|��'�	����=�Vk����q��~��q�ݤH���v���w>����������������;�tbvH�.���۞���B-�pG���A�v�y��S�
��ʒJM�a��W|�ل���K��8%����s�ϲ�u����Ae�1a_�kG~X�d4.��n72�<�f����d|xzvV�bA�Ofqձ����"�u�:��k*�N�A@R"X	�@�-�j\��<`�g2rٕ�	LEPi�(��q!�曃񐾽O����X!W��b�e�HV����?�ꢉKNE:maE�1.��Y���?��0��F�"m�c�QpvJg)k�����2	e�?��~��E��U:U�����Йg'3���1z��3���x�%���w/�E�yz���z�x5.����*���t0�l�4��č|�M�T͙.F.93��v���s�7������;�F���v�;?ٺ�y����7�FQ��b�V�St�u{�hq
S���!��.R�̜���ӅO��kPp����4)��,S�"x�x(T�mT�.Z�C��A���=�dJ�BcV#.�E^�:;�S��w
A*Bxф����Yv�>�K��:_��.:Cp*m�A��E����.����� ��mӋ�F��矋��yP���D�Z�4-v�^Ҳ�c�몚��#����l�޹}��G�}EJ��x���7�u�T���v׵�x�fN�'�LϧTʚ��=z��F����,i�}eueU���x�`���Rh�~���:ү�z?��3:έ[��Y"!��y=�	���w8拓%X[��WU�kðd9*̑�,F��	x/�n��-�N�1i�$On޼����LF`<���~�ǵ�H5_�Zz,�'���DW�H�%%�3"H\&F�.�LP�"9`Y�8Ad���t�� 4��[�1���Ni�ׯ(�?pS�� '*��?$�lM:�C�����ҋ�s�M��.�lЉ��/���zB�d8������x��@��W#�K6���?�v�to��A+G���c��?En��`�PN�ĵ��V)��vi|�n��$h����3t��N��q70�|��5 Ę��.W���JY� �x��Cn�W��~5��uZ	<$!��&���[N������K����o^�~��-x�Uj��$���n�E�����Z�+�����_���KX*Tj�sw.���\7L�!�N��*K*�+��D��v�:�3��2m�E���l�	������3���u���P�;�����~��0�b�r`RM�������4۹��+*u���\�6���aI7%3%�OP<bc�)*�������2�����1�z��ice�E�3
Ysd,\�,}=���ji֖Y��|��/�9�R�Hs)��5�i�92p��v�M�g�8�h�!��v^��.y���Vx��B���Dc�_�W�c(��;R��'�����:����*�w�hL��vW?O�0Ҙh�I���:C���~^��_��?���<��C��C��r�O�.�^{�5ң�ِΡ����M����DB(��,�㒆6�18v�L-]t2K-7������;�cH�Ykr�y��*+����O'����Sw��#�T�@-ges؇��8!*OsH��D0�<)7_V�_�n_�P�8��<�.p�y]j����1֧�TD�i��u���U4r`{N)����a���Wb./?P�˭n�t�/ChX5��-r�M�Ɲ�^O�_�^�8�3<=E}��Z9�cx�{�iefn�lPv�n�i;݉�K��3��b+0]�R�$V��*�l6SE6�U�@[F�M������ɞ=�>z��prFG���7]��V����wWߍ�5ky�+u���=���F�H�o�0���0�dLH���9�AG؅�$�^�͵��`ҹ�t�4NQGy���/�@N^���:ݪ��<ʬ���y��~�Z�6=N9(ī&	�H���J�3&�7wm�QެLJc'��շ�vR��܎��#�@�r�M���gy਩J�1���4ia��c��Tj�{�,�U�1|�.'�&�ы,D:'��
!����82K��:��m0A�[�:y_o��}-@���pdJ��UD�g�끓��4�WS��K�_��.�.a��g��_�a�L~^�콌��-�o��pVȯ��.tXT���HDI��G�tG��a��
_H���Bo�y�� d�t_(H���X�ܪ���A��t��z�DƼ���B�X\Q撕�dd�|p�ά�Kn�-�g!�_~E��(��ZP9�]�^M5Cg�0�U���숶�Z�H7n��S��mG�'��(�Ԣ�Z��U�ݟ��Ϯ�~��1��h��B�s��ݠì֤��W7�{�
W�'͜�����������bg�W3�s):_@mq���p�}5��%�1,W�c���.�$�(̷g�h0�3��g����wn0@J�4%ixu��a%3��H�5���%�+Zͪҳ
�H|n�"+�>���eQf���(
{��B��]��ݢ��5������9<��0S&o���p���l�9��5+$�\�L�)� }V6�e>*1A�U�͕|���ǻ�?�tW:M�`	��/�@,�gt�Y6h sQH6�b� �n�����:��3���R�\e�x ���n�׮잷?=����p�?ene �=���-w������S��������ի��h�(l@�(h0�7tǬ���
L�RT��Q\���:���rͅ]�:3��U��^�W�W��0m>{d��6V�&���A����;Rˊ�+MH�l�N�t�Ty�b���#8g���� �%w�{2ߞ�Wr�7��vl� �����ʸ
d�uL��k䖍!`���Q�fj�m�<Q�ޕ�H�|F�t ���v��d�n�-�<e�\�W�;�n��Is<�<$Ը���`0໘�Y%:���'�����@�s���詩ǪC"]f��%��f�D�Y��H�G����١�;�:�A�%u��sTȤH�W�Ʉ���ţj��]�Fl�Ε����Z�آX�7�=���+���30���!�X����C�]�x���۷o�J����e��L�Z��Zg�/#��O	��Ҝ<.R��p�_����g^���ˑ��`6.���0�@�hk�h2c`.9v��!�Ԥ����,���Z���*u������Lם;�gh�}�8>)i�R�Ռ�|���-(����ה��t
F%�1=��-Z���T �<T"��4->ܽ�Ϻ�T��/�l�����"�=��&���S4\ص^��83�g2='s	�U�7L�]�<�䧻\�D�=T}�B�O�PH���EU�)�U��"[�
��n�7/�����H��*`67��:.�A�d����a?63��^��F����y��:�{��o����l�7@�������O��ɷ|;m�v����f�D%���A�`�QQQ<j3#x�1 r��wp��Y�R��0/y�K��h`�%W�(p�!�Fb�a�O3s6��/8����؛�����Oy:��Q�Lt�ې����s�?6��t�ӳJC�1*��P���"������k\W
x旔U7��S�	�Gf-t��T�~Tq�t�k5K��s�$�(��N/\��[�����EZ �&=P��	�=�<��`h|(V͡Q[� ���g����g>�O4F�e���ja.օXUL���+�3!
[:�aL<��,nM=�7J��J�k����R	�C���kY7/)��o�7z&֜AWj8A�6��;5������ZB���|H��ڶ�&!�f	���<���`�t�E�����ǯ�|�p�d�`%k0���Ֆ�Dh|��&����>���42�oz.�]��ea.�k�o+3�;������u�����ͻ��%ʜ7�|Ez�̵��T�(Gf΂�S��,"	5���ϸ\|�k���bZ0
:sTb�Ui��y:����U�M�.Sz���n1��y�3��u�5e
i:�Q��a�R�C�P˴���g�I��5k
L3Z��RLxq&.F���bx J�
�
ɉnyV�?�f���q.�'p3�j���7����K��om]9��4�E��b�BV�f��/["*5��4�濠�B/'�*0��2h	3{ٹ��))��!{��	��\S��ǔvi褞5��QA]è���c�23?1�
��]8��R�1��x x�I&:�K&uD�B�����l�5�,�eGYl,��0���t\�v�]b�P47�8":�Z y*�'<���hKӺ���:���Jg>�:�
<��u�v3���f�*l^��XsYK�'�Jd�������6�.A�(l��)Y�|�U1���"s3(�y�?{`�rlx�;k)��?��ȉD4ϛDM]@�޺>�ʠd�H�ߣ��`������]*N;�c8����*�4>�_��G��:[�';.~]z�!sVX�i�$BC��]B��s�y-��:2fr����������x�>`m�J2�7��|h�
�������i9lQ��?�:8(���޹�4�Y%B�W6�ᴔ��bA�'N*� >�7W�f^C1X^��T�6.�È(
���%�j�^,򲎰�mf�A;��uEk�5�5�{!Ý�N{�a[)mK-�aD�$T�u \1� mR:�Qi"���*�|�`���*�Pz�� �m&^�=�ح;&e�0��`�xG�ܯ�� %`��a룙zq�@x�Ψ+ԋR�_F��׿<?�S��xl�g�1%����b*��\{s�֭��ݴ�����!DB�T���[͹Z��O��us��-��呱�9��a�)ɪ7`���@ibT2�Djܕf�
[N�иm���o��]���!�I7=T5�<5xjP;�k����"3s��C��."��'�_��'j_�eXs���v�������Kh���JX�a7"Fϙ'5���N�E(&Rf� ��H��r�,��5�d9*Lj�P8X�y]��+
��P/q�*#���+|��5� U5*�Q�O��+6}\]F,�R�F��9��H/�a zޫ�t��ܿ��[��0�$܈�!~Z���e�gy2N��H���Yv8WW#�gE��WY��ː1�vニb6Ŕr�o8 ��<q��\<����
5cb�`��œ����B���+o��P��'��!-JJ��'SCmYm�,�(J�KPmyY6�?�A,7�~����!7<1Z���wU�ԢX�Ew����� �='\Ǽ��c�pq���x����L�P�����NF<�0	�b�+��q�_�X��WV�˸AsB������-M�j��U���/�ķ\U�)��H��,:O��$Ϣ�nqx�����-ݜ�7t�8���]O�VV=;M��S:���R���T��eFٔ�4��!0 �+B���*TI��`*�9����d���'j:%�iq�j�hߢڅ�W���rk=Қ���Aف�5n�Z�.sK; ��n�y�?=�xo{���8�t��`t֘&Vɰ��<����O�GN�t��`(	1�\y��`
%���Y�挶�8�x��$M�Б�U	�����Y����__�6���ѕ���|��$�3{3����8O���^G��܌�"3��<���[�	ZpE\q��x*]��t��GL
C
 �az��O��18�r������GZ���d.��}�p�o��y������˹A!�]Bfi�AB��5���������y�P��Ns�r|�#�_r�D��G5
�Y*�@��-}���p�9$��+�t�5����m'j�U��OK3]�Q�B���&�f��k�8�4�[R*!��y�������������B`^g�Mh}��A���{�_RW��1����G�ѝ;w���y�#ڣy���J m��8��������J����9�0ٻ���<FD<G8�������7o�|��:y��޽{Wq2x�T�������m"�#�y��A,o�'Bkb�kw����]�����TT+G&�X�)m�}�"t�>pQ�w��=���h�	,[�FKT���x� ��[//�D����l_V��J��r�ԗB.�_��7�yP9w�n��$
�!�Xi)2DG��K��w*��A7�T�/,���7��&!y���&��g֊��Ȅ����al	ւGk�/u*�$X��p��Q�IfϮl+V_�H��[V:e�M/8��4K7�yZ������� Go�+C�O�`��<A��䓁��'ۇ�Y8�'+��8�3����\�z�����z�x��՝�W�N���/t��w��o\�5��m8ň�ۯ�4V�& [��d:;-f����UEn�0u�'��v��۩޳y�5�"��Ov��T<�t�[WW8����c�0jVM�O��*.ɩBm�	��[��e6r�G�8jE[bB������-S�mų=@�Hڳ��ȼ-�<ǣ7�+	�:D"�+�++_�;�S&,yt�D�4��p ���&Ԓ߿@.@P��H��efq���k��< MN�m�N�s���n-~�:�Sy�=瀕�*Q�,������1�v��jR%r�B6��lQ!�1?�r�%�s�t+y�e�P�z�}PwYV�n�#˾Η�y����IY˯��SZ��{!�y�w~�_�qJ�N�M/ y�����iܷ,u���wvv&�T2�tnͨ)�c8fČ��Ӥ+H�j[
�0��H��h(���w<��K�����Q�kx�)j6I�A��e�d)G��:��ܜo �m�' �f��Pn��E.��+���_'E,��k���GX�c�5�_Ŀ�F��I�Nm�-#����j~6uԝ��Ӟ�TS;����������>��6����7���:��n��#r�ګ�k � H��,��P���>�d?���?@/~�_0O~�ѣ�3���!))$A� �����TWךY��q�-QYU��s�jY��7������b�dg���ߋ�����j�da�(��01���m5��M�Y�<�t����������g�H��[K��2����T&Fn���4�[?w��2�x�ǚ�i��s�i�ձu�l2�:�nT�R(�:"Dib�U�BQ3!��оV|h��.���$�ԛ��Ʊ�9^�
��~�����z��w���ذ{��L���g/��򕧯�mwag{u�T��O3�u_6Z�A�Rʲ��[K�PZ&��Ȱp�V#N譆ٰd%QFD�#���{�'����"��%d�i��@��)x�*M�g�ICI0����d��X?��G�{̥A�A*�Fj�ņ�4+�5�P^��X�=A��,�wiԐB ��CR]�i �y��yk*�IpH��E@��HV�X�;�ֲ����dmm�q�o�B�`��7���H\<(ڊ(%aQ
��~F9� @�;��kx�ե�%����#R�f`q��~,�$�dFO�"�� �\/�z�zR�U�L_/Q���u�5�*�Jq��͖��Y5]�.;����IE�/by2�:�Ӎ7嵮'�.ozMp�m�Qd)c��e����C��]D�E�Co�gĬ����8Dp�[I�<��۳$�yk�B����T�LP�׀��8��+�.����ui	�c�8i��{��Bh�`����c�7D�뮚u�]�r�4����!DKm��x^����ȟ��w��NX����KE�����4��Ո���d.����s.!l�OI��MDE�l�@���m��3�s��䒥f�S�%X���������lb��p�:U�D�(V�4u{�ʷ�1,:���L�cd+���P��p����lg��ugkk+�E� w+Ȑ���ňTؐV9(�v��l(���9�G�gu��h�Qv����?\��t�ku�JX�(���;� �y�4=�zvSٚ��NF�$����@OgI��j���Gk��g��cdeH��0Sl�_L�~��G����^h,_:w;=e���O>W'�z��L&�5��/����f�o}�[M3P��<��e�q���#�P�`��3�E�I>��-8󩅅:�֙�/,�X�z��[?��>��K�����+++����!�N�QC�A�0�~?m~���RR)�Z壳|�r)˚������J9ƪIYៗq��@B�U��R!x��ǆPr�!�`g�
��s�>��+إL�̙�+���#���3�>?dߧ����3����`8O��#���&��>~f}��+�
윳g."3�#D��%]%9��o�o�$c�J'�;�wh4�4��J���#�8gg��3L��z�J�X����d�����g��E���Q�3��<r#7���D�A���	�$E��6��������/��s�����&=��.&���~/U���1m�8x4]������kkp'�!mh��?�E�oف����S��������W�/���(��b�'�^W!�������N�ON>�Z>E�:�p	�a�C�z�[��r� ��Y#�É&8A�ڦ^�sK���5��O����RSݾ� ��N�\x��ww��CТ �6R�ԭ��٢1��,�
�"CO�O�e�玅3R������g/!�)�����+Ͻpfq�.gz>͚���ϟ]^Χ�;7���5�P>T"Tȗy1���k��kN���-AM3ĶǦ
D�#_����vML`�Tdv�W��FZX���B�4R�5J���X9s��w�_n�ZO^�|�&rZ/z�'�=�u:��/wW�b�F1��Ғ��c��8i5}���Ɨ?���e8r4�����!Hݯn7c��m_��]w�Z��qpxz}�5��Aa_��<��E�0���D�,�V����y�:tK������½\�֚yS���w7�޹g���E�e���h�zR�����iuhe9v>��Kz��?xF.��æ�ԠE�1W�)ʇO�����I/��I�e�ŕ2\�f�Q�(��!I�Z��O:��}���(��}�(�Ga+�k,-���q3SgN8$����(�!�&��X�9��:gϞ����"%��꯼�
v��85� ��l���~��Շ��H�Q�z��ν{���v`D��H��4b�<�Q��klu�����������r�&aS}��_������SO���}��!�`j�y^2CD�8��XIX�/]�x���J�� �u������}S_�g��a&�m�=��P���(� �iC���g� �-���_�����]@|9�Nz�J6+U���zL�q�2ff�en�s��u,�c����S�U�B;4�'�赩��}���?([��9�����;zN��`-����AjǑ"�s+6������noG�fc[F/��Kcz�`O�����p�<u�T{����Bx�y��L�q�E����G��4�Y�[��N���w�!��v�΃/,���ߝ��޽�g��vfZZ<s�K�/�>z��� O<��*�f�*��+��g,u<^�k��j������H�E�SN%���M���
oܻ#뒅Pf�� B���^�t~a���5���4�����Ϲp�5N��4�ޅ��� l��å�)��NWw�MD��,,�Y�����~�#�u@��B%)����w�f@Y� ��C[ҕ$Y�kP�H�쏭����t{�\���>z��'�� bw��S�mL��qf�3�+�$�sດh�6dFY#��7b?�40��74��{��G�cJ�* �侗�O�j��ڮ�43��j�<�-*6۹���j,6	�;�j ���:b���V�I���駟��}���.ooo�z�k��7�|3�l�C�E�s[P�P�����'S8��z�4���$A{A@ǃ/z�#}����x��Vח�#�ʭ�Ȋ����ީ#���jU6J����c���r���JM�H�~���104�����m��F�GXL���_|�k׮����xz=XC$��V�������>�w��)�2�(��կ~z�&�L�ق�"�x�yn]�w�1�P9�^R�1��(P,iL�Y�|�Igm�~�t���*�C,�&�&�3�<�����{�"�>75���@��?�N�0B�Z+�q��0��Q�I;��)*^���΅�>��q�n�z+k������YkyI{�O +�&ʈs���Z���L4'y�9��]O���t�aw��Q��"p04CF��G���j��Ԣ0(li��
X�{Em�~ݰ��ֶ���a�Iܟ��׆p�7�.�(���p�l��A���`�Kd�ۀsU�!�R30{�K�-P����V�Tw�>����	N@
���bi����n�9�qt���z�5�WCi�<�5Kw͙H�gV���A?��3�tf�������3�X��~��/?��+_�J�®���^!��[���wߏвG"K���j�u�\"��J�%�Q0���5�9C`;��),��Q0���-[���] �3��L����(7��
��%����0�@5BA��P��AyR�O2�fψr��I��q�7E��#�y�B(K,�UgɅJ�?)I��(�PJ�K�S��C[�ú��#:{���s)j0�J���涓��}� �����C���?~occcZ [X�t����N��9&�"]>Y2��w�&[pΝp%|����e�����'��p�y@��e`>�|w�|�:��G/��c��~�[�����h��'�����g���Z�U�Sq7c��_|���W����1��^�H�Tx��52��|�g�2(E�5�_��+������Q��^CK����rxǠ���D�gs�v���:�T�mW��y�	�S&mŪ|0�T���P�E=	P<��)uQ��R<���	���ˇa�,�)%U��D5�YwC�=�yi��a\@T%���ĚOh�,X�s[��y��b���M��}[��kk�Μ�����=|����]��^��;���^���7
;�A�����n,y��2��q�WRV4ݽoem�]h\:}���5?g�;S�\w����{ (��/��Bw�$�,
SX{Y�6�*US6,����}�+�s��]�N�ܫ��q���Y0�4�3��ZE�U�o�4�8!oYU� ���h���޻�>��0�Fr���2{t{���q�􅯼��r�-�^�j���d�H6
��!���w7t-ن@3K�|z}<b��D֚� �!9 �i��-�|I��B�؊��)�p�*��l����59�P�%v�T("��i�g]���,�.zcSY�����V:A��򉝝z�d,�jy��6�
3���&p��ՑoYQ�yu���!?~���?��Z����R��[~�0�����:7��V]"����P��� �E��>�������q���*h�$ϙt�j��y�s��MVxFS.ʠ�?Y�ADnݺ�D�i؈��5l�6�ۛ9:+�f�15��7nܠ&;#������Ni˲�X�zB;A�r�5��U��'�Kց#J��0���D�^��s������_}w�P�
��*J�mk^���?>�z� �*'63t�c��o[>��xw�]p��Sg����.f�p0��aA����ɗ���ߢ�e6�#QVi�) �ڰ�.E�[lz�={v8����)���˞��6d+�$��q{���yRT���ϖ*�$~.�Ps��g���?��zR�=����&nYr�HOΐ�o�cPe���Æ4t���e�L3�����Z;&R�D�~���oG�?z�W�B�y��y�1szK���m��way��n?�u��m�po\�c�/��ښ��n��6��Z�P�w����������q�[M�7;
���L������]�{�ƗȞ�P��D8@����.Bl���Y�{��W�KM��	��(@��8�,�Ά`)@	?�f	�?���&�	V�q�D:�=;�n?��z�����hv��D�3���L��۽�q���Dd���-�,�cbn}�E���&"�Oܹ5�O^�<6f�n�&�8����t|#�<��$��#2ġ~�t���ig`�zR�gS�H]a�B�a�z���A�Wn��kDA�߶m둖�/�B'C�'����0��?�lzI���`"ѷL��Pr�$�D-0�@l#��z�	�b� ��f2.:==�Xo�<�<�j�i�;��rn��7hB�@XY�)ЕH�q���<�B%:D�z��;�e��	��nŮ�,�N��Y;� C��w��5@3/<H� �?Tr����fE�&~1�X�T�?��Oq·��=MO1jG�lX`ހ���Ɂhl�o����4l*�m��	1�do��ֵ"@��oC�5�����AY+ӯR�8j�k��z�N�c2��I��M�
��6Ҕ��X1:7�h�E�Y�NN�� ��l�M̜B޶<]ސ}�=���6���ށ��^젳��\Q��n�{PW��RŪ�4�B����E�Qa��Bͧ�+��rw�>؁[#�_��V4��cg����Ƀ��OӢ�7�OhrYq6���K��e{�cjQ&l*A�wӉN�m��P���n�8T�ŉ�z�9��Rm���'��u�HOL�-ʼ
���^CX�m��ԅ���F�ka�ӎ=rf`<7_}s����mc�SN8����f@HN���h��d2��8�S\#�oOxKz��v�g�>����Ù޲o�6�ݿ����;s�L�4�r�6f�8��D	�q�#gɓ.�+��Ū�pu�dp�މ�#\�`v�'���*{&L�}ح�yMO�(#�xǅ?�p��n�Eq�.�'zaok n�ړ�C��Vڛ��Y1M@��~�)�Z����RK�����y��]�8��>}n��8u�H�o�y�l�s�KO}�O'�K��Loo�}�����(V;���+�֧q$��f��Ѭ��[R�������I޻;֝<�Tl����sg28�o=�����s���^JNkE�kF�g����` 2�EifF�8Á�Abu��.ȉ�Ö���r4b�s�~%�_N��9�S�f]�.�vh�j
Lq�a?��l3�:���%d����@HГ���%zW�G����n��'��o�����A4�5�WFQzγ<�sr���w�Vd�ѣG7o�|����l���#��V� G��փsn?��ٓ� ؏���.E�#t���V3އ���OS��/{� �K���VČ��O aaw�L����K/A�\
@\�l�������It4����SO�m�sɴ;�)���ڥ!lS/-"����ƛ��F]m�AC�!oc�����%]�|y�zN�2�=�(S���e���9��ߖ�z:�"�K�5�{��"�(�HY_R���qD��k�$�Zi�ˈI����]J��Mț��	>��'�Ĭ=9�U`*�z�-�TV����yh�؍�N
��gچ�Z�N܏���@�s�,PF:6��5v���ƣ���ç�T�����-x$��^��dq����j |�'c�&6��\(0I�%
b+��E�s�(xs������t'��qUn?�:P�D��Կ��3�G`��y��� 2�28��	�(j	KgQ�z�p��ǩ-�v����<Si���S��M'�}��6���a��v����~gv�!�7IO�^��W`�y�I����`��[~�k_g�8�$9��&N1�cc�Yj���U�3�s����������z����R��ɽp:ݝZ8�	��`QV�l�#Q���y-l�}�λ����۷� en���w�/~��_������W��ڦ�.�W�,U�3�(�h��Ja�6�e�@>I�>�#�R/7��n��m��R+G�7�F��P�0��1�6~�-������Y�
u�+%�dQU:��ʛ}�,�'�{BV��z�J⹗����zc)�W�L�����M�U�&��T����waׂ�:"-ET�	��� ú.�W��s���[������G���mxƯ|�K.\X��u�4=d����3ю���s4���lU��P��9�NlZLY&��>����WhSw����+W��)��+�k�ȥb����{+����H�J�ZCPB82���߯_�~���o
1"gf&pr�)(��6�&�=[̭�.�狩�MR�����+��sa��Ek.�����V0 ]�����hJ��~�I� 8�)c�C�2z�����<w�sL&:�a�ED. ��q#��l6]��d���׼�U�!A( ��7j��C��2�:�r�Ea#̜�-Mo��Ӟ�L�v����Z����\|�?B3���K�O/���?��T8m�~fg�������E?ˮ8W�!�T�,/��L	�g��.���Hyw6�s��Cg
�پ!~`d�r�%��AK'��[��}�i����_=����)L��S6��4����=y��bީ;l�������R�l�~CG5P�t��`o����������C��[��ک�]=œ��p�=y��{ �����}?������)y�Ą�zq?��I���q\`�^4#�{�
"��\j���SʷAe[G���v ̧�f�4��� Ԧ�q�S��@��~�.�=�{�>��D�m��`6E� õ "T��3=ˍ���0r���e!��*�L��av�����2����<o?���2��-C�-��1IcQó)�C�J9Jj�T�$+��\����4"k�SɢRf�X�Q��e��:�WY%�B���bo~��!�G����/��2�6﮲TF�#�����t��i�S^\�g��]>�8��S�o�t�m#�L$�Y��V��K��"���x}1��S^�k���"�����w�yg��&�T+����1Z�m-+��NA��ESp�������Љ��1���H� !���"B�M�|a'&x5 �;;#��?;��#P��.�T�P�Q��hc������5�P�*I^������^���ּ�؇�y\�a�V������'2�\�@�A������+K�����Sy��u�s�?�c�1�P�O�YA�[���U�$Ah1B3F�f��)z �n�4�Ѓ�)u]X�i;i^tR/�����)�>��e�$
�4�Eϧ#PN�k�<���k�[ÔnR�x�9�����m9KBM�)I��9��f[��fD�kݞ��p4��	&�m��:,Z!���Ju����$�f�eY6;��ͅ��B����j�R������ ����!�1V"U���հ2f�o��3<���EM̵�����������lش_z�������R�L��HQI0#e��8�P �¢s�S�jZ��2������V0�Y�˼.>.��"��6��S��l*�0�i��;ӈ2!vk�.0�I����Z�K�4� � �S����?�*]��N��^L�\�b�"E�J�P�[��ޅ��Pn Y�A1��=�E��w.��d(�On�8Lwb�W���k���X��ao�B���(���|\�ҩ�QP!Z�fǒ�p��,aE�]�
�s�v.���p�E�G�����`<'�l惄+����w��G�$�l8��/�L�	��h4j�_'X��/�ڤU����cz��ެ�mu������ϟg�OpdFx�1�@i���/ B��Ҕ�td=T�sq��'��5��#-�8xN2�F��
򍘮
]�G�;8�	B����aQ �����O��ݟ�?ݒ��饘�w5t`�����3����1Ub�Pm�ї�� [u���	�2?����a?ON�� ��^�L0�䢢s�k2��y��Y��y]�à�?B�����@.2�k�uE}3\��O���HX<�T�{@���Wέ���h�2󌩉�͚`�K#�b�j�Ec����d�c|�d)B�Xqt�ޗ]�ɇ�"j��Ϭ^<����ネ�����vE���=��ӧ�|�IpS�=LCN'c�/���� ��NV=��WSФ%-�0wҲ�^��e�`Jl���j�<Z����ҽ'��\^�B�<Ҥ��:,\hd�J3���;[O�цUE|&��{��yT��������;ON�e4&����J^nM@&�%	>u�pL�JKl=�L1�@J��0����Ȑ�qj'S&v߫T��=!��M�2���5т��A �[m7|�&�
F�Mi79q� �*v��Ϭc����ɞ0g�Lv��p'���X�a�⠐'�+=E���,ּ�cu��n�W?��$�����<��ޣ�� �5n�t}̄�N�7�=�m�%;�G�{h�>���6<��D	�����雋�������_����|�o��^l���!b���o��6l �'��1D�EQ6�F~ӑg��Xr%�g7_�,8���`��N*�cy��<@q��@m�S$�~>�����Jm��� �������+I#�8G����t{ƶ5�i��-���������ܼy� ߀?-�-|v�|ss�IP�[�'�b�i�"�Z��8�nR�7mF-��%����
���9�k�������&��L����m�~�?�yq��^6� Q}��z�ɂс)ǞQ�����IZ����q�y��તJ����[��ï,,�n���NބU�c줱	�7�h�P�_x���x���
��N�y��}�1�<�3</�_���v�T�|oi9Q��
�����Çoݿu�����Dl�s(ʚ�6_"()�d�,��xUw�<�ID��*��.����Y�k9�8���1�#��y�#���������޺D����h8�<��x_��%����EJ�g9"�F��q���82���+ȶ��B�;#
�4d�����g����u��q8�3N&�S0̱1�r/F�6<�+N���B[�p>ts�S��ۣ�!>�}=B�A�|ai�$;��.g͍EG"T�u�4*D3E^D��"[W-'�������A�r�����CNa��x���j�^�(���Ɓ��B�?�+d�� T�xiU� ������n������5�)�ѩ���`��Np��lz��8>�A?rj2{%^�I I<,�R�lk+F�(�^�C>RicF"���Rۻ���%���Z��K�y��r=T�|?Σ><��G����H>�`d�w�⽑j/vA�[���2(_҄�����^?�/���2#/� ����7k��Qt����'��*��I�c̀ K�_��%�,A���周�yd��D1Faш�"	GA�~���yu����9��D�Ιc>����R����*ʘ���H��
�Ӳ��z��k�C7�g�Qfb�k��B3$l�q�L���&x�I:�L':m� WVb�2gϨ9�$�"��}���!�cb�/�p����#��!ݘ���9�%��`:�f�B�Ph��15�p8#	���Ju/1;٪��KA����yg�4��*Ie����C���_�ߒt�V�XeΈG�1�C �V�m
�F�I�I�(:�'�R�Zb�/W�8�kX(O�/6+�˂�-�ƤӋ2,�R�.�<mM��*�	���4�b�I	�]�hR�#�kC��l�*��@���	��aI�<BR�L���Jw3L<��{�Iv#����<��p7S)�e�j��A��:pr��\:��~A�b!����/1Q&�JL����h��O�+
VE��},+R�T�l���̋���4,�Q���Z���?�V99��PWd鏲n�w�'�e6DK�Ƙ�YK}�Q���I٤���� ��?^9��)}�c�A��ٕ�8|G��y�W��[�&ټ�D���-uw��C�X��[��t	r,+����!�'� ���ϔ���YN�r8�F�b�0N�����X3w���݆�[<��=�E�5�ģ�2�Ui��hl\�B�yʳ���9��(	��Q�V�b������z
��>�������>;��
�2��L�:)��+%b<��(L��1�IkJx��<a&K�cd�N\0V�9T�8��1(��H��q[9L���TA�Y���z�$!�V���K�ó�D�j�gtzȦ�#n���e����H�;Ď��
�|��Yj�D�I�|�aZ�H2�.���wuȥ��XHLF��c'�VO� ��X�vqC�7�V!�k�~�rȸj��L/�4(�E���7�㨭�`0��:���c;G-�P�D�PVE��~*M?4��+#�Q�"�մ�xQA,9�`)�㢁3�}i?�Գg�\o�vZ��Fr�p�F��$:VFb�&ṕa*�kL���_�g2�'���	�bV	��V�3$��SL6���S�D����"Q���轠ǅ{Q��J�t	��ʵsд�pU(�=Hb�7�3^⿢���$�sv�g����\��T�:�?��Y��Q���w��e(-1�%�<�MtN���%U}��ͥ5*�E�3Z�Z��+��S;��x̗c�?�����j&\՚�7+{53��� ���s�l�C��C4�\��ܥ��k�R,T�7�R��&�*�F�oc��O<u���%BP�B�1(�Ĝ:���6�ύ�v� >�kZ��o,�����!rݜ/��Z]���P��#�����c��g����`y"�����c%�9w]S��D�4��n�#�i��#/'���ad��7��8�g$y���	�0�Y
�PՉh�D�"��2�"h�"�[)uyym��؊�̪e��u�2��t_9�Z�1,-Y�l����	\�j�q���W%)]��LD!9=��e���u:'%ЅC�r�)�s��c%���<3?"������n.G�~L�g�8�hH3yE�'K�\o�Ƣۇ��L�M�9��E��Rg��0A` KZ�1N�iL����Pm�=��t<�U:Is^v������O�I�.�פ�������/)ʁ��:$B	4�0G��׼�\ {�)j�ٹߥ��ȑ @��
��M>vKu�<$��H'+Y��̃|���:�E5��p�e�A����S�|s�����,�QÆ�؊���X��D�nQ�/����#p%����y~���5Wηs�6='�-0���t F�fw��5m�q�J�2g�x����tA^xd�$��o�L��s��r�������/��륜_���&�JG�='��sL��p֓X!5,��Đ5����  LQ[pԍэ�e��f\ƌ53g�����H]��X&�;G��,�I^���=U_���D�[N=�Ĥ����
%A�"�����փ��:�������V��*�Ƕ���e G�Q �N�b��/ٿ��9�'�h�����|���[��E~xw�-��u}�b��`�A#N��X���13JX୶�ȴ���)�w��o3�o�p�'O"S�\��C$���rs��v��V!�`C��镞Dz_����@��9mM�)�����:�U;w%8��1��8���\PK�1��X?v伦,?X:��>SQ���D;1�2��u�vD�+��w6�_������2����a�2���V_+_�h����e�� �*?D՝�\g�g�T%��K"�t��Ԭ/3?��)8��ի>sx1�(-�Η��4>{b���˳�r����σ�a�QP����{ʕ���S�s}�,ㄜ���T��Ŀ�����D��>@�yު,���
�DUj����Ŗ�����՟�\r+f�N�QŹ��1u���J)����"��LQ0�?f�a��"�-<=��.��^�1���r|�	��wYg��6�76�����HK�98&��L9�ID;ǲ�f�T��	؊���O�!�����QF�U��v����q.?�X�;T3e��P�O98/sT����ŉF��T����2,��N�HjT�!��]A2�S�'Ј{���x�_S*$y��CH���D�<���("�������
Q+�Hb,]͒�L,�q�	d�s����MLT�Q�f��UjIad���4%ŗ�nO������9��~>���b q��8��K<�y���hՈ�|/��i�O�:�)>��squ �arQ#cT~'�497BR�S/Kp�6wB5��{�ۨ���w���P�躩��Y�Cu�͟���#�HTWX�������9�gӤ�{DD0�K!t-/���<�����"��87K,p~Jw��s�e&Π���h��`ο6���"ة\�V���r�J�Qgb�sa�i�Ʈo����ٷ�ˌ�S��O7�z���Kx4��0�{�"˓��Lb*Y�$W���m�Z�)�����E+���J�7g������Ҫ�K��2����1�kOq��
����Nm�T��U,,jQӓ��d75,�oI4���53O�`J��������ҰB�{�.2��2^�ԕ��g�iceQ�xui����d���Y�̶̂t����-�$J�Ec��A 4#�(	u]T��6��g���p�	��=�	Vk��ئ�Iyr����.�f�8��-�����>�A�ǡ���1�L@D��) �ߔ��z�Bw�H"saMT&�n.e�����#�R��Hl]�M��R�jY~*DF��6�3��\~��ݰ��G�p�$M�l9�p{��ȱ�,�D��r��Q�8�m@)��@sΪ��2���Re��(j�+�C����)q�Sɒm���驲�V�j�>wl�<�U�����P�{_^����+�.߹��o}�[��Ya��b }T}�r�v0o:H�8��r��E�1ڣ�ڶ�(�O>{���o|�����~������1p���"C�,}^`?�OYp_���[[[����űi���/���Ν��/^�t�bY;^��������@>�Y�G�)|�Y{V�w�w�t����`�����Ϗ��]���gϵ^t �8H��^|����/����������`�WWY ���I��nf�ϾW"v��7���`�GC�*��0�Y�R�WZ��$����W���1��A�K����/;����<����
�ylzml��q��
/ew�1wr�U̟�<��3�$��F=5/9����幇���7�l�+��$�sA���g��:�Q��x>��OX�U���Sq
�fu�Ǵ �����ݼz�ɏ>����V*w��5���"D�D�_��%����k:��^'�Z�?z����^��vX9K�/k�r�n���W�y睟?���ӧ�Z9{��v/���HDD������,(�O��A�V�777x�]x*�%5��TȻK}k��K+������ׯ�������K�k=�	}�Y�@fq�7<1BL�'WO_��������=ou�_|���R�'��Q��Y�v���{_��[o����v����Ż~�M#4���R���9����+/�K���W��i.w����{����Ǝ�A��Ԇ�@[�Г�J3I6���BE���,V�/�¨�}���D��&���6D�i���i�3����\�B��;��?�N�XBX���־��dF��۩�(�����O��c2U��e�/�[N���*y�W���[m�e�E�`�����c�1N�8��g�05W��v���g����� �t׎���m���>�79����:p�H�hx�V�����Y[q���M�*S��DA^��;��я~t'�7��L��C�^�n#�On�N}��p|��BL�|��_���P���Op�������ιw��1��܏p*>�yD$_�=�=�A8ۣ 9$��%�r*����F��>��7�Ⱥ�͛7�ze̝��$\�x��ҿ���:e��߿?XE���*YzYF�o��q�'^�;��jY�*�$ ��y1I�_�zummm9l���K-�?u�T��<X�4�"��믿��ޏq�>�&D��}ƫ*��(�^�������ö�*�a��x��+B�R��-N$I��9�T4J��A ��n���w}���>K�(؝n�<���.��5�����Qx���<u�wʞ?��ip��/��P`ˈ2��A�������}�=�;�>�k�5} Z�ҌB��i�Z:�S/*�)��V���������.�ٲ�8��w4;Pz�Z��p��ж</��KfI6�N�x�1�^vS���<���Լ")N/�6t�m8���[���u.�[��;�2A��J:\s�e-ǆü�0c�{�.��QSk�^�з����P�i�[X���}�y��z���ܿwccC��a&�AK2��*����/�ħΠ焎�})�*1����ȫb*��䟚�f�BKe��<'w�'���]���z�w`��C�l/,.��~����β՗b˱zm���E��$�2�����I���P�Nӕ�D���1�%���ЇR�Up�h�_�sY����f0�S��:j5Nn�y�g��������J�C���]Hv��S�]�Z,����#1�.//g���;8�S��Ȥ�J���~NKGD�,v������E)�ȫ������ɵ�� (w��l� ��3V*�ݧ�z
�{�_����C���?Z'=߇�sBn����}��~���'��k-F�b4��4���1���j�nٍ0�~M�>v�<�ey�6!|�̙3���/�66*����R�aY�&��ą)��u��P��s�c%zNN08^m.޶ �2�>�������%��	_]]��ᵟ��ISs����Z��^�f��C?�I�{��>��=Wj�廮���N� �Wl�k�N���I���mQe���[�����\a_�h���I�FC�[:��F���(6h�Qb+lu������,��(wvCs4橼ђ<A�15v���%f����BÞQTDp-;w��8@Ƀ�LrW9v��#�bcq3��jw6m�M=��v����h��Җ	%���5�U	�]��y˽�]�
'<��hjc�6*����8��-Ӊ��r��rw8̢���fÑ��M�E�y���hkQ������#�S�4,g�I��
A�����xF.[ݏ�A�iĭ.�j��GzL�9!�)D�ST�8��OǏP}�8?/d��kF�I^�}3
�kPyR
;l_��ۉ���#�<��Ԋ��O�6�y4\Y�nlB$g30?�cEin'rm��j=�g�$H�&Ռ�
'.����v\�&;m��0欯�O'�,iF�u?'��:Z}6��"潖r�U��ċ��ݩ�#�EY������(H��%� �1X2��jg�R�����Z>��`P���>.�ńr���j���.y"�Gp0��k k�:����4Y�X��.�`�r�L�M�9�ǫ%����Y�_-�[pV�ЧFTO���t�b�ΫV N�[����O0�����.l�Żì��p��kc\+NFy��.����m{s�矎<��!�:n-�iMzʪ��`ͩYϥ�e��`s �M��Ō\(��*h��`Ӿ��/�����p�E�k�.X�������O��ܙ��'��>~���/y�ǉ�1���`�q�L���%d)4&��
�n�D%"�#@#M{!��`�ȂSs�]��k�Ɓ�XS#���]x����떭�R ޶Ե]r��*+la��;�vs�
[�̩G��6���UQ�uS<*#�f�����"�۾�Ƚ�sa��(Ƚ��"5SD�'�f�-:�,M�E�H�M͘�U>��O�)Ql'w����m�7��D"�Ӵ�ӃO�\s1 E�� � �;=���t�Gz���_�g^�Rn�z&�`wV����޾�7b� +"nw�v���4�����O�v������0�-�r��TGf��2�
�� ��5&���vL����dl)&F�
�KI�K
�78�L�3=1�w��n�}�tD���'@��n������Gw���~eq�ܹ��Ә�.��sk�3���F
�@����tm�g H��C��ô�.���mA�>��Hް�X�+Ҁ�o������I �A�e�@:]f��N���ˑƱ!�ƹ�w��9����K���:������
.�� NJ�����#����Am��ŶO/X;x�L�V[v!�A�`��G�?#�O�3[6z��׆A���ٳH�>\�̴e�; ���]Љ�Sy�]p� gH�����(�hLA�+����p�3++O>��ým�M�z=�����ZJ$�)�!C�ݾ}{ii	��Ȓ�;��"Mq�,�gG"hӷ�z�ҹsp惝���5�UȲCϕ3�܎è�y�2�wʄ���-!�7���gC
oí�5�
 �joo��O?�9-��ay��Ӏ�Oӻ8	Q`,���A���7����8����������c���*�_�f�W�����O�y��;��mW
���~h�&a0�B̗yN���8�F��ha�AC��3Ka'Y�.7[�n|�k_�����G#�̋�R1�{,��������mY.�}�o��L8o�Bi�ͮm� XV6���,��y�펧Y�|a�y�G��ڢ���G���0��V��!���^�i��z) ܯ�2�0�N�B���+�ǳ0�����ru��h�py	ri���O?}�ڠ�Ȥ��D��s'`G����l>°�Ϝ>��f��7߼������ ��\����I D��hf���P0�AAS�	%��I�ƈ�Mg��B�i�M���N-�3�e��;���:-�����_���4���=��8S�ߟZ)�r�y�k6�5���`�q�2�2�U~Z���m�G<UA�>V�?k���e���9���_y��c5��5�Ix'!����^ +������/�tC,�ɻ��ֱ�
"x��5�u�k_��8�@�~��t�V��-cAڠ�n޼	'��׿��/}�o����E�rĴ�u(W'_]�^�|�s~�ƍ�t�mD�,"�����[��U?��կ"��y�(梀�A�{4�\,�vp6��}���/�:u��"������8J/8��o�G>��_���^��~�N<��#!��;
33pa���������?��W��|}�*+RGT%�Q=���j�W&{��@P||H$��
��(��;���R���7�}��r�����;�m�wge��9�I	�&|%5!Ï�ǈ�3=�U�_�c�z� �^\�\����u������BM�p���9���`�z��aw��mo9�����GxB���򿭞?�?�;����A.tD!gP���F���O��s����_����k�aj�]i�4<P�J�Ɠ���U����-��E�_b+��9?���0�۱l�y{{���g�ϻ/���Ӌ�+�?����)zqچ������x8������ؐ�]y��x��˿�K��4L5�����B�k�Z�O�}���>��������������}�3���AH���]�-�����^�u������@Ŀ���C�,Dx��x�k�F�D����p�:��K�e\�x>�i
�	�e���(��W�+��Ԥy'R2�1|FJ4�M3�:�OzN�<�Q�e�m�yqu��5�Sc�5�����޽�I��5L�T��ej�|!@�i�`'l����)�!����"�N<C�� ���C��r
��I�=����0�k�2DEIxrK}֩Ys;�ls�s]��4"�mOZX
�;a4}�8�,љ�͜��`�y�Q��A��ē7D��q���L���Н;w���>Zk6����O���p�@~σ�Y73��Q�i62�,�8o�|�֭�gPCghnP�pfm���{���}�!�-[�O��d��m!�'c����{��Y�OXP�O6X��z���&�°�W�^O.�g�7�'���+ ��&*�vQ����[gr+mE� |n�,x���$��)s�o��`B\�o;�7��9��F�a��݂��K|'ki�k�՛#	.����Ë������.�<+�\���1�<��+���
��>�c�8�S!j�S�"RV�+ޣ騿��^�Cx6�}����~y1H�Ly��!"-F��--Ǥ��N����v���vkk<ά�R��ChCES�dR�y|�+�~������캰��Y:r&Ы����,
���i���?����\{������W��WR�5�6^� Z�Y���#���?�y~��ga�,��ה��.r�pYa0����'r�_@?��Ê40(	~���฻�����d�����޺w<�M}� ��D���H��4���h���ٟ���O?ٸs�ې��C<L��O�����&=ZP�� ��5�,2��bB3NY��_�m�������v���,߳���vE0֢��V��v���w����ӓ�1чٸI�$D!�VZ���?�X�*&�)����p$�TG���(h(�R��,����cf�~����8ke�ĦT57�w�c�����d'�'" @�'�j!&�ٳgAe���n�w��/�K�\>K��dXC�q�l�b�����?��9����sbi=z��yX_��r���?��"[���
T�p�-���J��nu<���y�����@{-���!�N=�p0\��V>�!�p$���K]�����qr0m�O�W_}���������k�q^Ì�@����g�h>��S�ظ�������1��਩j�׿��v<���w���%k�?u��Hs�"��b��� G� �R�Ƙ���|���d�	�*,/w���I��p!S��T�e�N�����߿��T��Hxe�����_�:&��4��9�?�J�˲�E��sY����D�q�Y!�}��X�QD��54��0�r2I
*��3O�p��|���<@�IM�)�D&yŚ�S%���mn�b���^�:M�.�=+2���%�`���i�a|�֝o���<w�bֲ��׹�{ hP���0�k7��o<�?q噖���w��\��� $C"��,�\���st���9{����]۳�x��j�dm��2l��q~S%���P�����pz=� �zF`�%�w��P����,L����~h��Ͽ�Ⱉ�l`�(�l��fj���HDѣ��q&�\����{L���������n���pkc�e�9#�R��$39�	u�Ą��4ډ����}X\�Wq���߾3��������Z���&�t4ܹpn�6�8�0�e�i��~��r'���Ns��Z�*�(E6!ZIFlX�� �|��YTp��t+m��P�Z�䡌�t�\��˾UB�A�| �Ш��\C;��}l7�CuH~�%?B����7��y����CT``a�e1�!5M�Lo�p8���?_J8�fm���k�nVv�����w���T8���a��{Z�(G��F���{wF�666N=}	|Ī�5+�Z��7���Ç?��O N����eK��/����$��'����Ǹ�Kkg���q�Q�IB����b��cБ���ؐA6P4*V��e�Ĝ��m�����ݻ��^ -���&S��|EZ�Єډ>������ܻw���W���`p>}�c�����y
kyQ��a��`(��mf�EY�S���Q�KuB����II;z��sުjka���ɞ� 1Ӛ���=.�}�?K�
UP����j�e����=�p�ܼ� ��O[���p����B �mO�p�i9�H2P��$F����klcD�ϟ!���8�4�F�Q�|x¯�=��?�
�<�g��#��n���e��H�9h�u����X�ވ�4��
����l'��nܺ}�Ӄ�h��E��!B��M�����
�,��~���;�v`'G� �ib�-#`ްA���uB��4��j�&I�@;6>L#�9�ܟcX;�[b�6��حn�H`��>�pũQBV����y�-��>�Hq|_0FaT���䑃wb3C�(�`Y�6�d&Ϡ��~��GJ����2�}�c�'���@w����Vؠ��)��'1ʪ�=�b  ��IDAT���|�p�{��1�O�c�2O���e�5�i�Ǫ��/���PK�CYP�LCs��i�f�����ȟh��=F����
{�w�1�S@/���.���Og�Z�X��`��*@צW��'N�QӶ�#�)H��b��*v��-�}��s�$8p���pp�׀�Vd�|�r2��.
t�3����>�É^�����^l@�s�� lu���[[\��8�� ��:d�(��_jq�����򐴍z UqJ;|�9���k1��h���#�\jE�D�D�M����f�*
,c!�3��p%�� WTy������ZƎI�;�v&L��0��}��|?�옱`����$��z��P�Vw�����y2���E=�u�����(�X�Mp��,�@텗W�@[C M-OU
kX����c�"h�&�$�yͫ�^ ��t)�b�`l[�øa���"Ղd�7��S7�_z�K�#�a0�m�#��T��Zz�f���=|�&	��_y勠/eR���5�M��`�a��Y�,b;�Xdy�;T/��E3Ĺ��V�[������&�1��i0���fID��7���fk g>�r:��vo��q���$�M�T��/|�߬/�C$ �t���ާ�H�`t4�GTIP䌐�#���4��3J��:�c%��׸È�SIm�,�`��,4P�ڎA�9NTj�Ǣ����N��@���ɉ�gi��6~�ĳ��y��B���3�F��z�cz��K���LZ������{�<����'@�~X��W�?��ys0�{�W�%�`0�¼�� +6����_��5_lpH��e�!��W^�������b�E��?�������ꫯ��N�p������H�^0�A �_���	6��2�.l��D8����Va0_���@2����֭=��<@	n��D�+��n��Js0	7�yx�ƍ0�YO0c��h`3I#��+����m��G.�w~��G��wRL�Lb�C�3�j,w���.�����-~?A�fe�O:?��^%:��e�K'�������e�����pa8�	O�&���d�^8�p��=�����'���i����c�/17U�x�I�E��6��
?D��?v�c/���/��uQ{&���
D��5Z��mG5���S�%{���F�:�yw�:bO��ḝnsf9ʳ�����"ɂ�*�:z�)�'D�)���m��RCo�۝�0rL'H�*��Q�n�4�^�3,��o�4��<�R�����,d:��[D`M���]��a�jy�^�od��4��N�V��3S����Tw��Kۛ~ɑ]wb��s���P�}i���vsD�G�c�f�y|�7������9},�lI��t��4�
��g���.�QРƎ.Y��o����w��IǞ������U�XO �$�����N�Ӭ-7�o1�S�V��W�޵�����9� ���,Ny͵�>�)e�S�3�d�9L�����7�$� ���T�Oa� �+E �$�1�>1&�X.u���_AT9Gm���T��.�M8��-٠Ɨ[ChL�!Ն7��r�z�iU/������4y��2�f�{���������Xx�%����i��7�z|��;n5�A�\s)�eY��!`a+���|��́l6�����0��v�h�� ��Ν;��d���N8��PӦ�i'T1�Ӄ�Q��N4D�(6��f'��zH��	����0=�I���P�w�u�!��ى:_�uK�_{+}����9�9Y����d�c�P8��#�:��[F� C<�߻w��`v�V���g�Ú�2�r�l�WF��["���겠M<Ƥ���$ĜJNYaQ��o���0�oq6{3
_{��o������>IZ�h�J�U�_����r���"wP����L�OFhq)��(WK;5v�TQ��g2�	��G;_ >����Cd�,%޺��ɻ����}+	�V���i�ݛ��D���F�Zjvw�?���U|�i6s_}u/�����}t�.Z�Wh4�:�j��;?�����H֮������͙���M�jΙ�n��"��;[_���>�7�ĝ������oW�����a ,���I�
��1�G�������gA����������g�5 BRi���|����/���?���	:���Í:���e^lMd]�P(��h�~~��忸�M�f��<��KVkp0H�3tV�X]�D2S�a�}�ã_���Щ%N�}wogu}zfJ�3��D� �a���I��8}����JCl,TK)��7��I1WIlZI�l$�G�[=l4d�=���w����� |bZq@���9#`��VD���1�N�y��������a�賋�����+��ߴч�jQ�Z*c��F*jq:`Xv��oHY�&h������吽!�q:a]��᳝4ZO���� �ڍ
���j�y�h� �1S~oTޭ<�.zF(�`Ҷ;q��t�����ϟ��tR�=6����K�ޠ�bmSW$Pp�S�z��ڤ�I��� H����w�v�=H�v�U��6|{��ibν6�OX���!6�Ms&w���3�&|)���U�b�~�Ɇ��	�"��;<z(����0��O����]d��E<3�m��b���sR���E�z�stU}QV�?L���~;��wJ7��Ͳ�ې�U��l��� `���T�c�����!�n�%���h�/׳T?�|ʩ�%.{f���{����)���^+��T{RqC@��'�$ �ɠ�Z��c����n��kfu��<�㷰���F{ecR�������$tq	�I�Tܹ��%;�iϦ��}��bB���HZ��loK�:x����A�A�`�i�ua:L�h����d��K�Ċ�8"h�.¾�^(_�Q��ԁlo�}}�[*X��N�2�f�=�.{ �-xZ��k���%�1�o�٠]��5��K~bx��ml}��`@X-��#O��SE�h�*c�5��\;�>��4׌�c�̬;��֥�%01�(�؃���R�,�߫i�K��H:B=������q��%0-��ۏ0�v��V`�5'�9��q"a7i�<7�zVht�պ�q����52�5`���F��H)(h'HBudJIPywO%��ک�jzA�ՓPb��1~!�>�舣)��>���j��p8_vp��'�˾���c�{T��(C{d�� �<y��z���f�ɸ�%j�l�0����:��?�v�s���qU�!\}AV/p��� GK��^���j�E��pl�n��(fX�90��:(����=z��?< ���蕼<�/n0�:�&W=y�\��#�-��\�����	O���e�:�D�MC��>N�(Z�5�H���(D�[K�΅r{d�t4O�D�K�Ǩ��V�����q��o�M�o�MU���gP)��`I�&��t��[��I����þ\�?��C����E��TjGՊ�7�]��W���-M<Z�{�қ\F��A+��� U�k~���[�M�7;�������.L�;�x���9���< �@E�Ac�e�Ҩ��V,:]�yض֕(�ա���s�j��р�g��sU�+i�dC��+�s��׋I�R���癅��aݟ�vڏ=l=&D"�W�	�m)t=P]H��Ph��u�(&E�W�ZFQF-�;�Xؙ%��#u��+�'�*�Ѹ-P���Q(�Q&:���SJ}��P��ڴ�y`�������'J�X�.�Jn�AIAF�5am��j�F�u�q���V���.NFݧ�CЫ帙���a?��ڼ}��#(>/I��E��m#0~8��Ym��q�#�Z朙��9qu?�[Kkě�Q4v}*���2���2���_�P�i��>,��8ӓS��}�9+Up�b�ǕsW���"��8Ϋu�V�G	��"���r�u���1���4"�k�벸�-���5��
J}�:B�r����/�A��~�|B�g��
T-θ`��K_�9!�@h�D4ޓң��y��`��#M�E������rh�a�P7�3<I�i��"�<y޲C�N����|fff���eyI�D�U�I�A[��43�s8k�� ݟQ�O
oJl������>�H���t�����:-�0�������<|�3���f)G�Y����˩�8F>f���'9�9�G+�W�d�����:��}�tK��1��;�W|���
n&�ԝq&fT�����u��HVb�7��i�? � 	v�r|��0[X��rSR�55�e�Ȕ]h-� ��;$y�� �y�PD9��k�܊���p��ψ��,D�&5��!v;�W('�4��L�E������p�zl֔Z���?���[�XI-�A�'-9�·Hp`LS,&��)���aE�!���u[�:?%H��
�s�Q�kX�������Z?��2栓1f<�:{��;�<<<|�����S�1�fjHQXE`��hb�"�D=�a3��oŶ�˗��?w�ٳ�AoBF�.P8lQ7�O����(��gf,5c�X!L�m�{)m4�gtCǏ=M�(�.S��@=�]Т�����$hđ��������~��}��/��|q.0���s��q���ʦ�H!D�c���a�����N	�ߣ��G���PEIHͲ����]J)ZP�E�>�P��~Q�p�]A9q�JI�d~)��� 6��l�����aJ��V@J�JZ,�"&`�����b�kw��6�=�N�{���b0H�Z]���|�҅�߈nrۥ���E��J��U�k��:��z���f��+W�\{�:|׿>��ڿ�d���wR���ّ���Pk/�˥
,W
,�v��T{�y��J',���S$Z�
�=f��ۮ*}�O�E�1����9R�B��B�&c�,�Hb侔\R�:f����9�6�!ق�&�uEh�e��(F��Ș��q�ؔ�X{s�,#(:�Q���^���t&���z�$�R.��7@g��Z���J�i�����2�D�(yȞQ���Gt�� �qb��h6�����@xMT����:̼C��~N88�l+����
�6�H�nVHgR�57R%1H��Y<$a���n�>a[� i&�A�o%O�#���R������a���?^~��5�1� D>����%j]�u�6.X�Ke�����G:��3L��nh'Ȝ��҃ݶp�`bT�Fmb��\�4Ajn6�����%ϻ�S��	{"�'G��t=Z�,_��HY�S*�!螭H�p��Ab�A��D��,�*N �����vnq0���<�D�D2��|�E��R\�gU�_yϱ2��H�HT����|�܈��V���f^�KSA�8�dV1��)u�8ᣖA�,J�)��q��e�d���q�S&����jY�GV�X��ʐY���*ת��0g-u���G����Ǐw:��0g=MA{��0��_��g���C�j��L��@�ՕUx�~����r(�O?�tN�@���#��Q�`<��1��/���=~�~�9h��*�~k�L>�����׎v7>4�*�,c��(�B�«ģeBg��y2k`sC?V*�Lx���\`�"��a��
�7�{Q�FI%E�8o��e����5H��0\�Z��1�����/0���髬"Y�,n��0��p���+��qm���+c�Vz,�i���V���*Q������q����8'(�&�c羈��#ϗB�(��	�����RE�(���ٹ�AP��b:9�H�Ev��=�sAʭF0ݚD�R�L>���������Տ_��������ϟ��Nd�� �T��&	���S_��kͺ����'���}�YF|��I��eʉ�	��qz��5z�#�����!k���A��:��I7�q�j�F�~'����K*p�eQ��w�QM�z��b��i��54�æ�w��p��xe���>N���'<-Yq�BJ�,��ǫo�W������$��~Ҩŭ����] ��G[��5��;��Y5/�9;}���,GV�S0�=U+�y�g��Q��H���|������Fx���
��/��f�t��������͛7G���%Fؔ�55�Vc�g H�J���Ϟ=�m"A���F"J2��~���Z}4u;�p%���f��ZVp��~s*�z����%_����rR��Q�S����~�Ǽ8���~��j���K�|��8�ңئ��b��b�$fС�z���>A���0���P*#�Rs�E�����0��6�4�ӄ�(�b7O��nŔ
��K�>2�sp��k4+A��=~�υN:���:�U�ۼ`v�"�"x�����Oh0v�>>����������E�ƻi*\��9����C͔�'	8��bp/2j9�EL�>`  ǹu嵩���Q�����E4�����O��k�����{�MTZ`C�&&G���7�� ��0�ۮ��K�}���$��&�S�sB9��hNN]�9>p���������$�&�-j�<��� ۑ�*�7im�KU�'G鸒�;>��e����G�Z!^&�70�1&��%��/����9,�TU)�,����;�}�H�b4�o?��y����>�k�y��0c������y��ǧQmU��a�	�R��ͷY���6�6�7�r�(���\��s�u�=�bɈ�d}�o��y�t���8��Y&��?7��H#r�x�iv���5`����yN��|�FsiiIpM�% �oܸ155u�k�6�z�	�ZX�$-��ȼ��˗/�=��-��Zʕ��	��f�;Rbvd���A�Q'�G�,q�*�Q���ӊ�76�pU&2�U����"8o�~�S���4�"*s����(~ �����)�q��6A�`�^t����@O;%9���.48�ecl���w�%Lz��-7i)�5W�K:����$�)'زUaLh3D':�,L���	B�`�
�~�
���w�$�BcgL�b���d�q���{89�ee��Ag����>]�ȫI�ej�A~��V�,nDa3�K+�(g��pS1�.�Oː���~,�3�����K�X�	���*L��탞=������H{����<����{SS��!h�@�l����~��H�_����/~��W�_C�t0:w�\ZS��O5'��/��+���8�jx8��Q��+5ʲzd�	�� !1�F*끒���\K���[�d���k���%}�g�$z^g[V��e�\����>#'��a~6��Շ���2uQh`ySf9�ݒߘ
�a��O^'�_���ii�xO�1��9�h1).g�K-d�"wb�盜��"r�
b��΋.Sx	�,�.^]�cV82#��Ӫ�dƞl�vzW@]�����3Ϟ={����`{ѿ�	6O,�Ӂ���SЭC�l��g�]�pძ��S�1�4�7�y+���[�V������ܹsg���~�@h�Z @�}�G"�8uR���nk=1!�z>��'�o1^U�j�s����eVB<�e�j>�T��Ŧ�!kzk���J�6�ߜʄ�q�!v�Vd�ݬ�?SJ�R=�'4�Gy�#�dBw�ӱPk�Os��!�o����3x�����4�-���0�(��
�VN"�z�#�WPW1�R���к��{��$��*MJat��q�E	R�}�.(d�Y�� ���-<�a��������L��6�m���B������ȹVV���<L��vR��\G; X�l>��5�9�H� ά�̞�m�V�o=}�K_K�t$m�0� b(j^=����wZ�>��V$��vh~>��������w�-������׎��/��o�>��i��AjON� �������~���`m��8 fa��Ⱦɜ�~|�\���/h)M�w0r�		Qi13��c-�_s�`�E(]YǼ�B�c���Ό58�w6� o:�cy0�^�v���y�R�{+o�#g;��0�`�������	S�>_K���-y�|#�%+>QV!���3��{�M^M�ȳJwF���ƌ���������2�#B�.}�(��,N�T����EӔ��)�S.��H
b����pα��zՙ>s挝a�1�uƠi��p&���}B��b7����'A�ڔi����77A2<y���Q+"�܄O8�m�F�h^�W)O��0���[1Sp�ͷ�r�M5���i,)�V\�$4WC
���n��������?<����/޸�4g���pןFfH7��,ɺ��8����]�"4�yW,.�K�W�Q�j
�<���űQQ��
�QAs$��KOR�0�8�B�B�	�y�T	PƗ���=�J����S��y���$[*]��8�=�D}��~w��}����?�:�`Cx*��g�>|�'pT��G�Ҵ7���(F)�8��0�����/�,�@oi�20(Ay��O�l����7w캝d^f-{��H�z��}d92k��U�G=Jӥu���\]��͒�5�"���V��$���Rp�[��6�P�4�jm�)�i&�_���֭[p�<�{N|��	N|mf~zzZ�Q7H��%C����,�y�y��!�J
/�]�jW��q�9�(\+\/Xj��9�BV0�X�)׮��%!���^e�N��['�{�x��ZV�o�l�lܝ��H���"��$�`��s(k�q1�5�5�>}��������.p��97�8rKi|@ޅękRG����7��0�Ĭ���lcۆ� sTԔ-*���2�H�'��S;u+O��*��U�4�l(ma51:Eb!��`۞�1���������=l�ᛯ��o	,��-..����&��Y�o�a�t}u}k���RW�#YF֫3��z!�x��I��*JUZ�++*V��CY�L�L�!�Җ_��Q�s���Z~E5[�*1_>�So8��1}�O�ȝ,��*4B����/ElV`z�=���u���{�z�s����v�N<���N9����_���?_h��|�M�9�O#����\auh��F�l���$���̮��Aw���v4=�١�̰5��ID�� l;��*�8�etD���ex�@�rc���1ņݠ"Of6{sKe��6{y��3����m�#y���hQ0Х���)�\K"�DC��Y�[F��<��Ν�3y<Vwz���\U�+[:��^��%�<�Z�EՎm%{.W󘏙�S�l��:�������r�^r����d5L���0�Ɛ)��P��kW_k4+++�}�Y,�rv�m*8P'l�ݻw��ǰ��I�Lk'H	��q� ����I�I�C�?�Y�X"f8��;��3Sp���,,'��:N^�)T6Y��\'��,Vl,�Aa \����Q+4�-'`�❎���z3��lV0I�Ϡ���Y֝Ad�m��=����$CD[�\��!lu5��q��0�L?Gj�4~�e��0]�[��L|�@��uY.���KuE@�����J���fI��M:��_����Kia�3X		���h��l۩��+��n��V�>��ʍZ [a�>N�=����������#=LS���ul�ZvU����N1�޵��D�q��Ғ�xh�;��ޛ�\��B����Zc�,���-j��>g��ޒ���g�^�E�S&�)���"?������l�����O�`D3���LE�I��!��DUϱ0+##Agr��:���e���X����k&�L�Sd���_��&/�)#�8׌#)�%�WU6-��UQ��*C=9Yq�'���9y��]+ya%�WD��������F#V��\���7��^�JSX�	�2Y8, ���O`]���v�ެ��x�C��]� �԰�nU�E��Խ��ꓴa^AW���kO�fL�U�R�z
�kWY`�Rɵ�W.�;߷�o~�n� Cg�eR����N-ώ���Ȅi��m�V��\:s�Ν��!�[�T���U�c���+ΐk�+'(0�2۸Q [��h��2�\j�`2�2�L¬�<��^r��[R}������T���:�`�D1��v0cV*O�jF���z�$0���3Ak�`w3�u�/�	����;���~�7.Οs��I|�優�y��9D�Q�KF ��f��|��`��q2�x�%-;��7��<$�2�:n�$���*�j�WQM:��@����p�T*^7��)��Ӕu*�2��A��rq�!p&��*�\��cH��FNzW�$��D�yaAQ&���e
�s&hSx�Y9.ن1yy%'7�4T�9���|`�#)5ٔ��)��T�d�����'M�|}���d乤>���Hm�����������?޽���5��'��Ӛ\�~.��<��A�˿�ˁ@��3�$y�4�U��9*�P�U�� �r���%��W��o��M9���[$]�ڴչN��ޘ�BJ&^������+����-0D���L�Rdl��(�dg7�0J()�k[�0�.�:�b�^�'$я^%�#䳣����S˜}�|-jW�������,ф?�5�A����R�(�mWZ�|r�~��H���Dd�����$"�>�UW2Sy�<#3����������_o�[:۬7���kkka8�����9;;{q�"b$	���QNONyFζ��@&�Em02��ĦJI�rB��p)&��C����(N�(��d�,�/�g�<�HKyЈ"�k�8'|x��(s=(N��һ(_���A�FL����d:������Fs��`a�X�uE@�����؜�Rx�~�����\�Ѐe�!��7�g[Eg{��c��p���9n������X'vё�&�I�g�o\�:+��F)Iğr�K�����Ul>o�����O�b8�awyyyaaqii�+b��Z~���p�`C�{&Pa��X}�����\F��t1������Ut�yvaQR΢�:3�P�Ѧ��葖z����J���� �
O"�kiD����g�SJ�Hǳg눋��(CcE�z���.B���ood����u���;��%"��O�z~YݿSY׫P9;C�X���u�f�����E%���8��"vr���ʈ*s��#�~�����n�Gȼ�,����D��Y��u�|�8e��ᓈ��Ĕ� b��1��ʸÍ�=�x��Z����-���
&�-�^<l;��@|��?ܯ����^�6*Z�G�~�����F+�9��<b�1��X��3%37ø1Y�*��v����ǌ�s.�\�c� �Nȕ�+��q���f��{�V�Q���-�H��R('���,,,���f���,N�V`6;|�#+���z��r*gRc�SF�ES���f�pOD��e�OB��K<��\W���T^�;�����O�9aR��NR��cԟ{��#)��8~D��ܙ˗//,�Ⱨ.���6P�ӧ+�SD��<���֡���?�h��H~�)���N��>�c��i��#M�̦_���vrݪ/�<�����0=����3�jb��V������le���v��u�I�|0>��>%E�wnz�a�8�do1�0�.n�uJ��0��}��/�Iq��hi���2;�tb�;1�K�.*J��^�i��UƒJ��%Bfc-^ʊ3u>�B����^Q�^/aէ�Ѽү��S�H��4~��ؗX�<D��R¯˺��}n?���� &��I���ē]ջ`�w�6�{�܄�=̰+y���C�=v�Z(��iz���O���&�{�֭�g/9�����Ȥ̩�Z<��-��xP�o���2����,��N���A{s(;�����6�`VC'09��7��m�3F������>]!)����b*�V�YW�wJ�f��`»��l��<[Tp�Y��Q	X����.�
}�p�H#|�)[��lK�*}�ק���}�bϲ(�k�6�h .WGW�h�e���퉱��K0Z��DEL�%�Ix0*Z�U�ơ�B�P�ut2����:�ו/x
S�);�b����R�-=\�N6 �����a`?�t:���#��p�츉q�١�������lmn�֜1�5��*�v��ԏ,��� b�nC�hȺ|�X���nG��)��PKv��@��9;%���w��M������N`���z��Q�I�`v�؜�1�[ؾ�e�k�L��|�5��p��I�4�v񒻓�H�~2I5���,㫘#t���c�|�+d�8��Cej��ك	I1�BE^,�`�:!(��p3��V��n%یD�i߁2yp= �[�!}��z0t�d�a~�g��#3���bj���P�ճ:,���tY�c�øgsQ�l�YJρ��ꐛ�t�T 8�/��Gm���N�L�u�P��zI��p�t2.��y����f%�ւ��]�1mQ�0%���Fݎ+=�Z�=(�Ȝ���	���C��ֳg��Z��V���(�h�4rO!�b[ū]�HL3��.�cq�2��}|��V�� L��=%�/�W�e�8\��2W|]���J	I��~�I�q������'�_�~����LD}2�'��{Eu��w.{D2%�i���j��Lp�"`��>�o�J@�°��CNM����QD�h4x�2Y�E�Pv������7Z]:��FX@	"{Q�-egX��@OF]��{��DOȺ�,;vܮ��Ze�����p�	��7&vw@��R��"�I��^����p���I%�
�l������ι�!A�>�;�w3o��8%V���mP��D���w;WPj��ͲZV�(|�l�k/�W��.��^���{�L�0�yWy� ��˪�V�4j�������9n�e�:�v",sb�MYH�,�7��fn�=�i��	�hĘ�� ��`��zݰ�K:�='�Qn,�ُ?�		��Ie]y�E�ةf�Y�1�`�HS���MV�,�NJ�����X�&�[���߆�;H��A����eG*8�KSu.��qf��'���h���)'�|/��|?j@T'f��NU
1-�j�*�r�������)� }5��oG�9Β�y��T�<�򆒻������ߦ�WWF�p�T���PhU+5f<HS8+��ZV��ʯ��(�J����� �u������m�Z����n6��
�gff��C��~��կ��$�ʮ��B�H��h�ץd�w���`r������#Փ�ͫ�K�7-ӸlAe��no����K1vaz�������0L�X�Xe��IFV�F��!4G���"�>2\���y~9��+D���b��r48B�D��;Zj��+,c�ִ�����]�=ִ�s$�����ж�f�`��.4����ǩ�U}�z���Z��#�\F�ɨ,�:���T���*!�%��{c��P��!�7��Jò`�H� ��5��i���d�#mo�k�J��͵�Z��͍%qa��=8�l�7�x=9���Oڈ��h�`e,��Y5�[%w��Y=�/c�X���W7X3�*TE�4�t�2}�hT��V�ݶ}���O��8p�WVV���m�����~rD5,V�L�9v"���S�b��e5̹K�Tr\L˲��!T�DY,JI��C�4��+��*�gr�nr��>�ج�\��<�דo����#B��ھ��{T%�x��?��^���:{�����t�A�����K��
�w����=z 0z]v�Q�x�W�������o�Ҽ�}	��'H����(�C\��ך5'��I���$Q�L,c;F�V"�Pf��;�������Fl���H䀬�Z�Z��O�U�b���I��#�'�H��~��COӘ�O�t&j
X6�����t?�������"O���E�8����T�[��=��w���)<�S��E[�gY��̍���n�̃�a堜y��SCǏ�"#6b�l5 ��΄�eb�++���t��������Z�{��\[�|�Z�G�Qٷ��ܚ�7=�\y��_�½!�-��~�yo�/B��.UG�8§i�N��P]IQ�XJ�P�%d�Ly����0L;~̙G�=^=��/	�;M��l�L�x�����0�X�F�����'�q̲*�+Gˑé�oh��B���ShaL��GU���s�<j&r��e��瘞gʢ�J�uA�?�ѯ>��8�)�ʼ���2��|�]
Y}��l]�Q1�'�*>�vvv�]�6��m���fͅ��d��ӫW�>l�Į����v�/K@��*�w�ت�]��S���9�l�$i�h}Rc�]Г�~bk�Bk����|�����:�{}��3���kdi�+S�&N���I�Ȳ����^���|Rs*��
\��g$C4��X�k�ܠ�Kͳ�*dO�Y�Y��{�j�XEJ����eƩޒ�#�L�ѓs��X��g���x�eU��K���uR.����)�Y��IJ��'F �c�0��Y� Lr+l���!���(Vɍ5g	�(�]OvX#��<�,���D�Gj2����Pu�}#kӵg?�^^������|ӗV ����`�u=&��x�b����ޘ��:�� �R%�`�NH@��EKYD��S8V�X���{��*�yZ��(j.qר+�(T�q�by� ��{����V�%����I
��?�%�������.�A�ӺL�.�oɖ���1Y�x\��r�V%C�X��h��y<��R��{6.Y8�EL�۔o�WK��	�ir(P܏�4�/&�27�Mat��p9��ey�!�2�p�W�P�#V\XI��`�7c�^�I,Ź���>Jι���@I�;w�ܱ�^w��ʷ@)�Qel4h��Ν6���gϞɚ,3Y�+ס��W��;U��9M�����4�;_ܩ	ۭ
MZ�\���ۉ���(rjV,�~-�ja�G�qj�^E2G��IG�Mt=�|�tqg2ð�pF>oQ$���R�B�QU,|��\Z5&_�68�9+X�*���,1��yBY~l��Fő!�=�/'#q�AOzz��|0
Jbɓ�9��_d���	SX�U��� E���Yb�� {Հ~0ه����9X)�p��~_�'�fvH�N�!-3=�����Z�J�����J�eL�Qy^��:�dB�Il��G�/\�+��������$j������E���=��m۞����������~"�2��vy�5� hq��s���ڝ�s�X�>��T3o���~����aA<���@�_��{�*�}̘����L�����1&���f�}��7CS����Y�ⷑ��@R�Z�NM��8�:v�x�*]�uQ�&*�-e����Ӕd]�	3T��9��(�b�s�M��ԉ**��P��#������)D��h�E��<AV�F=����Mм����U�K����|z~�|��1��;X__O�����TkV'e*�}*ټ�:���q�c[� c�F��7P�:Ha��_%<f��VX�X^��NbK��$�
���x"�'��9�p9 ����1��br��x��a"��V��b(*DH�9��y���a�d_�MD������r��z�7���ȡ��$��av��������"eâR�)k�p�M㎲T�܆%�oFI��o)��&�%����%��pg�%��٦��b�%�]�1�<��q.��:�H,�
iI���A��K-,ٔ�A7�bly�۾D����O>�����s��;;1'����8��FbT�lʭ�6G�w�z]y���I�:%$jt,[�G���8ʿ�9z`J�-,��̌-+��y����En���S��R~����p9�t��/�l�u���HW�={�W�S�AS�M�?�?��*�,�$9f$���q9MS�
���>��X�N�<٧�n9Ӫ��sU3�/V>�� �ו���[��e�^��z؂���v����ҙNb��n�Ǵ⇰��ch�u��[�	Tf��$��DCm̰��֋��������[g�6��4��w�����?�skV�����uL���ͼ�_��O`LڦL$lʥ��L5�*d�X�i;�ͭ�([�{�cSԶ�rܠaO4�A�P/�J�5z]9N|�8+b�):��V�/3��$;�ݹ�>Ie��b��f��;����Oe�5��K�?��[qA��Ƌ�2k?D��*s]9�B��Q���*��`-BR�V�, �B8����r�1��e~(�� w�F�����4�m�A7r*�f�M�:	��P��rYD�I���W;r�A8��{{b$~*�5���!����A:D�����k��u���f����LeM[�G80ؓ�^w��/�ڈf����=�s��!��L�� �/��>��_B�U^^
@K����X=��*���Vy�'��8��`�
�ɒ�[T��I��G�QX�N�����(㆖�Ee��B�0�����4�E͖9Uы�	�0:.��xq�1K��(��a���2f�q"da��>A�rR�W�w�'P�v)�s��c��S�m%�g��,( �>C|��F̆Fl���xV�A�2,��\]2��4�+�:��d���Q��C	��t ۏ�q�����Ç��ϟ���;�"��@�aFG)�%n�Xu��@����߿��L�J�S)�Oe�'��X��[Hߙ��A��T��N�Rop�W/����\�ϴq��R��|�C�=���Q��՛n:�d+���Ϳ�}շ�<x��?��"v����_�����
�j�X�2���og���r�����۰�p���G�W(4�w���g�ܸz�j��̻9��؞�u9d�%�jZQW>�-_��裧O��:=������D} ��0x�P�)�����O����������:Ϗ�ı�M�yf	��� G���o��<�ډG��LÇ96�ZX���db|��y����66���>B���	-L�r<d
�8�w�Y���ظ��x��>���zҞ^�q���˺|����uw���1�H���!�M]2�����l��5G�١FY�X��kٻ^�;��աe�ְ���tf���_�=յ����Q�~�֧N7}5�QM���e�<���><��"���Q�:#�F]��^|ib���N]ޠKX �m	"(��9�H>���i4�G�VؓO;�O#� Uf&���ug�W����)�Jm�l����:���3lt{�>��ES���kh3==��=��h}g������C�P��������L������j�ܹsk�!�
2p��bA�lG c�m~���sW��֬M�`?��{8��?j�����|���~�3�T������#�"�<���҅��?|��7}[n��އ{zEF�{86V�K���-�3��������ﷷ7����*�՟�B��x�Q�픊Y`A~��_-?~k��Ǟc�{ۨ���w
�m௬�xB����7���������	�����������z�ʀ���������x'�I)���͉�d�ĝcu�`�`D����*Z1��Hq&I��ɴZ�I�yGez�� �#���J�{��{诹��v�KV�p��7���ʅf�EV.!��d>*�D�&�N�ݞ�t/ ��Ry_�{��y�H�v~&�V[��o�]�;ǂ�����w.��:�Q��ٛ��gwa3;A
"�k�����ܾ�'�~�1�*��ƕ�7ϴ���<\M}�"VfB��ר�gg�xs?l�T<si~����� ["�p�0��I�4L�P��^������fgj��dt&����`Y�2ŰF�E�	=�����oY�;nq��<�w_e��-�m��FN��Bez2@d��������q������ɓ�������-��
C����+���7�{8=����t���b�A<�j���db�̧'�.�V�W4v4Eo�HA����1(�Ι�mw�b����J`��4�2��ٳ[�n�k�O�v}���C ��tGۛq8J����%��7@tMNN���y���X��;�sR������.�:N�\Q��?v�\<�J&��1Ʈ<ۃ��������i��EԀ3+�"A����!W��p��U�'�0����*���?dA�H�X;s���Wძ��?���AߘQ���h�.KQ�\���~��d�����%�B1*6�l��]�o;�o�|kg؆1��P��$!��N�eBg�ƍ��.�l{���Qe]���H�gTg�s0`�⹳~�C·h�QwwȀi��6������:h��%��W��s��Ht�¡+r��7�V/(x�o���¤x�[�Va����<�:���L�v7����}�Ө'3I�S�܂��;���L6c�����$k����_�_��T?X�n�W3��9�S%E��Dp+��/�b�D8j>9�@�X�h#Y�w���G�R8r�w����ΡiG�
���hZAVx�������]�������~|ؓa���2��1VCk����t������m�Z�Voo����Њm��d��!��w��������+WFݝ��A_��p٘B73v�������۟}�%,�R}v����t�0	��&��0?�<9��_����/q�h���LL�����00�O��zP�&��}nj6p���A�;0Q��[&�m��؞�����M���W:J�Xܣ\��2�~�dE[�(\Y�,D�	:�s|'C��.�w�V�&��Z}+���b�5%|�z�Ecz��>��������j�#���d�,4��S#�}8�W���Q/ !k�h���*tNE*��Z�9-��T4	�s��1��ؖK	�*���(S��g���TO�[��C�{�����'-M��]�1B	����'�|�����]���~�.�<[MR�|��_}讠^�Z�A�P��Y��,�:�O�7�~�郈���f�0}Iq@GM�#��8y��I��~��Q��
�	��&�!.H�`��|�̓0�1���IyJ(pC,�t������_��:U��5`�������>�N0pa.e�8� n�Q�M#1�C�����`ɂ]F����'j�
?io��F��V���&��[F����<��S�y���;)��mD�3X`KG6��t@G�b���ވ&pr�I�� =M�B,'U`O��I�1� �]�ъJ_�*5�s)���tzD?�fܲVT~��y��La_������X: 1?���:�S�o��E�յ�H��f�7��s',�b�#���³�4�-�?��]�n�y�`��_魁��=�5a��,����l����� ��S�����7�a<Jm'!";%Z�p����F�Kw�l8
m��V`@]��IL:��=#B����s���s{;��0�T� ��dCE	v�f������.<��:��}������,��+���m+p�����v˯���S���.���:��Ȏd��=�^���z�<NӨ;�HF1P؞Y`�g�l�ڝ��P�z�p�lLd�#v�Y�Bܒ��1E4����`A<5�����LG�`��¯�iG$*��n]�t�:L��tP��\[9nA�d&����9`��Hc{P+��(#�G�rhbO娂HQ��e��s#Wf�Su{s�6}HI�&
��fu�u*��I���&)�R*F6��a�`�wR�
!��E����#���!�$�:��E�k ���.�������&�����&��.P�"��J`��~�^���o�=���SW����+@��X��o-��0�40���Ğ$Mףa֧რI�caa!�������n�;�h�"�\��Ơ/����)�	��e����{Ms�5�7�-�7zT�?ƥ�)G���Q ��Ӎ)���k2c�eL���:�k���v��4.�x0l,�죟�t�#'��ԧ\B�J�1�z�k�C��Д<�%zv���ۊ �1��K�@9E�a**QQ�+��"\U��S��Qv5����^h���Y`�\a�QT��	���냦u��;��|"t��@���04����Y�Ǿq�Zv&���w��:ș�_�Jl;Y/��M,o��N.N_��:�[�nmg��N{$U�pP���&��-0�ݜ�����M����w���%��Z��1/���e��A�8������f�ce�H�����-�v1�%#Qd��Tck�ѹs�.M�]���˰���p�R��Z�A2r�^����zq~�ڵkqgO�x�:����6i��3s����QgS��k��/-^@y�ۄ'�'&�S��t�4�5P��H��P��h8�� ; s��G�~KZ'�`J�J
d�:g��O��$�}�ǃR�U��a8�o��"J����`o)p(4��,vŌ��@]�e��q�l+��v��Ԉ4�A a"�I�3(G�E��E ��b�K�7����I	ƶ��c�$�4]9�?z�ʓd�(c�b?%���م�>����+p���ZF�F�S�rXh��v���׀&f������=Hp��sW�w�-�5>��Ï.]�w�w��>��{��(L�j�fgg������r�ƍ��)��í���D��¦b��Q�������gW��aH�Ã,����AH�^��R���N�^u��M�������߁F�x�.�&(��>��_�r©�����n߾����{!��  0l�ᆹ�����Y)����ջ�����Rh�;�W�֋����4�f�슆'��Sd �h���Ӏ���U�@؜b��G)D�'Qz����2XI��d�8u����<G�҆�E�{����"�,�n1�Vk��4��c��<̍[J��ٺC�U2U@�Q�ӧ�L�m�&���o,����{w������t���}̻uT�3�PcL滶������ [���ʰ?�x����nFI���c��R�k[�sv�̿���8c��}�]��u�6h���zqĭcJ��o�p�^��7�����\=�ߟo���zz~���<��v.4����h�u�V�ĳg�~x���d��9Q����3�?y�C���ý��婙i˱-��/t�A��� 6ϭ�>?�����7e��έ�.�OA̓1sQ8Hah[+-.�=�g����`����o�c;^9(:R���
�tx��G9`��)��D�c�$�v�XJ���t�@�v���M)���{�B&�8�mm�D-#�ڎ)m����� \,a��"i�"�R73N��"���(�@���J�L⚔Aٙy�����	��Oq�s`h8�����?���Щ�����e���R�>|��ɓ�.v�yJ�g�h3��䨌j�,�81�X���� ftPW�d+�e���*�����@|�]�(Y�:p(��}�}F���ݻ��!6��V���#kNx�k38/��o�����c�0�p�������(S����ŋ��O���X�&�]�g))�)P0 ��)��@:=�|>�����!c-���eb������C�-�hu����(��y����	!�9c���
�S���DQU9t�m����������s�0$��a�x��|JO$��Il�G/U ��e�����2���*��$HI޶Ɵ�r�2�F2�즚��c��� ��`��m�v>|���|��<�|u�9h�X��`�\&�'Mc0���ް���֜h��'{����;��֟O�xU*�)	�<|��?���gϞ���,?{���!E:�]��]PAD��_��om=��ûo��v.^�|��_�Z �	�<��N���̙��f��?|��W7�]����.����}��GQ��$�܇�
ff�����_�ݍ��όξy������/X�����(��8��.PZ�Ds��N����}�qk����F���Q�{ӧ��9<����g|�����K.~�����~�h�L[e6"�0�U2Q��ٕ*���b�eA�w�.���a/�� ��t"0���F��VC��*M0ґe��Nc0�ف����hʎCXl;FfiP2Ld�f�ȴUױA[���Ka��$��i9��'���d�!{W4�'���)���r�L���9��#Xڦ�M@y����A݄�o9�;w�Ȉ���$Ƶ`�#`���Y�	��pܲ-�)���8wn4��v�;v:� %�U�2�\Ry�T��3F&�@4�o�|�(�@0�ޠ�t&��!K^��h3�>{C)��D�հ�0�3g�`d~��fF���f�g�Ⱥɇ��av(!0�&�`q,�ا�Ð0�Ѹ� �EI�	���`�L��
v(JLH�@ġ�~��ʧ�N��䅅�00O�>���p ȓӷ��%-��P��Vܦ^��)�6�)��S�2:7?�z����
X)�P�%3y�Ϳ�5v�P���%���SX�_�'�h;���khI:�I�h���BHS�A���Ï�~���w�	�����ݭ5@^b"�[#��b3
]۽r���3g���?�m���j���l����*
.1qdr���s�~��O~��,7���m��)���c��c_��ڭ7����������zm��x�Yg�6Qcn��^/�W:�����ř/��s8]�W�at�"��P�����j���]�~��%�o{��/�4Ms�]�$!��m�,A��7o�<��xwy��>[���f��n�I�>Т���p�wΟ?������'�6G�h��1�r$Is��\��mIּ�5ڟs�,����M�C,-ˢx���d���`����=z�h���w�yw7�w{��z�����gոV�d�
�ߞJp��ȡ�<��h��'v��V-��o,\�?lvRVư�x��p�6*�F99�@EY�v�_�x���O�W�t3tπ�OE""�W
�#��X*S�][� ^�l}�������̈�H9��o@�bC�Yu���u�~8���V��|�&%���O��}>,�S���:
���� 3%Fpz�uYYY����o.an#GF���E��w�	O�;���������Z�:y���Y�+<xjj
�d ��Ȗ��RY�R�q{mF�ȷ������ߏB�jC�a�G}nh�N��6���@1/�v���(&���ׯ����A;��n<�9.���;a;������q6<��g��%34�>YM;M�(L�}�tв(S�9�P������-�&+�R�U��G/�o�T�ۑ�.mqV��K��@Yˬ8��H�ꌼOi����N!�5�UKb����D��6<��sF�%p��;�&ѵ<D�{�Qw���NSr�f{1и�k����Q?�X��i{�K��o�n*IGA���H,v�逈�]�L�#"�w]f*�P��u�P�*�i?^�f��'����ۅ/�K+7L*��&�����)��ڝ���l��m9;������ƒTn��L���g�V�Oz����p���V��(l[��NJ}O���a�����~7	�F��v�f �d��:����a�z�b�e���i�f�g�d�kt|I�ؖb�}��C���یd �Ks�g���f�y�9�GT�j�����}�Y�t�bC��KWw�֓�mm�s�}&�����D-�����9ן��"O����<""x`u0~�Ě�W�M3����ͤ������=�=̛�v'�h4�M5m�����\7S.�li�D%I�Pt�B�@����i��ߘ��U�1E=�T¥�J���wJ���"�s����� �Ī����|@r���(�d�Z�����Jb�c:�����F:��)l����]\A�*5Q�ww7*�ݗ��2]�!���R� �-)4HTt�0�2��d �_,�N����@��N��)���^�0�mXV�������h��O0�����D���fB&5 ��pzn� ��6����%k��X;����O?�d��y���[g/+���O@��H����TK����#�T'>Ąa�r������r�Q`���g�Q���V�&����E#�M��\+:�y��)�4s�ӕ�z��/.�,���!��"�"r|6.�$$fj����ZV�L �)"a=����f�G��C#�أ\�� Ǘ!�dyyR3�C �w�t��SydY��4��b&��A%B���&�c[�;:B�y.�w���i>�`��~
6#)KQ��E�07e���OB�,���_b9`i.d�.����Q4L�ɕ�
qz��� /"0sPda ���Nb��N�U8��1g� �-��s-;�Qo �,N����y7,�����G0�p�m߁3�:={b��~I���O'��Fb?_ST�7o���Ͽ�#<�}p8r��٥�Ý�A;�9��y����~����Sn]yC_h+I=#<��q�"��ԯy�Vc�x$HG-�`�6X�ؼ��e�%��4���?'O��M�-� (���l�����nIݡ���П�ѳ���!1�1�6��!A�A�*���ޥ��ַvfެ�!'�q��7�}�Y�[�[��p��J4�(�ܥ��4s�fϱ�
��5 �Zڱ)�R0�X�e�?�Ԕ3	Q�m�}���x�eif�WsKN�U����� 䴖��}\��&%�h�З~�#Apm��B��uUy�� �a܃����O?�JK(ܬq2�|��zz�Q��Q����MG����+�1!�8qB���$���*U%��=����Lu��׸�$�F�Pn�p�+3T�����H����l�:���	l�Ya6��)�J�73���]��$�/y�9oY2�^���I*�8�=��8���ީ���˗}�6M�ݍxf4��p��_�x��C4n�8u�I.�v�'�Fҫ�#��W���_��O^��a�4�?ո1g	O�ؓJ�*G���L#������� F�ȕ�m�V�*�Mh��3�=�Rӌ�B���-d��S��HPH�1�
ae����O�V��(4J���Koaqix���U��R(�8��ti��U��D	��!�"h��ڰ���,KLe�s�:���9j����$��(g�p+�$D�$&���˖")��S�@>��Z�Ve�y ��V� ��$Q.c���8׏�gJ�h�{eF�rB��~��&il"֠�����(U;����X�G�J���C7�]�&3#����_��B�gui���	�g(���:�����~�pD��v���9��v�zx/vF���:]V�B��+K
8����G4������N��$6����j�><����q���k�r�����3�:ol���̔��1Θ�� �|����qC��6Ƭ���O��W�t�3g#�T +����IIS卡�K��h4��P��M���[L���0QxZaq��W2�2�bo�3sn���̀t�E^�\M(�f5��v�[TS�DN�������9�T����F�S�J���*�4]�I�n��op�Z�
*�ćR2�=,�4�a�~d}Een�uq*�=�CY��BHx����ַH�7�W�\�=��5��p�����t��Q0�'m>�pT�L�����vv�lHb8�M&拑-�͵��
?<����GXh�k.e9�g�%�T�ڄ�hl���Y�~�w_�ܳ�fv߫���wD��@���P��`>>��WH�Ɏ�U���[��,2��n�p�A�6$=M���M5��uadt-�1����,�n���+�hF����8�j�R$�*2����`�Ed�	�L�͒yQH\��}�5�&�^�\m4���쵪�����4�e&�p �MT'�=0��m�:!l�0��PڄlttECs�
�e{A�I���g̶Zr4��U�I����%d?$���Zs�ǋe��4����<Ú��$ Ims��1��3
7u�s$\l���lּ�me�.��޹�@��cK��~@쀮"���ֻy���_��G�EfRV,5��Fc�kD];:uj�R}m���'�"ZEb�c�:|��(�k	��t�0�^���Y XuP}<?���Z�[X\��m��CIgQ�� ��2�V�ؐ6-�Ц�G9��M�����I�7JR ͠^*_en�I��".SU��LS�5[��E0}�8�}j���]��I�@�������$i���T�q-���O�k�`��@c�Ѳjڎ���<9�\+��i�Y�cMa��cR���-��07K��\i!�I�y%�!b3������]��
SA����L�3.4�Vw:�-�;�[�RQ�0��R<��R%yӣAUZ�O�I|'Y�G/&Q5*���?��ƍ˧�!Y�N'�^�v����F���?�5}��1��s�x��R�]S=y�_a_�ԭ����	@ҭ)r3�z�-�G%��ippp@r�si���5��z<��MJ五��7�^����'�~�TǬ��sss ��iNbE���LB�z�d�^Tn��%t���߼���J�6�Nw�4�'��b�ݦh�����~z||����\�ꮡ�F�)�S��ˠ��2߭�v�%�!�ak��Y��Ql9HcR�$��0�d�҉���+r�ly(�"QA��1עSk�,�sa�VQ�S AE�z.�V�)ꋭn8 ����1ñ���yP�Sx�K��FI�|�ƻ'��H[rb�B�X$!������j	��,�T�eC��jC22�x�Y3]α��c���4K/�z��kQWCp��f��2�K�U���~t�t�2��?X���~^��o��`�ih������K2��!d��˗/w�h}}}nqauu���L��H�壧�w��E�P�H1��dj��%����������w��pԚ���+���$��O�f���F"��]=� Ȓ5��,�Egi����
�tԄ�O�a�(g8x�;sFު7��YᜢT�cbG�Md�����$c�{����R��������:���s��,�q3�'4�ez��腅:}�/<x@���j�/^����#$E<O(0�[��Ky�]W���;ǄW5���k�i����Ī������ɞ�������9Ʀ�g����������8k�\�RȰ0M���<�v��?�̙3�\-��h;AJ����8xs��z�V��<����-#F�~k��$]ѕ��#�D�D�W��$�\H�h�:s��N�ui�mV���ǁ%Mr���^���Fx�7����^����d���=������#z:��u��
���U�̬=��=�5	�o������&Iest5�F��C�"p��=�M�r�Ŝ�T�[)�j`!�F�w��	+�8�J!�� �j�`�I���sk��l��ׯ�]ؖ�:�G����+s�ߕ�ʃ��^�Fg�9}��._��s�<�����E�b�\s�wNk�ۺ��yR&e�����d�RgO�*|��)i��A���o&Z�l1 u��Ϣ";���W
K��~��A	�Z��`a)K��%�e�38���������6�(E�!;@p,c_l���d��Fn�)\E�[�ad�&�[Z5�PxD��3����=�)k����`��Z�;��'U��\3-ֽ��ͣ~��;̢���yW:w8�j ��M�$�G>|#A������¹�LW�Zeo��K��3f[���D�/�[��(2Y�o��n\�|�������NC>��V��|w�U>�W�+g�οum�\���t��T�]�f���
a��څŵӫ��W���OPL�Y��:�����"���Z��.�>����zi]��<�����:tB`kr�K�)/�����W���?z�W�����iq�,�Q�+�Bz���h�q���������>~J�Ld�*u�4��g:�Gi����s���T�y���'9D6;�î����'G�	ӕ�A��W��;7�YYYvc��J�s���z�j��O��Q6R�H�n�;���|��)?���=~YM�$���Ɠ���#Us��٫/У�˽_��Q����ԃN�M���f�?��w��O��{~�� ���JU�B���sq��իW/]�B���ϐBXI�'�8Y��!��n�[��ћ�Hhr��������r
)�E�ޖ��G�w�QMN��O\��*�̑5�����/�B��=�Ju��j$�#C�?�$Lej��nӀ�D�hB����2��H-�hc��Q�sz�K�.)��`�Z1i~9�d�*{q�������� ��C5�5a�+!hw���(H�o�	-ak�L�?�����1���wy�2Ϸ��sK�u\a�N����'�v��C�"�}�\��[ ]��`�v�G��0g��6���[a��;x�>x������_������>���I��#uജ%|͆f�qr�oZK�~1�����'O������l��Me���ls�,G����h�ִ�|����������~�D���#�Q�[����[���wiB����띇w�W	Z�'ܲ\�Ȋ@��ǟ�z��y��R�>{����EPŤtn9d׼,I�I(����#�����i����';Ao$��FVJn����a�O�����p�;u�/�tpԻy�f�7(@�c�MQEO@�6���y�0�MU*A˪I')ݴ�|�=�њ�lB�%}�3����V�#����3�D��2̦�: �,|q����;W�Ө��n�l�	�ģ��J��w7�m��C�n�3ҡC�U8d������@�X���kpX�(֓�Z̼>82�x�K��lq�"22��$�_Ꮭ:t�$`�}ojG��E��R�t�U���Qc���~�3��$*Z�d7.��*���<ԐR��p8��b�+U9�%�f����{0���¹o!�m;?�'-6gF.,Pu�<鄝�;��>�eu�Q��A!��4<��J6�GmB�{x�3O�wUV�-F���'�Ӧ�>����;���\��ܪy�:�reP�e�~�)��\��B��$}?f�s��&[y�J����%^e���#x��D	c
����K���}q@���-�&xq��A��Li�;�T�+}�FC�۳L��9D@�OcX��Dbx�2(��cf��e�t��x���H.(��Q��l�IsL�-&ha6=pv��!�c�S�_��~E�m*Ø4}G��O	�]����6��ԝa���V6�K+�Vz|��Ξ����/xKC�+�ѻ߼�x���緞�17���JYlfWӂ$��Cf^�vj�S[���Lr!MBɽ�ހ��<>��u�;Z!�R��*/,.}���5<l�����J�<�
2�{y�Y^*���e
��i[�0��G�eM1}�M}DF�.��A���g^�g�_?��ݝ�ݐ�6��W�����s����Aq!���cFZ�H
K���z_T���1�����h�N����C��&`�z�Uy����-���gF�]�[NXEe�2�
�0�ʄg`��v�9t>��)V����;{�8h.�v���m��~�OF�1����� �ӭE�K�Q��ɍ��{蔆'6�ǟ�=�3Kn���O�w���9�:�zi��zy��AR��21�"�
:$U)���
����'��ȫ��9A�� x)��ʊ8�B��HC�'�j�GMg�x���2FH�i���o$b���1���PY��Ҿ�����q6Q��2�TГt+x3�Y�`+�V���P}��0^I�U�0SSXP�p(���,]���VO��@�G�-�qȘ��X`����"�����v8�U��q�s�=��z�y��RЄ#|��"!�?�`B,+�X���SLZ𽘐�:�'��[s-:!��MZ�c�*g��n��<u��DX��st:
iB$�PLd*)���5'f21�$>@�&��@�V�Τ���ۺJ�!!=�F�f�
iLA3�Iv�݃F�X;E�"�BϮg��Bwi'-z�¹F�X��j:*��&��s��Q&f1m�ıs0��(|�3$�>��=͍*��XUe�{���ƙkMo�/W����ovww{u�����7��k�O���p�u��*�#C��I
�j��$%����4��(��F�I�Mɐ��p���a��� 8n,�2%i�c�Ib64�ҵ�J!�dW���!���Ti��n #R����%�����P�)��u��8􎅳�W)!��j(m	�"�0%<�����z7v�F��Z���ep*+ͷ���l�Q�6�l��=g���b�	j��|�Φ��t,�,R$u%46S��˨����Э�˴����O~̀D3E��J1.g䮪v�Q�Dv�����/�d�6k�3��~UR��s��f��QA���ja�G����Ե���U�U:�����!�׷MX�Fx�f�]�U|��c�2v��_J7+��E�pT$�ˍ��5�P�e�q�-�7+4R'��B�]�RQ�gR<:�5L�E�9ϙsę.���>韦O輦�-g��O�}I.4�u�n4�F6���t� 	쭪I(�.�TD�����nxغs�J�P��p��Rإ��?�d,�&�CW���5V��K.��^�L���+H6R`T�&��k�:�/J�� �aP�xR�<᱌+�5v�p_���{QLoئ��wT	�����Ă�*�4��2d9y��3s�HC�ǘ���l18�C�OՖ�L�7�|���ۏ���d��,�E���ׯ������8��P5D�@
]A W	+��+������:Ĳ�OHp@m.�A*�{G��y�
N����W��ҵ2-�T�yU���"�8��<�����򲐛/��z�
�Ko_ �UϪ��9EZCK"F�;w�!�W�g+�[�xs��;�f6(8�c�I�׆32s�҈�H��<X�E]�NRą�c�9r8jq��Ȋ�<BV���ts�j������ƴ�l����b��E��ü�9��e��g��H���C��a�ia<"ǃfф�	"\D��hVYai��ܣ�Qݯ��!#l�D=����+��.��k��\���Q���l�kb?�|�q�~��̘�R�Q�B�.�h��\�/���/Z��;�n�9�C#f��q�j(��x{sg��v�bf�v�[���#�&�p��-���e��8��*uh���������i$�8J�D��J�R�F}<����}�^W��Y.�?�5�_�W�]M6|�*3=���Y��5�:�i{{U��I,��&Lf"��~����>�y
ʺy����y�����@W��=`^-8�k��gIS9�x�3�Ÿ�'cc �-UƎLqv�����|���+'���/���_�Hı�.��&f�^&�?�:���d;�@������˓�P��Wu'�z<���~���*>Q�Y��I'�|�q�¨P�v���ӧO���i�>�;!~L�����%�{�n?}��3b���W,�P����*w̖2�Z$'ŭ#�bK�[���X:l9����fʟW�]�����(����$�xZnn�����q�%��ӴrS�pQP,�umy����,-�xq	�K�Y�,\�x���t�8Ib2RÅ�ҕƺmx��[�O�y�VV�73�>��22��rd�X��5�^���^ ]%YeYKI��IIw��r�-�R�ա(XI���Bcܰ�y%Rܡ	p�B�Y^╱�(5����{��Ld��� [
5�d"��d��l=O��$�����ܹ&s"�Ҭ������gSqŗ@���]B�Q�kɅ*.丝��p����z��06�H�Q�De4jѐ@Ήh:}���-7?ݻ�����<����o~SK+)��#��ೝ���ppxxXyV��*3���W��;�I��h��:Fd����,�Lj��F��	]�Uk`�����E	����2q�%��������OV��/����F~�k�NW��4�9�)*��y���	�4݀wX�:������������H ����,��J4�8+m"}56���N��l�0QlJй��C��!��y�O�5���,$&}�f��s��3)�J���)rl�O�d��'��$o^EW���N�x�2i�G��lnn�M���;�~��aL67�����_����H$�Rgj��丯�t�ڄ����7��T��=���1P�"��t�^pZ4�q�}���J�5[�bH��bњ�E]23:�t0�8�$;��H���i$��Nf�����I��"K5. t�����&��\@%�S��d�+��i؇��ƥ�� ������g�Oѧ"�hO�Ck}}����\M�-,����YE�������5�zVD�PB�V_���̊j�\Mk����h܅0n�j�"l��K$SS8�j�I0@&=�[\ۯ������@�8�0ҟt�ԣ�!��2*u�3�u�p�9O��s�A?*�[��h�����?�ЯY��]k�i�ֲ�f�FU��[�k�%27��F��ȥ�J���:�j���j$\#2:��ͮ�t-3��*���L�RF*\%8�A7�*N,���E�lY5Z��б����˨׫b��~uH"�q����C��H1��+G���ÆN��f���
1P�̪����=�J[㝭x��.������gŴ2�����oC7TҶB��>h]o�P�R�}�;���f���r��?�b���x��B�Gt�{�g�,Q��]ZlP��l�8�f�a���E���O�
#U�`�v{�����3�+�}⇑�:yu%*���DR�P2�����Q3��� x_�C---�N�_z�HV"��k$Hp>y��`�ƥ�h2�|���ϟ��AE�GUR
eZq�Y�*�3 '�x�g��6��ЊGaYɀA�����I���y�N�A��08�"�V����Q��U�r��Q�ϳ'-�<(^�*�WG�����ə�+�\�$*�A�
�tee}����K�R�jv����ʔ�QoX��#b�fS74en"�(O��|����9e�¦4S�E]�[�t�c��a?�C�%IG7߽l�_��6e�b3Thb`�I��O����@��q���°h��H� U΀��G�]%���
@З`6����s����1:lHO�ee�(`s2UÖ�*�%�)��cD�>5��S	��$OK����g�DKjf67�a�os�R4����w��:�޽��	�����k׮������_~t��}������|pz}�ը�͒ �7Ҹ79	�,��BM��ͪ<������Y\��JtC>��gy֯2RO�Y���"�Tr-�7M'��V�tUš�!5;`�3��z��$�� e$%���%����d)���b�l5�C�C���H��b 6-���-�ꉮ��2z�����`���=m�)��Q�8�C��#��)�=��W�G�/�����q�I��!��N?}�dsM�К� ӂ��>��������U�A��O��d�=��\p:��N�PA@GCR�8�͚�1i�njcT	Z��y32]9;0;���L|����TDM���y�}5%�`�N��M�yjߔ���B��o�b�fT����˱�B��$Yl.������?�;n�l��7n�Gs���3������i߻�E�7���H����E���ZoNb'H�'�I�����`~z��2e���E�g�!`�a�|R����9�鎾�޳��k�ѷ�Dd|&`_G���Fu�&��ERp�i���D_cM��W(���fl��� ޕc�X�jeS5y�n��^b���Z5=&�����*��+}��%�)wG���85;
5�TW��5����up�qZw�Vf��5�(v���3g�J�bkt8���Y��"�U�Mɑ^�4�5C��h�\��� $n�lfaVI���|Y�VK�\��<ֳ&cn�m�/�ƄҐ���[�&ź�FTO ����=z���|�����b��,���١�(S �����KC�4�lܽד0ݬ���b�u�=(Q
�;Z���Ui1a��@��G������a7�2�¥������y��Yr�Hɱi.WYw�r[6�s4�Q����b֞Ƿ�4r�r�9�R-1n&	>�u�R�s���>r\#4!�=T{`s{�@V�
��U����S��_��ϟ����݁?䆔9J���OlB~��IWAF������B��BE#���S�YN8$�j
��k�R΀�IP��.��1]+�_�/A?��M�D˼���tj�d̒��'�L�I�$כ�5�T�p�����yb��RJ��Lq�+e)�x*//	B��?x� �H�iR��ViΨ�/j�f�+Q��V�Z�s�VaV��
7���S�H�,�cG%�F�썬D��d�c2oeRe�Gδ^���b*�o�<�QUK�Ȟ#��F�a��wx�'�5	�Ҍ�lu)����T�x���dN �PQ����(�1����uA���P1}Ғ]<7�b�&?�K_^^&;�5��|��@�"��X.�D
ԗ���	B�r}���Je4��`3�Y�mV�O_Jf�q��[&��s6��|8���Y�2�ev[��=��j�	�48�Dr�nހ��B�Y�*����`�6g�ht��gߪ����z���<��O�Zs��ЧIjd����B��kK�����3�J�c�趨eZfX�iv���L,Qb(c~��k��?��8b�UR��oGy��~ 1��B����C55�v�˳��/F�����G�1JѻP�����
V�rLO�Ęމu4CL�Hq5��Q�{��^o�A��ͭ�~|���F-�Es������DS��S�\IU��԰���!#����d� 9ϖ�\����'��Ff(�w%
���t�"+�Ƨ��8q^G����죝U	N�V�1G�.3��#��#�+���y�u����֗�]�Y�H!��7������f�lkz�P����a�i�WV'l�x��#S,V��W��:�r�;�8{��M94��3�ѻ�OT��������G7n�X?�����6S����ٍ��t_�x����`(��Ob�dӶ�j�b�<2f21��B�?N,D�R���\ç	����,��|�C�g��4�t�Fe�D����ZV�4j��|v||ܗ`u�㴇�xÚcH��R��vCvɦ��7=�z���"i�b|��$��b�/�[���~��;�؋L��?�!N`�g��G]�b�R��꿷o�&��2�H��0b��򁤺�]�'������⿜�H� c�SF7�M���K�����M��b~��|c�A�u���4I���B��:��tW��R�f���:�W/�����%ꮮ�f�t������h3��_�'2~���PH�H�82�N9sr��n����gOR�X,O��*_їV�fE),��r���uo�E;��pk�>ҹ�Lrcc25�(�2B���F�	G�dQ�ɲ"�^T.��h�q�w/�=�Պ�:癸�4���f��5��Q�s͹���>\����z�n�����6��}|7k!;����*���s�c�H�-�<�T�HG�3������|���K�6\C�q�Ӻ����z�Y\\|����!���Mt\�����7��od�ʱLfx,�Ҟ��(�eH����k�Ò9l��J��V�q	G�R�#Sp��q��tD��$=)M?���:��C�{y2}6�(��q���=�3/�a��Z�`f�(=�X.I[Eoɤ�����3p<89',pφ��bd�Xs���;{��G����>�5�zT�$���UL2����;�r����W|�K�U�K������WE����D
\�eIP��x[��R��]���ٓ�,A�#P�Xp���dM̞<$#-��"ȧ��qC��&���]h �-�1�sM)����'�q�dZ����T�Q1y��E�� ��3�`�_���I�va�r��Q����"*H��.9���3g���׿&I��U�t���	���.����\C��SnB��@uyL96��+�����Uu\s��z�eye��Z�aU�@��^0W�/�����q6���|�ota�	5�@�<�����L�TG1I�)���D���zy��&�7	{d��:���Š7�11�|�~��*���%'�*(U2Ŋ��d����
9�f����G�L�l�L���q��Yz�u�B#J���-͇���+E�b%�[^�ĪK�`��"�d�Ԙ���I&��#�z�բ���U����n=o��Nڥb؊����aI2�� cFOT
�1�vX�&�Ys�,�,ᖺ�$��m%Z`��y;��[=ٳu3�C7�[��[�a�hFP[y���B7`�§Qϰ�S;�7�eմ�yw/��3�j;�_��g�������wF$J鱲�t�Q��ۇ?�M\�)}���_���%�s�7�$j�2=�T|xi����{��W4k�X��5W�g���{���0���w)Fe�1�E�n�OS��-�,�Ef���ڠ4�Sȳ/bt7_��������K:XR?���XZ�s廰��$iP� Ű��X��+;^pL�(PU4Ob#3��n]\]X*gA�9�1�A��W�#�%�H�2�y���f�fs>�m��\ CS+d��cH���JW�O�ӯ��4J�9ǀ�JU;MhZK��)g�)ob��rM�2��W��a����^5�*9�xJ��N�����HIG�m����K��UѲ�jU��v4ը�v����9�.��2�>#��������aG�.*�vb؋`b�?�҃�E�O��-����s��� ��֚
"� [�:�B�'л~��cx�U4�zt�݁>��Ƕ��$�})/]�t��U��᧿�>���"��S�N��$�W�Oת������!�X�V�� 9�2gu4�U���0�#��׀z��=�bsԤ��>��Pd��w�d9|�<x��Ӈ�i>C�Ë:��2�Oa��7�6�����B��E��d�>�kHKRT�\��^�U�������U`���{�QE�C���Af�\tN'�K�TݴH�9�hT�^d�3u���e�HҘ�S�5�mXt���<pq���*&�-L�[��>�rmj��+��xqs�+ၒc+'�d3��p$�_���"�tO�V���,+J̝��C�-����iz� �Q�$��k�\�&�M�%�E�#�c�����ʫ�,�붳V:�z��vh<��s����"�F,)Dw���pW���D2_K	�fbE��uZ�(o��峗��ƀ�1�`O�rPͯ�K��Tg����$!n�~�Y�Q�nދ�7��X߽��k6O�]x���O�-Ш:�����������h���8�\��8�a�W��6�gK������-Z
�J����i�%J��7._9{�XYY�-�͵��v6$����}���&��]^�P�BBtP����?�6@Ɩ�8��OF��=��U:1�vX\�a�q�t9,��%�Z�q7z���V_m��7�,��	Z�/7]B5�1� V>��W�kH)�TA�<f�+&���;
Ѓ,Dg ��K�h�$Iα�"�W��JX�"ƒ��Y\6v���YZZ:����_cg'2Xl[��v:�v
�syjY��Y���x�ꬃ;��%��mҶ(�l aZI��~��"���v���]a񕕕�����drݦ�zM�@o��k�־�rթ�_q>���3N.��ѐ�V#(�駟.���
$i�}�Y;�VSY���.6jt����"��*�r���8�Oc��T���y��r���Sq���#�n��Z���������C��LC���(�ܐ�����t��9�,u�\����ݚ�erji�>�p�1D���L~�����K!�x��f�Q��3=�UH��ҬL��MKsL�c�{|����rXjAV]det�<�8��U&GR�p��sU�%��VEU���^�'����7-!�UfW���3��d�J~�]S�?���q�j}���s�K�皖�u���ޥ���0��ZV�Uv�j�6mV�\��d�L�X�Ш� cZ���JۯoT]<s꭫s�*����u4t�3��p�^m-��w�����Âz쬒�.x��ԤYi���a���`�[�7f-V�8�eЎ3�ekh�10L�B�g��']�H�5-�n��vY��s+���Wަ=do���烧��gOO���ť�N�P�n�G�&�w�U���gh�I��V�!��f���y��ײ��V���#d�d�$��Yz����拏�/F��釉�����7��ak�%�������|�����B3K�n��	�y��?��K⇽펙8apl)�]�
�RH*��/\kI�-*U܃����/�,gM��~�O&q�qb8�B�Az��N'o1Az�-�ߛ�'�;+�����@���m�����HV}�˨c�A:�|��ݻw�/ɲ�G[���ᙉӘ����[rքi4�����#����&9]_vH{�6�i�HFҐ�.���<���/N���?˩_����a�;w�{�y��,�_��؈�mz�@��O���몞��&G��%H4'Q�l����/I�%Fa̱L25�?ڌ� u1�I�d���;�[����x��`����C4�4�4!�G�����T-��U�*��*�J��fF��?{�Ņ��"�2P������~�������YY�E��t]�$0�&�����i&�Zz����T��Ƨ�z��D�~%�D��/j���&�>��UϷ��?QFM�����Ku��n���;Gk��\��.��tT7��5��ৣ�Ov�:Z�7��[r�S���Ф�{�����4�7֯��[��/�J��{띫���{�'�H��t��L3OZ�#n����SM��<R;�v��+��o��������[��VH3�>|����������-,@.<��D�y����	9Y(�0@�`y�3���ˋt�����<l�Ss� �˗�z�z?Mų;`�c�χ%��c�����B�`��ۨ9�N�G���vO9��LG�L���u���w�{aa�6�b�L���VO�4B�%и���r�G��%9~��\}q��tqc���(�6VϜ=s�ɓ'I
�5�"���p�V�6zIO����r��T�c��)���(i̻� 05}]1�0���i��O�=�����Uz�����Lx�2�]@�^R�D�u:)
Ȱ<z��u�/����&#1�
�2�G��n�*#U�`�ڠ+���Z��j{��K�d.����;��O`�M�\�I�5��"R$�ΊE�����}� ���5�+O��_?���;WѨR�\��ʺ{Oa�_=u{{��I�����eo>���ov��~���Z�;�*-��WG<}�%<Q�}��	I���gi��ٳg��n ���ɹ�ѡ�ʙ�M�+��6aW?z��g��0�)IBR�`�Wsi��4����>�^J�a%Nܾu�f�wI�3��! ߹_G�[S����;ή��S+~@:��ϡ76	z�4ET����r%^�|����U�:��ƭ�P�B�e��̉,��Bu��I�=��]�Q2v$gAӊ�Y�M����W���E��Ϗ�#��AN�\_GJ��J����0��L|��ҍ���[|��N�>��؏��.�q��rL�0�8�LK��%����U鑬zi��d����_ܺu���߬���M�2i�kz�jH�%��4j��X��l��҄jA��L}i���_��\�xm�t��	�c� E����L:~��4Ӭ�m��^0������� /Ȍ][j��������^<ݬI�@��A*�z94�|�Y&��Z�Q��� YϽ�N�3h�����I%�Ņv���'����nhs��˗� �e�j��58��$�w\���~7y��:݀��� q)}Saz�27���i�E6�������X�A�3�t¦y����-�8;f�:̭ O�ǒ�v윔��G�4K��tk�ً�"n�����#.$��bӐ�j�N"|�U�)�K͔aخeښᣒ�n��U!@N0X	�,]��(�,F�V���Aٔ6�`8
\]����˃��|H�����'�2M|ǎ`^L�9�Jm����T�q9�ʡ=)�+��s2+�<k�ήc�4�j���W���O2��/�$&��I�wqn��O~�Z:��ɹF�N�D�\JR�LoW1/J[o��ѫ	$60��W�����_H��6=�0z:>`�[���L����D�UY��z��Q����ɫ��뻄�t�C�6K'9DB�o��o��.xS��Q���	����MKf��ϼ8��ۿ����gϞݾ}{gg��'������\_��gfd�������>]�SmؔvW�:�rGՈ���o~���˵SM����"���o�
1"D��b>m�N��̧O��IN�t!�����LN�6R��^������Ȩi4�t�gh!���)G�B]Q�h�z��T3��D.�'�f�J��-.���#Ä�����L�������r��s�>�j��ZJX��2!�}z��*�~_�ƀ��g;���4w]|�kz_��)t�\g�椚@�aJQ�^�<'�T����O�_�z���Y:Y���w�P���a5�m�=�	���n�ƥK�wg�����m-�u����������	Mv��E������_|���ٟ�ٟ��Pea���
'�͚��� ,�JO�:ػ��)m�����//�'aD`Q�A�	o#_������h�o�}a�o�xIM'qӢ%�<�mW'����Ư^�4�y�ts����W��������ӧ��N���!<��+�e;����q�������}�����s�d�f�T�kNMXd��:��|���,�t�-�l,/4�g����4��������p4�k���꾄wի鑧%��yfa�!]M��ш�C�}��;o]���2G�,@�Id;G��h��Ţ���wQ8χ.L�e��%shk���VG�j��yU:bhXQ�j~1��n��S�&s��N�>@A!aNT��~��������ց�Z#B�G�c:�F���w:C���s��2{z�u��\0��,2�(�V�|9��k�|V.�v�ي�Y�I@�N�vT� I@*�f��:	���NO�����;.��"��N��.z���tpI�\Y�H;�w|�7�����*�x������m�rRġ���D}@�*�}��?l��;w�ݸq�d�`�����׼r��G}rC���bBK������h��j�GO���Ew���Φ����Z4f�J��;��1�!�U���$T$}����x�hIq�������5�&7�_@�n�t�:��F�+T�zRU�� �p-}�f���5�$V�c�l���Mhxʊ@#�P�� �Ms:o3^�����$�r��A�WT����ƥ+̌ 4ˌE̟V*{ M�F�z�Q�ԭ�]WB���G���?�^���9�.��xf��T߼�w_�M������6�^)}0�	Sp�� /�n;{��߽#��V���K��2;8������Jz��ƚ0�i����h�]X���,���'y��*�g;/h�m��^��{�y��{��o��.krtP�N��б�Qi1�?2�tZ�8i�uC��0�����LC��;w���h�-�Z���}���~��v���G2�	�f���WVZzajG���ڝ~o���'��
9IeN��Ե�w�<x�dee���yvlo�����ᆍl��K��Qn��8J�$�$<��������������ݵ>����L]\�v�l\u�	��{	����gF:"��a]����Y���V���B��?�k�ܿ�����K���a{���'�Q�s���]�yD3�̘"��H�vo��5w%�KC��,'8��ߴ��&T�ed�thY�ܬ��{@�c!	��~�*Yd�F2^��(���5j2׻t�����p�K��0���r����gHD^�?Su�g\~�J��O=��b�lUn~ƃ2u��鞞�\�bB,*T	�$��u3������QF��ޤ����~�{��ϟ���~f�\Z��$U��`΀d���\Y����������u/H��^����Ϊ�V���a��Ί	��+(�1�'=��b�,�!������:>$���ݣ�HaJ�TV������N�T��t)�����L8^��_:���@���fH݂;|W*?���|^z��]�,��m��k�@bvM�HF��|���6MN�b��
u�5,�՜7GOq������[��B^��$U��!;�+vl��fj)�U-�
���`X Cq�n7�d<�	x�.]�D��d�)�a�"O�~�9�S�w� JՐ���ۢG�Ъ��V�ت"I�� �iB@e��Z2��
��T�o�o��KL7L�����_c�3�J�w�w����;�g��w���X̻��Ҟ��?�]��lq�YV�?Rz�dc6+a⸆C��L�O?�����Ο���
/�|��upt�.;� ]�P������t8�%*�+�s�I<�l)�hm4��:�,d�F$
�a��d�'�VIG6\�u�v��(��Ȭ�d}�処�,�-�7O���m-��_^>�
�68��0�yZZ��k6z�#���&I�D�+ˈ
��w�H�.
��(��t�^�[�X���gE��t��?�V�f[��;�l4��,ы�]��*�+i#G�<8���W����뛟\z��S?�=�|���%!� ���a��%[F�v�eq���@4�.����kaa�������z���tr��76^�|\|��Ooݺe����)hᷦUʴ�;%�1h��P�3�k���+ת؞,�����`A$뵥���P�K�j����6���W���O^����
Ϩ===� ��L~�� �'��]X�.\�a��������8�@flQ�I��J��p�J�
&�n��=��>�}�e��'�|B2�XA�I �4b�0湛�3NA���$ h��M>�-t�Q|�
�馍�&�OY�	Q�؃���3������hJw���3��"�DO4�!sڮƣ]K�)�ȷIKD4[���pnZu���S�L�ԀI�):%����?x��|6J��������Ç{�\u�P���nVe1��>2s�Hn�˩�d��U=�I��������D��
|��qs�\ ���<'+��;ߢ�X3����EF��LZ��k�5��O�C�<)y�n,��Q�M�m��J��A��U�UY*_�9N��Dr�7	����z^L�=*��,�6�r������̘�����o�<w�\�gq��v2��ڈ��sSj�AMG�&3����Qӛt6�Q�6�e��G:�fJ��J>��C?��7�F~m}4��Ɯ�D���[���,�T���,ќ�$=�Na�n�Z�jz�0,2]e���E�K�6�JC?KD�|��<��c��}�8���a�ǺkE���9������tTh���>��q�w���\эЙ�E�w��t*�)f��8o�օ)�`@���G�m{+J-�������αY�N�by��������v���ޕe���P1D�@�<Oۯ'��Y�i�p��t���޹�˴�����9>o�|�%s�6V0z����pn/��E��n-��-�t�3i�tv�[�8�C�Z�<�2�0������ג7���$l��ڤU�P4=I�4�W�QP��`�w�js��d^��w�#��.s�N�0A��K#1i:�M�@6d:;�T�Y����˪�޿�V�p㐮@��Rs��qTu��E_�z�"�۪ꐩx���M2���j�?���$3d���<��VA����Ȼ�!��t%�$�o��Ejl�?z�����Μk��C�֜R}K��� �R̃�>�8~��$Q�%3�<'�����i�u�\����G���bpz̏��~�s����s%�
)�"���b��_~�̍ 2�ק]��!I�´[�z<t���o+1	��/�h ��6�(o\B���T�F�lq2q�2T�A����l�䠛��=�@1�r�#}X�%@O���?�#d2����o�m��F��\�ދTEg-����ӤdrS�<�X��4�H��^�@7����{5������O�F��TM��#-��:s�]��t /��FBg�4r�sNeU�"{
3Ƹt��.����u5���tR(QY���h����{n��f{� �#0c8��k.�⸐�~��X�)�-)�	;M�ˈ.��'d�I��,H��ߠ�����T�*�	����<�H�����h��#�腮g��ʪ=�o=|F�5W5��	V�He�f��X�c9C����b �g/���8|�%~ͨu�Q�I�z�9*����T?F�t���
@���Z�t��9=<�G
2J�Y�(#��vVh'{�,27tg�p �㪴暆��e���*?�.�#��5O��R���*b$$j<I�<+S���p^T:�Ũ��J&z�hZ���A;	���2�ΛS_���NZ\�� 85�SE�5=7圢X�]���a���E�I5���y�af����9�H+u����-�u���8>4�bWw�+k�{�݆��"�c�ኅւ;?'yu�f)r�r\hS<�-�y$�箽^�2���M�P���q�
>��P~�F7��&�LB����2��t���ɽ
����.'�+n�V��Xe�'�>��6��CL>�g�I�ٱ��/ڣ���={���G�b����(�E�u�����$`�Q�a�[�*8xT�!��S�<��	��0�~�G���bBM���KH-���LnG�;�_���JM��WP����={���H�-:��ޣ��~X}��Xq��s&���0����{6D	�~�k�VWU� }�G��"����/4���I`x`�dw�b�v:�Ω�P����Wj�N}���ch�Ѐ��N�q8����H�[F�YrX��s��w+�1�]�L��"Rz��Բ��`�:E�^[[�l�,��vE?KH�n����o�Ω)'�i�WI���k�[��v����Ya����m��A�.�ܓ���$Lt G�B�:=-Ԝ,�zn	��,G{Ғ9CL�bof?1-��Ma�aJ�C��wF�Bu.����X��D,�Ls	�'��Af䃚E1*�P��W���m�E��7���t����7yE2C�x�<=8��J7�Y�5��,��Et���[��=�D��";���4�QXZf�%�4^>s�o��=Fn�Y����q���zv�P¥��2#%[ 3���`x8h�_�����������1l�yX��'-�p�7��J�}����sQ.�[��ԢLb'o��#�;#�!A9�]H���+U �I�S�,&�4�.H��"%|{���,R�ِ[���RK����z��k,XVW���ݬZ>�9�д[z�,�E�l��N�iUӴ;�^Y���}=;j4_�[M�if�x&tj�(춏�m�)/eX����{�{¿�V&S`);0�˩���l��B~qs��JN���~S��i608:m>�)�ћ�՚G�+3U��! "9NP�'|�Q��MH�\��r+)�Se�@<&f����B���Q&G��ӧw��c_������v�v�OtT|N����Tv=����TJ��?������;v�]$i���09cq<K�:iR3����8%�_��#zEG����H��C+A���ޤp�$�(�5��k׮��]1���%R�hW)N�E�h�ru�D��(�!��{�.ǵWSyV0��Rs�ԩSKr`��X��`۪I��ڈ��K��v��xM��j)x\�g!C���6�B=����Ƽ\Hĥ��{���W����R\.�J�W2¿�P�y����+L��  ���&��,�n5	I����(�l��C��rQ���!4'۲=��%�4�_#:�c�Q�y	�{)��P�9Ii[�~�]���EͱL�ayM�v�9U���	�C�s-fi˔$<>T�g�V�UE?���}~�������˗/���?0,���Z���10=]9kH:��Q�G���庭��a�v5 �	�SN������-DXL0�2&TF�b�Q����=C�"2G�GÚV�ⳏS��ԫ!|�OX�e6W�K���4�̺����;�>�3��a)ʖ1���²d�@��p�]�����m���6�	���ד���au�zH`�Y|LR�WdܗP��LrE�j�����7}�#���=�<�B�F�M	�[��8;�H�k�c6��V_����Rk#�4Ԉ\��x4��hܨ�̬�3n�}��Y	4Z�m&��"=<���{��m�m^��jMQ��.H�<�
�ʽ0�VE��I`��U�=�o��B")�z_��t���}u:Z�Oĩ٧9�v�J��~9��ix��e��:vI�Y}�(1��;�f��\d�f�l��"GDYϜ�g_�i���i(ۤͪYV�t8ө]����K1��d8d>Ռ<�d�9�6�m2�$�<�����p/؆�t��;e0(�l=��1�5�]K�Fm��լJ�ڿ��oO�a��������^z�L�/��~�D�zv�Y�M5��0�/�G�g&P��	�_�OR��o�&t��g�#-�,sd�&�g�)�!xtF���ns��ŀx�+�c�@�&EW�;�#S�;P��$��b�cZ�f�Q<�zԜ��ْ�s��+�\��9,�4�GŘ��$�f�@ͦ���fF��T|~(��v >��=���z�>��4Ӣ-�
5���rO=L�|L��2�(3A��&�t��P9 ���Q΀ċ�uD��[���S��{�OEX� 3in��f����s�	X��O`!�la����Om���@Xܱl�u�:�'T���(	�*A�=8�H�=����'!�vg���Fа�����p��� u�i'<�V4ɳ���R��� c[6��n���^���0���rPdC&F��҆Qu?���4�A��"'=�9�;diB�МjZ<�ڗ6V�]��������?�_ʯ}�k$���	2�%��䒞����p�t�����)+�|:ä;���BJ���B֕ʤ����xgg��4P�A������V!�T9�;��ƌ⨧2�)�Ұ�#�LH���
�%E�DNWѐ<BM8�g���Ǐ��Я�E��	8-\�ƪ�(�b(<FM1�+����x&��oz��YjO�8�v�(��p��Ѕ��qܝ1�EN(ם���`5�4l�z��1R;[��c�Vex|���h�4Ys��\�j�L�P͂�B�p����0��S�3�I.b!lZoL�P�ūd�W3?��z3C�L�	N�q������6�����d.�����4���')�b9����38�t������0 �99k&#h�:]��)^5�tƃ����>�����J�e��k�̞�Z�M&yP)�StЯ<��x<�������O�O�h��7�q���lmmѭu���L���`Tgn*?r��r���M�w��{��XM�Ι9Krf�@ߥ@0k���0@�D!���D�y�e��$�7�|s��+7����HF�Q���O!�=��B:�3Ń0sq��^s�?��_Q������h��ItL��.�@i9�q?����� 0�/���Y����Q�g19��$!��i�S��r��.�R�ы�yU�U�����Bg(��,��ko��5\��,�)�heU֌=0��<���J�u������b�aU�S9>�"
���b�݅^!��k���D�vm�J'��A���C������"�����X��<��/�\lu;v�th��Ir���5(cJEo���c��T�۫�ӎ����5��Yi<�=����lӳ_y��^�79\QG#:K-�|�?��.N�)���օ�욮�9�b�a�+ffr��:��s����t�����	��Cuy��3 ��l��Ъׁ���%&m�?.�׌Y@�,��و|8�����	r 2Z&R�d���1�i��(L*.m�p��KK<��Ӆ���f�΢O9���Ј������� 2�do]���ǝc�:�N0�\����X���bk4�ms�ɉ,o�*j�,��=a\����#����B�@�H�=���7�����q",x#�D��3}�a����+7���&/j�������s�U���LlǴ�;�Gr��Ǟ�O1Ih�a'����2gg>G��:8��E
�5`�N���J���^H߼yS^hA��񫯾��OER�:��o�Iwt%	H
������?6;f6�8 
r2c�+�ysHhf���03�,����f!�A����F��Y��6juu�5�d�o�̐T� ���Aܧx�Cn3u�������K,���8g-Ɍ�}����d�(���+�~�-�".��������.�^�	>V��JR��Wo�2�x?��U�ݸ\�G,�v�^1��kxd��&��d��t:m���x<$�NBg1�Ɩ&Ղ��0�wJ)יdӭ���;���J?L�-1��F�um�"��8�w
:�Wy~���b�r@���� ���z���=�肴�~�|��-O8^�<`K�K�Kj��Qa7�L�I��X�B�!�k�[�`b4�گ�|�=Ɵ��oܸAK궺'z�g���	�[��4u�V��[�]^�>��vg���I{��{N_|~���wK~r�ʕ���ե���F����c��wrm���ҏ���,z����ܥ�q��V�gi�ϰ9[.b��œ:�2@pbJ�Kcol�c���'G����j���ʔ��23?;8�PI&�1V4�@��yI��k���6؅"+����]��W;�fgؓ�+�d���p�f]��C:�ܿ��?.|N�����j6m�s�Ԛ����S�|v��@k.<�xK�Z��5#��M?b�+�ZY菊' �s"�N�8k�8�|R�*�+pY�}�;�!������-��S4�����ښ�[�nݼ��������^k5���t� �m�&UK�$��7?���k[�G{���>�������0��/�x�b��(������^����#t
{hsA��%V�W�n��~�hm�:��!}�ߍH/�-_�t�q|f�,~�aѭ1�yA���F��0�MKB�kȓ�~豞N��9�!X1���*jR���|�?�<w�n'��6o}���֋�,��m���4[-Y�p�ԉ[G�~j�lT.�y�[�w��Wv�͌C�
d�HƋK9水���IqT��� ȩw����2�~NC��WL,�X0��2ۛ�u��lR�ȾMg�T6�h��`�F�2@�1�ÙE�v#��Ѯ p�@낪I�td|�<�i�`"�0y���
��Ƞ՘��w �q�YB2�I��S:��՗/�e����:�*z�V�'U�A�*77׏;;;�0��� �S����X�r|;�nU`HV�	�˖7P�2��V��QC�G�0hD���FA�ˣ����a�7n����4�E��l'�IR����)V�\I>�-/��v� ~��i(���ӿS���sզu����N�/��/� c�>=�mml-���T�����f�{V�i��T-�O-��\����N�8��Jed�����������2-�'x<�$�<�h7&3OD��g�+������师휠��+�Ĕ�����m�T�{���t-5�/[mw��sh��lO��mx�ֻK�[�DM�� ����x|gB/Y�g��>�.�<�e��x��μEHW���I
�9ԦJ>��S���w;�OO�
���G���}DC"��D�J���/#���/t�Yw|=��a�;���@�1ILk�Y�Zά���` �E�"�U�oR�d���+<#^��<.���WW�st�M���#'OL��5�$�B����<���E�w�H�ֽ?-ħsnY�ǡ�_aZ��߿o:;����ݳ��K/�DJ���� �����4�&�I���1}�:`:��Pns�D�,Y��v�A�p 挿����SC5J���˱�z���a�׹��ʠ�+�U\�.D=���N�~MP_�$=����M���0\=��	=��$�q�a��W�Ilr����^7?�F	^>۵}9�2|��n]�|��������c1���PO��{Oßk��#���9�2�~i=}��a;��4Y'�q�.!(.r죉}��p�4!Ѱц��j�$�W2�J :E�d����i*���v��J?� ��˟��[j�|�=������������4عC���3i�<�1�E����s�4.Tӓd4�4pT��0�#'�{��e��������x+�0x���N5x~cu
7S�k��A��i�{�d�����0$D6?�^�X�;�Vwz������|�,	:��O�ٽ\X�t�ei�+�Xe.X���ԩ�9�w�;�����l�|�t��f�rX�(N�i�m6��4RN`��ÿ�m����mz������50n"�Px�A�E�����>�Ѷ9eWt�E�Rw�b{cz6��d�T������xD�G���V3jEѕՋY?>�0�jh"떉a8]��a*1:;�o���9�Z5J��U���l0��a=@p�Α%*���3y+�����XS�}����^��)]=���'>t�#��ٸ�����ֱ��8�|�r��=gZ����T/����B���zt��)w��!]����r�xBrF�1��& 2���]�����ޢ+�p�1W/�A���F��������ѯ�s�	
�9&+��D�2k�Mb����W���l!V]p���@�ͱy��5% t;�}��'r9$W�/�� >Hj��W�a=e����ݻw��ʻ����g#�أk\��ݭ�1ߵ^`� %B�Y*q�%�J�2Z[i�" �3شQ�<AF9
�K�YZ�����`�i��EEw�B����JZd�k�z\�<Ӿ���p�W��|��>y2��gֈ~����=�����$ж����1ﳥ-�Zs35?{r���"���6�_�n:�D\k�9�~�}�f�y]���W�s9YT�sk���%�yE�ƮU� ��̭T�Iў����ݻ�#ld��5��Vg/\��
"����Ջv(I���7G��@/d D1-��h�E�F[~dE�|('�����1�������u���h��a�ju/Ȧ7-�dx�5��]�g��� ���`|BrC>>��O�Gdȃ��אM�!�ޞm�F�3"�yY"/C���Q��*̬�͝�l2��DK��]K��
�ވ��Γ���m�jDe�Uh4u=�z�_�N�Փc�I��Κt��7.omm����~��ǃ�i�6�p *aW�� �dp�{r��Gth/�\_�����-���?�����XZW�^%Էe��S���9�S���$=
�	qI��d=�R����4�ۍe:D�E/v�&Y�?X}s��������q������/?�V��zk��+��]m�7��6�/���-u�1a���6Z����?Vn4B���A+n,_p-�q�Ќ��$�9����Be.�_�_�Ys�����t��s��JU�	r3�C*.�����x��H2�j��<y��£ӷ�~{}g�-k�j��ƣA���S�DdiI��P��Sʡ��tQ�o@��I�iU�&��z�
�R�1n!S�ѻP������/�YY�Kv�#5r5�^��;��ˠ�*�hI-�����>664�R��&CR�an*�%X�W�=EE.�G�G��(�>��Ͽ�����i㩙d�ڕ+��D{�fS�憘��K�@;I{kHQ������3Pړ<�}�'?�In[`%�y,��8�0Fa�AZ���y�&zRs������Q�����ӟ���Ѓ�)t��o����{]���� �ӈЂ�cd
�n��<)
3�Ǭ�ߍ�-��[������2�2l�
tIR��Ѷ��[��W���*�"&�+��x�T��ly��ӏ>�����Y��)H���������.G9�M�"R���k�")�~�L_ٸҜ�b\�g@iI���d�H�V;�S�3�T?|�����?��?�V;������@I>�x��*rI�#�-z�$|M��ˊ���ZL�3�J�&s >Ҙ�����$�Yk�I��M�z�M�P*�&Ř�?���'�K��(�����{���7�t�����8H��;h��?��b�˾u�-?�tS������_��D�m�rɖ���+�A��ۭ+��ͯ7�~�[�����O�<�?�_�ݍ���icx6rF�f�9�Q���ZYA��4C����kV^cQ����H4���I�`�Wm�@$?�׏�����Wz���F��qa���V�a!�9�۴W�d�NOˤX�,-��.�b�?;�c�To�B�J���\O�Ur����c�vI�#,��E)/����:v��p�mNz�63l$H�9�E�����D�/��,�Q�[�����-o��w�#]N����S3N���ґ�vh���u�q�<㪕��ܨ��	6s+�W�nE۴���В�䁁U�H����-�ǖ�`m%�
���:֗��D���S�`�}B'�U@�>ז%�.'Ib��-��=��q+�Y!�N5��y�d�N���a�����������=L���k�CPΪ��B���ifm��im�Y�F��������'��.����@n9�����o~��}�{��;w��J�����:���^.]�I^�a٥e������d�!�ja6����Šݕ�= g�_IR�u6����~����1zL�����ǏON�i�k�	��pe:�C����|���ܵTb�/��N�:��Q֊��J-���HO&��S�ԅ�p���'��MUA>�t��::)~��?������,w�j��]n��~��@>)���1�,�����S�\�>yv���IU���R��\�x�/<�9U�L�"W�S��o�����ͯc��=L���8�=�2����_����)"��x��n5u�q�K���7}#�ј�U�PAk)��v�ݟ�=��ގH9���9�6��q��>�샿�+�Zq�T6��$�W�."�����8*N��Zm�p�N���Ĵ:�/^#�Њ���m�<���iٍ�n�K?�^{��w_~o�Y���������/����~��B�d�0X��e1���N���>>C����@����?��|p��	����n8��ݵ�L�?{�Kk���-'qZIw��.�o�m��y�����եNg��1�Ď����խ��%��][�����8M�& �aI���+�UdY��<x�@�D2�!��̈́sZzxx vM�dhH���'S�sa��x:c��lC��Ф3/]��_���B��N�#z��?�pkk��>H�,K��g���_��5�*�� �Qf!Pm����y3E�&�1W���d,�7ވ��'\DWvv�	�m-]����+�\� �W�r�Cg��6�0��k3L_!j_�כt&��u���+W/�C�G�t`x�ڵkdIֶ���"U�����]����F�� ���R*iҖto^z�������"r��S��=A�D�c�&n2��g����~��}3�'M�7�b�n]k���S?;+�R<<> �6��<n�����{:u�86/ƪp}N�:O-sMi���ݻ��O�7g�k�AXY
����y�i�G쨹 ���\�p��?��z���"�AD�]��Y9��Q>ʭ<	�L�CWc�zW�TR4H�Tna���{���������ۗh��J��_���#�t���:���<�Sr�r_NX��З��k�L1G*�h��oS�q��$���J��,��t⊻���+�����o�>8{���{�?��2/"���\7}I�H���#�����tp�3���Pn����A ���Ɵ�ɟ<�sHZ��z��A�j��T�pt:��r��_���K��V����q�o�n���"ou�����M��pN���F��k�d�J�m6|���.��v�"��V
��%�M�&J��(p�����%��8��N���+��Hc�mD!����`�*�iL�q��ptZ�U���Kᐵ)2r@d<��jb'���0X��^H;����\����Mr$l]Ge�¸�l2�Oǿ�\]�@gm��^�/';;;n7��y�*�H�ã��ə��8B�z����g#�HA�\���՜��wkW��[b��T�ѻ8�\��y$d+���(~�T�oa�x�%R����H��p�F9~xt������/�~~��H���/��;�6�x�Z��pWOk�P
��<���9�m��+��$B�t::u�����-)�w^�������H�,�[�c��Ą�]A~����~A��{Yb�'e��DU̴2�\,�#�B��7nܼy<[�2��*�t���Djs<@�Q�����|��_�;ྊ9�Mo�3d�h�mD�˴#����RE�LoR�Q[%�,��t`�g����sF_;�c�3�|��݆~B���=M���)0|��Gc`�5q��Υm��>��~��;��-W��U�����q��HLb�U��F�x��3ۄ)�o2@�#���!L�ޝ3��AW_�gt)�	�{��t� ���3w�ZB��f*��mn���v� ҈
4:��F��^'�++�Gr���
�*"l١P��j-N��KA����N3N&)]�Q_q�����*4sY�����|	��)P�����-f�Y�H����`���p���� ׷��|絮����S�*U�t<X�N�g�?aÏl��7$�'�����M4	f�*M��q<(J��G~�L�r�iO
���8��G��Ѻ�h�v��o/<��S��V+�*�S#l˅�VڍBM
]�����NP�NvR�qK�	:��&5�-�"cw6�����M��-�4*���ӧ���H�ڎznS�����Ӧ��_x�����i�߼��~�ӟvDSOPl�"�}��+1h�'#�X[�`?I�4��b�ǉ%��*+�|M$3���|�^�'u�o#sx���1Y�LV2��8Ά����N`�m�#��.����C��w�ʑ�\����b�p!��:pz�.R�U�8X=�sC`���=��w�}�yNF����h��C�ZJ=_�i�4�c.h[�0�J�n����f� �8��6m���:��8����G3�;��GڎD��N5z90�z��<r"�`�e�;�2� ]����]-t�!��!�cMʏT ��L<�QO"�������hB�uk����Іx!bå�B$�W�)&u;��;�}�V2ӎ�bI=���B�x����;wЋ�!�Y��-1}\��<7�Q"���%�"Ep���x2D�Sg��|����^2>�eJ��	��қ/�4�2�VB����P�����j����\��r繻~N��y���1�X�/c���I6�=U�Ϳ˵i8����[��
U�F�����6���Ս����~�f_|���|l).n_�\'��K4�U9We,�jBi1�di:7�s�Y�㈼@UVb�j�VA��W����c=�$V"�D-9	�	����DY������ӟI�F6�ϊ,�����(��i�z���b�=������IR���{�Z���k��Fz8���;|rX��ZN���׎$`�f�"s��d�`r�e���u�������$dL�h��Y`e(n=%L�ͭ�:&�nў�Dm00O���p<
y�z'���H��8���w||w��
<�;�"�r�:[ĩ�S���ӻ�&���oa·*�<����Ԩ7�$������A>�+{TNߋt�����^[ik��YE�(����I��U*ۥ�!-��xR��su{� ؓ��O��{�k�]�p�J{�@�f�s��?IǇ�X����z�:�a�Z|FmlM3�����ke<C������� ��Y�uљ�g�ξ���8�9�6�"i6�!��v��~�����<(yaMl3;��Y���Y�<M;[1AG�Ռ�ŚMn� c;"\�W�W�p�����:Ӿ�%����'O�&s<4���G,+CSm̅)�3��9c4��|��G=�A|�������+��պ?~Jz�
Ѵ����};6���:��S<�63�
��)@�Y4���t�Y���#�Oz���a��.�e�N��%K��M+5�TVjX�?���y��}ڱN�� �P�7"M&��q�8vv��N��p��-�4�:��yZt��0L�~Nk#�I{2uQ�xqm����D�j08A�:?T���y%�</aꂪb�)�_z��4
 h��69����-����գ!q6I�9��y����YۑA{j������y��y|��o\|�����/��on��@e1?86)RG�� ��B-(�q3ܥ"8��
4L~�r�P�N2k�N��4�'ON��������%�M�Bv}o�)��t������^�s��-J��b�Lϲ�5�Zjv0����P��XI���$TEw9���O��t$����l��a-�@��$з����t`�N�i)��)bO��ʖ��M#ϧO� 	/:B9���8k��W�'\�ON���Pˎ�a���,i����j���<)&��ip���?��ٟ$����/ONzd��r8.R�`�*��ђ�p����[8��(+`��5�<}�{�0lD#;!�c��p��_&�z8>TÖg#��Yd��&;-]�j�������h��N�I��#�!�zU�FN��^�����#�ۋ���H^��S� \oR�]�)c�T�WQO�{���;�X�O���jb�kYSc;�A������ӻ�N���^z��bD����k��ָ�L�~�J�a�Z��*s~��/2��Y/�ЦfP09�i��S�{�R���i�	CuI����(4<��'�L��O%@9ٖx����*1�,g�۔����Ç��ʙ�q`ZHi�'���?�XD�~��1Pu{{����+?��R��������+��O���}�6w�A0�,_���~��h3ų��ȋ�s!����޺�Y6�wH1�>��@���1wn
$Q�;�i�z!Q��9� �b�ߢ_G�G�v��늴>鋭������	��l���͹N����Ҷ��`TU;�h�d7�sd3#����$�<�s�O!g��$ͤS3�K�|G�����O�o)���'�,�&l�����W��V8���dR�hĔ����L�ғ�������&ѓD�qq�����{j����~��/_��7~���%^�C�9FEX�\�F����Qs��Ԙ5Vyd�Kv���%��^=;+�Q6:�W|:d��㺓�}S#(� �}�H�)�ȫn)}�1�b���Q�d�IxiM�2���#o�ڥ��<ȑأ+��a[�!����F%�,	�.nd*�,�[�S����~�����h}����V��0��-y�;ޣ[�z�������R�k�4T�L{MUc,�)9?.i�n�9��[��Rr<�4;^�\��X_}eel��6-~%���u��k.{g�*>��|z|�DV��@&���yL{�zH�IB�����W�-Fqv����vc��K-����;�Ȫ�Q�9�pJ%�$�CO���2@��>�����\D��kX�I<Bx�ן�ǁ��`���W^'�z��&���)�1�s%Z[?K�'c����	^;�	�_<��|�y�uAvN��Я��Ro���I����</D3�V'� �~�`0-�y�S:�g�%�K�}8��� �h�Ţ��������A��SP��WP;��0o�IFj�i�`�6��e�\h��Nx2��Iy22(��jE8:<�t��l0�Ts� �n�RG!l�
kp{g�\'>�r+�}�9�k:�d5I}�z�%��	-c�i�sӗ�G|+~�w.tְ�<XI���Y�"�lSd�g�]d@��8����5훽[S���Ǐ����N��+�X2�y��uV[]���_?KZC+l�z�LO���z���̰�@���l��-e5���G?B�t��
��|� ��x��I=�	��i15�1�N�FN�0��'�T %2�K<S�@�nJ��,cZ�Huo�U�%W�a���+��̡|&#�ͫ��E�F(e�&���ߗ��:Y^�>F�,�^+�̤s1����q��A)�s�f�m��������{�L��:!o�W
m:�v-\S��9��fS,���� ^����a1��rdR�)X'�I����ՙN���%'xysg��Q������l5Ԃp0�U9���ᑲ���E������u�͵�����f��Z}�}x�:��sǾz�Rsu����(�Rh�`��⋇��mǷl ��
R���h�W��Ii�/�d�{���~ק��t��*;����P�ja��0�Y0yrP`'�TV#�A��*ؼ����F�L���TAL+�*�JZ[Y��&e�fEX"��&�m���\�����fx��s��<��f޻��A����jsխ���T�r"Ih������&d�	��Ώ-�UU6���V����Q!9\2n�fb�"5}�����_�\��C�sE�ЙEU�t]`&Cxb1�q�%O��9�!u��E:���[1S�&p�y�#M�֠��� �37��l;f�P푘�JxfE�XA�0Ϡ�*����Y<H^,/���Xnb|L���n
�<9���qnG|wz�SC�q�BO�B��Y�Қ�C:17to+Ԃ0=����L����!�n�	���h=��<SA�=B���Ê
��.0�!@I�A+m���m!�K6ֈ���1@�$E݈ʙ'?G�5A��g��	�e��y����z湧\�͜{���.s��2š$	K��9�����kZ{L�c4�Yt���6�Є��� �
�A��$���|��L ����se�*�f��\EX*��#+�ʬ��#G;^�~�>A�9��[*�d�z�R��P�r9�fVd�R����dťr�N��
��h��~#�)�3�,���B`_�2t
���������u�]7�e�Z�8`����&��~lX�9����g�9��+�a��C�xf�F��$�&��<H'�M(.�-�7�NX���.�!2A�$�%��
jH4Ʊ�Q�I��@O��qe��Lt�:��R�(ؾpe�CyY�p/�B�3u���ioU�z��j9&�BZ��m2!��)��������ak{e�L��1O�
=���l�66O"���*�'�-��B��U&���Y�LA=9>"�d��$�1D�(�ہ�����@���D�^��T?Y!W��H;�B9�\iXݮZ��O�!�*<LM-�}�j6�sN3gQy�����e�c���20Ae�H�U�U�[~8 ^♁���|&[�C?ݾ}����e��ce3��������|/p���ON\� �	?�pe�|�����،7J�����e���hǸ&����k�=,�P�c��Q���%��h��!��G&(N�Kp����m�S�ٶ�y��O>���sZlf�5]Q׮]An�{�Ѫ=B|��1�O���%��*�1�=2�����t�5b���|��
vK�V�vvv��˽��3w{�I]Y229�~�殌Q#�����ӔnĽ�&{uo�\����k��qx"�
y��������5���}��z�����R�X�Ԭ\�1�,J�����F��ys��f�y�?Us�q�N��-�����ȳ�K��:#�}߲̑�U��N�������UJ�Ym�	K�2*<�`73�I>J$�h�����d1 {�*&�#>gҜs6��$��2���3����%Td�|����u��\��d�$��R��?�!w�L�ʕ{6�� �� �z��g��]zr?��ն���:*�P������8l5�m/<Ir�Ѿy����nO��h�b��|�xz�v���.�u0���`�i�pJG�,��<#`D�8�Sd���v�#��M��˦UH��(�O� >�H:D��㨚ؑ�8��Ԍ��1>��X��]�P%[�ir6�>2e�����I���v�n���ho���)s��n>J>�N�V9�t��Rrz���u��8����v���_��u-���V¡��v��{���3ZqƸ@oQ�Zp!�6#:3�q��b�g1�\��(k���Ņ�`Y4���~7����D�;|�/Z	>K�͈&F!xMeX�u����a'pT�0iϦB �r�Nƪ�
,3�VRb��)�����ڐk�9�qy�M�9X�}.9O��,�ڳּa�Fg�B����x��x�Ȼ��2M�_�nzm-��^]�V�>� <�63��aűK�&�c��[#Ca��nt��^��$̲����3��H6r��^slcCL��ޓ8��X�3���ݘfh�t���7]�H?�ty��F�:
��Ә��Q�z����S3/���)�쨦Cx������HpN��o��O�����:�Q�n�
�	�	s�zZ��%_�3f�s5(߸.�g�����ˋ4���[G'�ƅ�K����D�A�U ��3�u4Z3�ݘ>�T�Rf�؄��d�[��&���\R��/�*mr@b���)x�r;�*{8?r��7_9߸�iŌ���x ��K���aՉP\��r�4q� Od�\����j$$m��]��e� v1V���Y<�t:�
�fX%�)(��������H�􆄋[���N3���/���/��@�Z��a��^A� ���j��j�tk�`

�����&� ��:~S��h%\�\����g�ϧz2�%<?�A��
�U,-[5T4~p�1�Z$$1��m�5�x��	NE��q<�K����o(�\u�5��7]�<od�{Ȅ�Қ6e�D�B�$*6�䶏�ǳ�:r�H�%{�(.wʱj'��5��������@=?Y,�;��V�J��հ���S8��s�_�����N���s�%�Mq-^���:~d.��ͤ껪�H����s�lu[]e/���Wn�E�����i&bB�K�G�i�9���V/����6z1�u
��+s����[�25��u��aL�j2ˠ�2S/��s��7bH���~j�m4[6����c�H� >͇�W^�sonnl��0�$�#�5X���oS�T$���Yj��`k�l3��,�����{r��0�ڲ��������j���W�_��|sQ��7����swΕ�0�N=��*sDj��p�)Q���-&U���Z�'�¬���0���</S��P����D���Ϧ��į{:��L�F/L4<��uAܑ���7��f����EU� Gd��}��_H2*ݸC�����構�Y�)�LT!��d08�� �e��
\S�TA��G�({�w��|��V��Te"�RC���m�@��2��_#���:<��̭Զ�1Wէ!����*f������q�{�C#����q�hk��,�^�oNd[�c��m~l5�r)/� 9Dm��3dv�:<]��T�+y��6J�硱��"��8ak�-��kф|w�)<�	�a�}�:�������FI��?� ��Y@���eY_>3uz����$M��Q.���=�n����R����YN�����Q��S�X͂�;�TJFe/��p[�e�aM2u�4���$`�����hS �W���������y(��:��`��{���쿘E�ė�������Xe/ͯ��8�sz�l�?A��,�ϼ���~Bf�@�
E��X��5�`��w�hr+Q��"��F-@/�����έ�W��s�o��f*u׫�V�0�P��Y���tM�y�Լ8��F����|vM΅-��Pmfk�|��k�b���ʬqKԕ�6]w��V��[����!�m^>S��謪�2l����d_8�Vg�k��Y���r�)�3��/�����2E?�r��+�rE��{��ۚ�o�ǹ�N�F7%2�a|��G�C�Ӝ�^�z\Ue��UY�;Pǂ��)+���Um�`f{�x.��~�Fm�s1P����ñ��V24t�V	��S�$���8��g,4E�����R3~�&]_�����Ia0��m��o�����r�u�k�<������zϒ�72���r�I���s���:��^E݁��U�Gh��X���|	���.�ʾ���Ts.(Q�y,�X����	6���Ns,Ă0>��j����ԑ�s���Q^<�s��|�r�3��x�\a���ṋיi��Q��1���������J�*6͒��-���.�f\A�7D�ไ��s Y����g��⪣��r<��,t�.��Y����f%���`F.�H�2:�������|���,̓t��
�,cm����\�>c&Vk䛑I=9�t�ޫ�����3����ӭeôY�si��^�y"iR�w���Y]��~ϯd�s�+�"~T�9��Ѣ��O��WT�e�(Oʂ�+8���j��S�@`澐܋!t���5H2��?��L�>;F�*�A"�Pw��u)��mÙ�O�%Њ�g�(��X�/,L5v�`�v-����T�HAǢi�C�� �*"��^U�q�n��}׭L�!���� �ED�7�b5s��L�q�B�k�,�,p,�f�����΁s\R�U3z���8����Aŕ�Y'S�	?�����A��l����B�Ԥ@�@��	0�@�<0��*d+$e�2o�ፘp�d���<�M�UU�bG�	o�\lϜ0Q8'�A��_b=n��M-����찱d.D�S��^|���9B�4�g�=�����^��`�9[u4�rc�l~��U���/��~����Pp�`JmxL��(*Ӕ��t^$#g�����@��hs���^�m�U��O��>�Ĺ%
3�����/����4��E�(��a��4�q7�$f�D���\��za���?�s��Z�qG9���'�s��В�"1�K�kW�]��")\�Z��x:3�=-�γ���b�os���$c3E��j5��9=@8Įf���X�֕���(��T�*�$�H�:7V3a��;5��r��Eb� �j6��lK����!��eOV��6�	P-Ǩ����g�Y�]�D����I�7�-�ue��	�����.�_�E�%�V&x��B3�^Ꮯ{�F���n;�R�{�(7�~��~�;EB��2[	�q����^�SΚE���F�U�R���"`�!���.{Z��66��x%�(7Z�mfq�p,�YB�Uy,��Ԣ� c8!S<s(e�¤f����X���������]���"c>o9G���3�~�b&3뵨�24\K�'''�a�i/Yd�b�<��C^)����|>9F��FX��GY� nD	aFx�
G��2��K��>I�(�[�U���.ϊz�]���I;h	�քN�-p"2��%cX�ӜN����Ɠ,4m��I�����]DA�|��C�t����r!�\��ՋW��J�\��s������[�6��C!�����I����mլ-ϕ�w�q��ȷ@N18���k��!ru�
��!w<h��7+��@����!<���/0�*��]C/	v�˴�o�ceZ
f$x��U����X���)Gm�g��l.�i����DpY�'G7�#'6�9k��ܩ��e���ʘ�!K��ȍ���W
�b,gꍍ|��Ν��ؠ�f&1�a�VC�Y�9M�=��_L`��a��MLGi�g��_�\�Y�yS6m�3��g�.�eq7��FĭL5�ȳQ��![eg�8c��������J�G���Qa��fS�d�6 �l�[T$��J7%�Ғ��]��5�!���Kg�D� �=��́�`,a��(��e�.p=�«�ȋ����O��5E�XZJ�ղ�{g�tU�h�bq����>��t�r;GC=s�L<�xr���{��z3���P1�9fW,~,�<���^K%V�N�Q:"���D�,m�@R�r��U�_�WH��<uIߺ�|+��������Ԃ`�Ռ$=�K�����u����\"��9�[��*�U�cM%r���+�����CsM��V�"-S������iX��F�j��[�S5�m�"X��]DM�49&���)㫒��D�W�*�NМ�2}�����bz�D>���M�A���S;�"��� �f�[��=ZU8
�/� Y�Y�hs���(ГNh3�9<��N��g�����+|��V�PFŁ$㌓�<88�=~����#9�<A�N�E��	��y8ӧS�C�|XD���{����o�㧏QbA�y1�o�P�Z�%u��c>Ƌ���Q��z���")�YOq�r0Q�]����,T�u�|(K�~.��]�]�J.g+p�l0��Msځ^��wa�C���`I|I_�J�8�"�L�v Z����+8_�m�5�5�o|����!����+T��L�`n9�� W���H�50��g�BD���ȷ����մWqa��"�_�w��:��\�k$�d:#�O�T��Q�.f|0Z]��5���d����#�r�{v�8�z> ���a������f߶vV�n.�?xhu��f=k�	p�l*����$��t�2$�C�v�쟀~Ws]���$�Y��Z�8qK<���ss.%�] ��Z)���\�nx�I���}|2��W��c��&+��@]=f�����U�#�N��i8;m�=�x`�O���>'~�A�3�����Ie~rU� ���+zS��TI=�U�� Ⱦ	/s����t5�c��?����
 �G��0�4�Wž9W���l�rL˞��s�]`W0H�{���r�>���	3B�,#�b��h���l�
�Xrc.bn�_�s8O���U�C�f�BeՆl��ܨ�s�'��Ǝ�i%߻�f�����RF�G�� G��'Fm�Br0~C 1\R���b;���Ex��g&A��Ѩg��g����s����y�����4?ǈa����!+K@���>o|��>���R�*Ű^�3m��s^��4{����`)7�[�&#������|��L�"���H�m��'�˘�9"izF����w�kQ��q�ӧMA�^������Z˘TiB�f|Ͻp�j�;�h81��aTuX���8T0����@�&xK�6���;��F�Ob���$4#Ί�n��˘{S�����C��0������B�� JSa��&��U|6
� 9�&�v8�窱����H�|G��^u���c��g��5 #90  [�IDAT��^P�$fqǺ��3���������wX�[n)��P;!OEj� �u�(ϑ�M84�Bo�ՄV��^O]Ds�jWU\R�Vy+T�5	�lU����XOdq&Ӂ�N�|�P}���j������D� �&�0�N�B�:Isk:�r؆�G�Tw�<��b�f4�3~e�i%�%7Qz�4e���1-��*s�8�
�z�hFR����m+#�$�AL�v�C�J�Я+�ܹ�p�a�M�����uA��-qĭ'P&5�O�r�U�&#�S�i�=����@�CK��C�q�k�k�����b�锑�CY�8�C�W���N�y���2���#3���^�h7��s�S�CH��!n�
<��窾RC��-����=�:-I���N��'2�cq8�i5s=	�V�����$fe��~p�+ �W�f~�b�_V����όN��C�0
���T����WS��D�r��0��mb �BM�V9+�2*�L��p������F	���Y�{+��p��Mxi:MjuNW���ј ��ڨ��3�-����@�.��U���l�f6t��3�����bޛ����+ΞInc��%*�m�
h�}�G���L8��Jkv��n֠%fyJӠiɚɄ��Xl��d�Gj6������
�����d}N�'�2��@��l�$n�ʡ�φ�2F2wc#�8��[`U�-��4t%���`�j�#�$G��&�?d8f�����y���rͯ`�Yt<B�nV�#�S�F!1yf~���/�AqQ`T0Ƞ�y����	�)�˳��*!%_:�+��l��陸I��ښ�>>;8 �M����v�'GG�h,��ȳ��������oD�wSxqN�N�̺��eGa����U �ҩ�`=�$#Ai�EC��7�O��x<�lO�)I<]g8�,'�,����ݴ�O&q�����,E�"��I(S�u�d�7�V��Ft S=�j�� �)��67��n	��~��ɸ������D�4Z����⚓h��omV.!V��7�L�I�r���Z����ɸ��t�;��1�H��~�	����43<��O�6��\�P����Fg#qvww��\�"᷏��H 0��p���kW�*������-0O*��j�<��m�l{9��8٬�o�S��V�����ӳ'ǘ��O�>퀹*�\_���t��.����b�̏|��rME�F�D!<e�qZxl).�(��Ճ�p<n��̬T����á=l�E����eQ)�9�Kf���dK��ͅ�Џ3|����0�.yQ'���.1���j�D�X����s@/f��O�y3"���������"��т�i����$j�H��[^[���s�M��0G�y���>�rs�y�6�/�g=�����ߧ�D�TZQ��w0�!��G�#��y�?�sp�N;���T5�� ��Lǅ<<<�{0�n@��PI]���d=�?�v5+��˪8���Rĉ�/(B˥��t��T���Y�g�>�+L-������Ng��Z���\�
Ҙ2P��s�ƘMP����v����>yD7��]yi��&1s�Y�������˛�>�4�����Fqİ����s����M<D����
�m��4�����t���e��r�L�a�a��%K��O�3��I�ژ�ްL�y��	� �\Y�G甮?"rt�9�
�!f���b�ܓK��+��@7����5�=�0����}A_���k:t��r�h�'�������������*vB�+�T�Fۻlw�q�-�V�1������͛7�x����������b�r�	?��̪����+�ь�"���
�3��������X�9f�NB�ﾎi�>�p��<������o���i�Xg��\�=�;n	Tg�.�.WYYIv�S���/a��ڊ�`p朊����o���;וּ0� ���?�u���������U��qDg�Nۊ|��R��e;/#Wmɠk7:g���{"������!�ڡ+����O?��B�Q���i:����n�5&�Vi;�HO� ؞��vҺӤ����]��^rr��rl]�p�k7�|�ך��H�=z���~u|v��{������������Z��}r��ze��V�h)X��{����p�\t������o��Z�ܠ�~��ݏ>����/������=y���~�L������-�g+b"�a*-a7R�U�7�g���Y	��Ooe�ͼֻ݊S B�c_�<��$I�ba!~b^zƩ7���l��\��?��e�I$��E��ҥK��{���Loqܺ�Ӛq\`��-����TL���/��6�>x�S�����>���Ï�^O��n�qR��u���������!��z�淿��׮�^�^M�1��7��������x��x�9�Ħ#0�@�C�����#/����\~yiuU�N�
��������o��o~����N�8Y���9��1x��"���ܧ�_|q���;��ޟ�ٟ��}['��ׯe��o~����t��?�1t�0�jZLX0��"w8�N$�t��)�������?��? �򥫤~ ���c���7����w�`��	ȴ����ڛ����5���x3:���������?��?��l�`M���������_���|���,��ӝ�Հw��o�P-Ԣ�O2��9< �	�r 6$:?��
�F>��-�5a4�A�F6�������9��4R���|�:BN*�l?'G��t1�B��Q<Z�7֮�����78x�Op�ge����v�ʳ&%��@8]���~��쟍���k�������]�C*�F,�.tW�+�f�����-�1ɸts9,��J��?y%�������;�.Ek'G'ӣ��������J֜��K�#����Ո~���j�����>y���,Y^Z[H���<f �:T�s�e����G�Q1H���������W�^-�5�L�<�����%�u'vo���W{���	B@��HIS��2�,+�A��/����
����X3���4�H��I� ��޻���z[�y}~�d�˪.hF����WY�2o�{��l�3^�x}�.^����|��?��?�u�e���Y���cf�*y���r\O�x��Y͝?�p5����ڿ�M��`��&_���}��Wo�o��n��_�ܢ�d�:��D��+��me*-9��,��!����O��+������ɤ��������3��ӗ?���������w�%O���n��z�?<Ƹ�2��dT��N1�zN�ؙ=|��/^z��菾����������fup�������_���O�ݏ���GN�pQ�ܠ�Y��ɕ���J�Y�)�5��s<O��$�:�ɛ>��xcXl����g<�S��p�Q#���7�4cjg���j�����Z���W4��g�i.��x��òR��ވ��2�h�a�9\*�I����sX�'hC�����x��B֤�r4���&KCNa~�K_"���O���9���t�eճW�O�U�>|����7������햾ߏ���B���d�������Ox�Ͼ��F4��񼔋"��J��c&u��G������{��{W�\Q��������2X�P,�}��;�C>��c�7
��8��ˌM��IP���B-�w��k���k��V�Q�w)��v�qJ��ow:_�����?���t�L��mI?Q�d]��!���꯿�կ~�HL��O�]�%�6+˰�W����к�~�j��H&י����;�^����.�[��[����
0%�q-.x�4q�+��樂K�}���bAr�/&E��X�
�ZufJ������������q5�pys�,J���A�E�-��7���& $�� |W��|�w��	|G�ڦ�k�s��+�=�<��(�G���\a�{*9�/�K���V�����?��������)�n"�0f�և�����]'JS�&�}��~����c�}p%썫�]g�� W�J{=,�m{�囟_�_(t���#����������#7?�ٛ���֭[=��I��b*:3�o����@9���٪��ڗ��/;T��b�>���J� ������/~�λ�ޤ�F��u:%Ay+C�c�,w�H�p�[�_��B��՛_���u�8
�?�A�}E�PV�)Z�x>�ؼ��_�o~��/��{0)�W��K� s	���k�II�:�G��Ǘ��ڗ�2���-�	�1'bB��HJ�-G7�������l� d��d�����r��`�c��Uُ�(����tv�{���W>�R���H�<~Cs�X��9d}r�������ɣw���}�Ԛ�a���fZ8N�t��,ԂF8���&�rJ�óӍ~�:JW����%�<��ܰ�k���l�
4�&�z#e�Z&e�� ̫��/S0Б���S�' �mL�y��X�x���ECDF%T�ӏ~JߵⰗ_~�H�[�Ya"�խSw�7�|>?�ϐ�"�� O�Zd����?!�@g�ƆD������ @�S+���Gj���{#�ss��L�W����&�������+��"�Tu���m?��!��	:�юC�%�H��Qs��I.�T�rct:<~LǓb�6�'���H"�c\��7��ss����ׯ��Ge9g=g7���ı〞�K�탃��|�+�k&�E.���Rپ�4����/|�����%-�8ѓ'O�s�3���#�,�}�@ȍ!�o������} &K��R�ޯ�����~DIf:{��h��\gY�ϐ�A�;�''0���-Qis����xT }	�x}�%Y�eHA� m��*�*���\�A��95�5N�Ý��J'��k�����O~�s��}~�L�v��O���/m^{�����vB���ҕ�S��u:o���<	|�;6ݎ�����wh�Q=�z:TաӉ�zh�̢���v�����N�H]X�a�f�C[K'�X{�Az�w�F!�4_�B0�"��|I�����D��A�2�pe�3v�#x�Ɂ[L,��c��>-�"ټxy���h��9�2��]��v���GG?H
s�@V6tz�^y�wC7��7���Mf�go�ɋ��y�LI����Z'V��vn�xu�#f�(Wg(���b�Y�L�eiut�o�(mf��:$|���G��,�O��x��S$��"�D�ZU1{�����t�<p�/����߾}�7.��Yo��Y9w�������J�w���������n�k+PzS��0�9I�mi��I���}��Wל���x���,&zA����25�ż�rNr�ı�-sΧ̱H�����o��'!T,l�jF�%���]�k�fs}��<��k�LݧcK�����f��z<�����O�@L���m�sӝ$��"�!`(Ia�o���p?H-���e��P:tl�\��gBM(O�>ım�}�"��j�T[/�O�>�v�n�U9�8%��l�3%��hn14��}�NWVV[��g�U#_GJ��:D�2H㩋GQ�Ʉ����	d��p��ʤ>��p�F�n�?s_]TZ��p||,���U���v0��ۂHÑK���D�V&/��!3�l@�p x5[Ij����A��p�H��ȟ� �ٵ�Z���.�$���Q/:9'�݄�I|]:�������V� ���Q�%�8�$��M�)x��;ZbJ�L*,��I(��{0�CB�G�<A�U�kWCI�F<�~�0H��5{�o1s���%�Rg����<��.PE�c��Xe�F�,�dq�G�҇����� 0>)��#�iN�<�`��5����0�кx���g��EL~[�R����k�<$J��/���̥���M����Y*[;��F(\/���Aw0������xs��(���\&1U���\� Pƹ�S�K��i�
X�ic�
�����q����ݚO��`lS�<��}�I< �D��tz|�	:��e��;9�z��6 �<2U��|�~��_���G�̋����CJ��d��<#�g�x� ^��(���*7�外���$'�0�㦪�ᥥ5=8�#��X��"��ia{v�0��v���݃h��Y������T<��³ߌ]�.�m��"?N��S�h����Lim�s#6_L�q�Q<ɬ"��<��N&+�������-0Igā�{qV{z4�k�ĵS�� wn�fd}͑&ج����)����ZAn�'A_^]�@>������,\@BPA�F,�Њ�l���m�/��K�L��\���Ç	J���O�ˉhs�m.{4<��z���A*�1��V��Z����y]Sf:�-{{{/Ўwm�8�>��Fŵ���c:S�{��}:�T���,�
�svM�z�9=*�x2P�!��s/�8gK�EjT��7 f,�*u �MIu�E�3�'��en�C~=��s.��7a�I �L��;~�%d��qX���P�>�9��m���l6}��1��Λd�ɘ{����-��a�������6OA"����*��N���������#���,�\^H7;l������!���'	��(ąy��?���4����چp^�K�Z���#7��fb����jꦺϜ#���ps�Z�Z�խ���G��>}>�f�ePY);J��=����_D�������0}<�z-0�ѭ�+N����'��,���������Di�v�&��URr �8 a��ރ�=z����(M�V,��VG�^��U�v9���<�G=BS?z��^{9;�}CL@�:	���X��l� 
���~��݉�"8*�����"ZSHˢ��$Xg����y�v�7��z�W_%-�����[�R��<K�ꗹ1>���ΝE�ݷ竫��rnf�~������бƝ�?���d���go�y����Q��r���8
lԉ��+:N���G�n���O픀�2<�5���ѭ�0Y����n���ۻ��p�tm�(N=���������H�&'?�O'���޷��O�����s�T�k�I���$�ׯ^������_��_�'H�L�%ޠ���TRJ�M!�E7�?~�9-�ɬ́Y�8�i͌���Fd^�;&��H���bFa�����3�ox���إ��8G6 (�s���T�Աd��k��
fd!���Ź<�pds�C�Z9�̎��!AI	����=�W��2"��p@O�������	�o��W� ��Zq4@�J:=hⓃ���@��`��� �z����2�=��ŋo���[o���_��K��]�@����(�^���|�����!w�f��3�Q�~���]�G7�ŋ�|�ͷ��^{����������I!�2N?�;ߡ���C`"Ym�2�)�'b�*}ō7p�ޢ�~��5�*Y5���(�v=����n��?x��	]-=Z��|93�j��3�~�w�ܡ�]��︌c15X�G6�_��|���*8�s��Fπ��Pu�z�/�o�F��IC�������/�;���Cx8>�߾���Ƒ����[d��|A�icQA?o[���1
��M���Z

K��z4�M���*M�j�{�1a��MI�%Ā��F#^Jv�����WYI;ͪ3 0:����r�,��5�-zNo���
�M��J�z�f3�pƝ������S]�yp���/������vn޼����^+���N=�w���������ѩ��� 0B�@��cr3\���Zgk�7'�f������|��˂����Z0��s��'�ÿ�۟������:fkPl��~�ya��� )��+z�'�����Kϫ�����?��������\�\���s�V��0�{��������/&!�|���$("��(� ��c{2?za{�~z����;���;��ο���?���	�x�tr�j?H���I��Ϳ��O_��{qx\�Ε�Q���<E_Mf{��Ӄ)#��k�$�u�b�3�����o�d�'��K���u]�%�㓡�H��#������o���{�.6���H_��qn��0$5f}���DG�zk�^����{�o�{����+�M���YBeJ>�$�4��{��w��?��̆���^\�	���۵�?zqV~��ͻ�r�:�͹9X����K��18��p���M������,�S�keY�(C����ƽ�y�|9<7��đ9�8������;���9,8��r�^�THߐ���ܤ�_y啧���?��?��׿��+��F�N��;ۍ;�n���?��ݑKB� ]���\0q�Ŕ�.�)��~���� -���[��_#ʽ�`C%�z�����}�����	k]F�4`Ni){��ٙ{$}���������7�7���>�p0�%-�5�o��.i�'O%�MwG]y����b�h����p`��n�����m/�׾���=o,� m���ݾw�ց�G�D��	.G^i�U��n\���_۾��O���?�������#����4�-@fٚ�4�����������.���by��N��&{�F��
ɍ�\�p�������:�?��|y����Փbno|��_��_v�puJ���+��u�c�$J�l?P�%=M�����f�V�����Rڒ���Y$��t��/t��d1��~D��N�;ߟ�Us$`-�Id�(�-�/o�F�t-�t~D���Ϗ�geV���ҳ�=Ydq���G���o�������ML�?|��1At��~�L��,�A@?O���万��f�!��Uױ�i<+��5V�S_~����w�}�w���Fryak�D�������vH2�/���d8�YQX.Lrb�e��] �98ʓ�Ph��d��m������7>|���/�}X��~��n߾����ɟ[��˫q��Y��IMN@^3�!k��Z��#�c����+��	!����w���|�μ�=x�`��$Io|�jz�|ڙO���6��'��b�(�sP~�pKq�S��.������]��%r��������_�ʿ$9�X��x��!�҇ￃ�������FN4�	�G�&���)�UZ��t�ŝ�x��{ǿ�`��������_��sϿ|���Q�G���i������O:���Z��z�K�_�̳�v�	\���Yjl�C�AI��|7nU�2mF�ɑ%Ԓ�PU<�c��aH�w��������K_�r�d(?��C�|�#���JO��s/�/�� /����޽{��j�tr[6�lVtq�>�`a_��DM��?��Z��ˁ�\�k��K�D &�Xx|p�=2���F����z!��+kd�y@
�{���O�X�[�UP~����&Y\�@�k�WB�����0G�?�և���{���k�*v�C��������l���Ι���bb/�{�>W�A{I�L����%4���?�p����׮�
��<��~���W*�tjnC�&N�e6����퐣��.X�=��i池3��,���!/{r��Ç���oѵ}��F֠�s1iYȦE�E��\CY6�A��9hUc\�W���^��gɚ�<>"o�����c����2'��n�d8]��1ڎ9MnT�m�4�� �/}�U��7�d,������n� Ў�.���oD)��	���+48P]蠕t�����G8cş����9�
��\:[𐐾��ý'{��F��7@�cr&0TsV��^��{���A�͇���<ÉT�1?N��9q�9C��:jѷ� ��ihRn9٤�V�Py��~����~b�;8��w�>��B穔fat���q��꿸��)��VP�5[�.}��u_n�8F��wn��B[�+��0�<z���N��s��^#�h�	��\���D/R;=ҠmMY�Yt�0�c�A���v�(�Ԍ6�k���1��<�-�O�|b-��]̄)/��ޣ��^2@sA�"o��P�6���
ŹS�]5�����o�_Z!���9r�`�����(~RN��Y�k���mwE�cZg4Jb��c�T*����w���h�a:{���`�z�t��y��N��W���v'���޴�������:�O�b��N��X���-T�:A�e�ә�v9�+�i(�x���j���
�������˘I��J�OtՀ�)�]���f�k�n��/#�Nn0(�`׮9�uM$�
��kk�E�CV���˨	.
�Fd�}e*�lGR �s\�Y&�Ȓ�����BB�\�G�l��{��k��L|�s���=�ۃnf����Dq�Z����<��j���[Ω�n�	j������s�=�6�IW�J��i��=�GZ���\��U@��&���eD�)�2�蚯��_~y�3!I���[�;!*|��e �D6̓cc�%�G�T�G�9=�ħ\E��]?w�2�����}�6,�����6F���`E���z]��"�d�eGH�)�ћ��ܾv��Iq����f��%{l�ҙ�d���F�SQ�W��|7~TSM��Iڡ�G�P��������qп���B�C<�53}�|��'�7q��bH8��P X�lvr���>V���;��eP����!�&7`�*�Sa�Ճޭ�;[����K��������n�"Ɇ�p�)�.2���f
�X*׮��U']����D�ʅ��3d݋Q�#����F[#��f?�p1qE�ݛ����=yiXg`!�޵��.�-�A>��NѮ}�\�a�ȎNz�=���$��y]��8#�-x�_2���PK��O\a|���M���n^��i/����V���A��\XY��E�b#���q��:z�H K:�=.�PЎLa��Ǆ�X���c���8۟�Q�}i����.}9��؉&O�'�)��v�7cL�iT�p;L�S�W��q>�V���q���B ��]��+%����Gsr'6*2|�8W�0MTo�P؛)M���M�B��0�1�e�sKXx�����|�58�
�t��mGV��;��O�4����*��3[��ϴ�,�j'#)m��#�E[�B�k���cϲH�<�"�R�H�|ě����e��$e��8S��D��ൽ�$�mt��6}K�C���%��Zx��΁9[䈜D6��;ݎt�F,�����(�ǻ�YDxRX*�@��t�����<�L�s)�o�������jj#4,P`>�}M���I��̧O��ƵX'9���2�V�Ć�h��ˮ���g�Lo�"�����١O�A�����c4	��ВT+"�D�T�%��vŉ����0OUX�=�ϹFͣ��'^`?8]$�L���ı2�]��V��U�+��U&� �fWs���a}��HV+]�pi�a�/�㐇B��@%P �k��͑�t��ֹG��\8�vT��&�,��$r*�c��0��ॗ_��K�o�3Hj���e���1K�q$'e�X���K̻@V����N;�F���h���W�0q����Z��P�WΑF!i�g�|���D�	�tՅ�x�.��=���5쏡�K��H�%	�r��x��!�8%g�#<��&����b5���}%$���IT�L����lh���Dl�f���ǋ5�d�@�}���(���e62et�I	҅!�2z9���.S�s@�(���@�璂��e̽Ov(���c|�7�˩�4r*���@mB1��,�;N�ƞF�Ic�Z�?}8e��^��![G*�O�<�mY��#��do��dZ���Z��Y3;�*�.�]�-�[�W�]Qr4�}���t�K>�bծ8�(15�j#}��&�xRK�J* ��K��A�o�QJι(&�2�b�`�u�8��d�%��L҇t{��	���J&@ɖ���t��<���]�h�cdœ����\���'��9���	|	�5VUȣ���#�nE��2_>��|,�9�.HH��
}�`�%��>B�pǐ�seC�p1���B��`��c� �B3�)%~�슅Xf(pq��\���3'<g�f�����Ȅ�	�F+�S3��|R-@���cs��"c�S��������(=F���/+�<�|�n��� 5H�>I�l���nyZ9��Yd�<IՔW�ll�3�i��򛟭�A�S#R����%�Ѳ��P��cE�`�ʜ���G�6U����M&�[)��=x��U�9��4+�Y��7���Ǽ�����h�io\V7�=��wQ����Jh�[���t��F	���G��+՘.`ً<%-�@�ڵ�4A
�[ =.=�c#��"�5t���R )-��9o�^̥B�T�W�),r*e]���Z�N���.��pK��
p�̸�"�XI (�����,&o���-�=��)�ztS�_�ZCY��������y�,+�Q	o�ǌ�)�K���R([
n��m�����R=�$=��9��7�>YL�3���gdK�͂z��}˪Q|2���Z4���n��7d�X���x�JcF/� "�;�`>��$OI�$e\���5s��
)'a��c_����m��d+� PVᐶ���l�e�|{����F�><�w���[t�|"kΐ�0���A�������5����T���=Z��,H�>�k���"3�F��">�9�S�8���J4�R� �^��[�@u闣�%h���Ak������C+R�$�+
� 3��6q�%���y+� �q6��������7�����z�.��� c��������G�LW�˶|c��1Cn����΍��"�}�m���C����\�W�4o�;�Lu�R�ɖ>J�p��&�v��$������m^�r%��{��=X�B��%O��8�m�j<�������3�ڸ� }�e���Ã�!i�ǁ��rŢ�$r��5u����'�"~����R��'�7�U�b*AγG�8�42�l9���J����Y.�+�֬��� ��Ah��K�v$�������E��n?8<�͎��k'<��+���oO�k�H�D�ti5�j�τ����Xy��''�w&�S^����,!�����3Wx��7o�zd�\�o�8���p]?\L���J�9l}V�	+��y���.��j<銍���� �Ƭ�	AZ?�t��̎����~�A�� ���,�_�\ظY���R�hK�\ ��'ő䔬��f�x�?�{�G
q0�8����}�=�7g-k�n�u�U�2 �$י�|�O�6�;�L9�����~xe��w���ɮ�����;*x�-�ty|ʳ7rBHc-���CF*[-;~1�Y���E�"�SX�ϹG.�˿�_I�Fɬ|���V�)��/���z�*ŵ����1�[�#yYX�B��Y�:2|�)l��lbQ��"$LD_ΙS��<4e���a;(S��2R����n��S���?E�"%	�#Z*�����1U�7��9H]4:Bl ���Rs�8���Y�5wrm�	���e�R{���*-��L�l}^I�G��UG�Y�{��Y�I˾�FAl��$�-���հq�h�R���H�h�ga�~]�b<�������H�j���:W����J�>#ꦮ"�B���V��ƻ�9$��$eE>�3+j3�M^��-1^��2���Iω�V6Ou�WPd7�� �t`�v������x2����-;�k$M"��pKU���'Q[��f��w���3�{�'̉�s�ũg����cjVk6��G:0�p�W����F�����7��C`�pQHƌ�>���c���V��0)�;�ق���U����hL����|�E����v��[���|2����d�Ȅ��.����E�t��s}�'�'iEڬj��_H�Dn:r���n~�.2̄�J/J3��9�8/fehF����8M���������e3\�NQ��5UM�u[\u=�{�XT�'����R�e�TZ��UFb䭒�Z��f�if��dW�����AS�����r��Y�H�U%��\��E[+x�O�F������ũV�% 7��t�XuC
8�;��o�j�v5s�hl��gZ�z&�i��T��K�����K:�-Q6�'<p�tgI����VVVn�t��Ar<40����a����)as����÷Z��|tr�2	��e=�P�R@�3}co?Q��&��*N �����h:�q9]]4�� �e�F��KQ�Xݪ�zY�'���ߟ8A�
��9������C���jinS��ʂ�hI�Z9& �n�N���dvj�@	o������;���ʾ����e��ө�=��%)"93hg!�e,� A�������e���6��b�s��<�0/���+�bf�LГk�%��z�T���~�\W��X�����I�UN^V�r�fr����s0��B@�9�8y�'��"�	�L�s;���^\�c.-PApQ��{�&��F>ؙ��\�鸉�6bDV��D�`k���1�K�]��"�c�	��uKt��)�H����i;�f�Y���&w���mB߲�ۿz�ʵ�^2�q�z�9gKa~Ց@���c��$}9����͜o�oZ:��Ŋ3D�N<�Ş����?�$ק�74G�=E˕l�����ʴ����
�z �������g���� enlm����Ы��g�{�Ad�1�!.����(�s���K������P]q��-��Mj!��I�!����n�yUZY"'��EkJQd{�*N�j�<�\]���b�M�D�s��锼�A>D���l�Y:�k>��i�/r������[j%Qf��ʜ�	�$�
J�U��@g9�#4�"m��%��1G�����{
��K��x�h4�
�����zt�-���Xe�8I��2�)��z	^h�����olAu���+��\���*^P�Z�^�]���I�"�4y3ptI���H|a����WV_�u���[���qamks�~b�&V������#�v�@n�[Գ-G�4�c7��,۶�q$�̭ T�cn��t�=T�ڜWJD���F,��m	��ȠDc�e
�e;^r�l�qT�Y'L�E��49�|Bǘ3�(�a$HB���	��UI���4���>>H�z>>�\E��n�}s��d����6�H��������b��.d�q�,��:��C�k�AH^{B��}nΡ�Ԯ���t�ό|�[��<�Z$=���f����Av��a������i��2��Y_��[�E;��-s�$B�o[�r��{)uZ�KD�NB!B�������Vn�MS��Dpy�w�3�ƴP�j��j�X�Uc;�<O<!nG���t��qI������G'''��ufNB?�J��t+q}E��M��$�R���pJ,��9��J�3�7���>6ܩ�ܑ(E��D�:�|��nY}��jH�����XPF�i)��)ו%�K-(�Y����3 ��s���Y�0Dw^�R��΁��Q�bi>[�W�K�nɽV{�V^�� ���;L7��=D�>��@hS�/��R��Jw�c:xg��׆�lՔ�V|N�D7���T.�t{�H�8T�«����Z�^+l]E�Z�U�]�Y����RD��&_��V�n���iAX�'R��Yi������I���;ʹ�w��~����l@ib�$K�L�ƺF���L����F�Hu9���]���|{^'zN��v{9$ظ��|6k	xА� ㉪f�כ���y�Y�C�$��,*rcj���k�i�㸴{�ߐ:$>�[�_pP���D���a�K�JA�:N�鎷i_8�cz$�E�
�� Z"5I�E�� K�"�m�n�R�9���E^��#6<=�3!������f�˙�8Ke\8���ȧ��p��1������ �na�;��T�f�F]6�"4���F�Sȋ���O��f��D����� �^AuZW62�ȺŕK�QV��j�
�-��LP��ɩ����%�N�C)�p��#�'��ܫ'�Q�R8�Ԓ��2mo���7\m�����H��S�4bŐ����(����F�k��+��X��0�F�ͽ��0>]k��V��w.똫���ݦ+����@q܂yE��"��S�.K/??��n�/iXLL�D�e��x�\ՙ�Kb�uĥ���0� ~q��ȜK�~���enNK6�9�f�j��&���f%�Bݥ@��xzOT�nN��Z����g�CT��K�;\9*9 n|�|/Uy�\,�C�
���̏��'���r�%����OI%#f
#����F��-��M��'�[b~�f����\<�/�|m�Iz�� dh��k�ٔ>T`��c�qT)?���%N��&�myR`�\_=��'��{�w޻�滴K�6W�����D�QY��>s��/��#����*�ĝ�2)W�dq�h�?�s6�E��6Se���2o�*X����K���O*0�׏��^4}4��V�c�Ջ݋;
�m7F���c@)z�ݐ�M�B���ՙ�&t��N�ثE7��d?�i���^�t����*�f`'t![��9��!/]Vv�-M�"���f�e�e��<��)o�����ɑ��0�<\u��Y��N+l}:fyAC�<�!r�f�n�v�� ��e?�/7�	��<��ZsA��s�ʕ纫t�k+��ǻo�9<<�(�h{{[����OP�|���P-�x���S���u���}�>x��(�g_�t�w.\���W����E5V���s�y�e內�	O&k��yIە�+[[[��bgg�(��t���D��,��F����Ll�8��\\����y�֍7.8i��=Z�����J}�Lr�X�S�`S:���Uzj�O�8N�+�z��_��oOo!Į+��9�*?_�[�j�<W���L=D��8+�O]���r%��0�����z9l7�u��{ip��kZ�G��ѣGw������:��.�nyx�����!2�Ah;���{�b����/cF/G��Fg���t��L�zwr�8<94�p}l�ζ�+�Nt��%e�5'�**��DUkqy� ��+lr0�G���i�]Ǻ��e��h_ͭr�/�O2Kͣ�<�\d�U�Qc�7��9� �91�aͥ3���V���= à��
0����1�Q�B9Q 6�𢗜0�!����HPf���_�l���_�c��T�r7+~�"�g�\Of1�Zh��t�\�8H|O�{�F�vm��5w���e�V�.v�Q�� �2,wwwg�(�9�18�,I:{�DK8V�N��[rm	�����,.�|z~q1ˌ�J�O��ϕ�柭��E��?�6J����$�����_D��9H���%�|�3�@8�"@�p���a��8f�5JU� �I\V3+�Ç律PS.$%:�^\�1��7.H���pU�u��,]�I������[��W�_��0���n#�FeӚ�ZJd��j��� �6Ơ�����Gs���p�:�H��i�o]�M�vr��$���W2��taoll��@�7�d�&�6����&6�0�� x�c�'9�V�8�2�C���fd��+01p.��?6���x^}[r���Yb�j�>Y۟��A���i�ti�S�%�����*TGp
���g׸�����ھc1[�A��8%۵���Eu���v��� ���'G��E���k�ir��]Lq,�q=e��0;����܋��U�@egx������à��܎�ک?y��݋/�!�D��cUև~x��_�~��{�F�F� *-+=��ˋ�_�ӫ� �|٧빡G��h=\��F቟������d<�9yݢ�͢����,|Mj��x�X)���Õ�'m���_	.]\��a���%obR�|��'''Ȋ�*�$J�p�p���褫E.���s�*���{;�)!o������ŝ�O;��w�A�������GzjmF�q�Y3������2=ףM�p�D��I�]�QQ�<�{�����2�U�ŭ���EL&��ZuFc���1QhR�
Ldt2�� ���a��8fT�JÜQ��+Nc4��
�E�s��U�e�p�Y7�[�v��X���gy��VB�����������?Y����<���1�.�;DA�~�Ġ�Z�G�w���/F7�J~W�J�&�,|Kk���a8D E���''���u�K�)!��r���\7�W�rv��p�
���>ct�-gC�}���msH��I�(y��|��~I��|�|>
Rr�ݸJ��9�,� ��)��v̷womnn�6{��2� XY�%*b՞qc�u�J�'�Lc�N�����r{tI� ��̢_㘛�����<@��r]+��P�=yB�*�������?�.�߿��U�$t+��~��7Mumۥ����ܩ�/𧅚�T��O�F�C�6^m[ ��MlE{L��$��^�x�����;�]<�^�#-�']T��4������++��M&���E�sph%�g�����@�*i�ʽ�l)��%[^j����^=�'�����ꮭ����m�����A�T]���y����Y�W���J��
8���w=�U,T��b����Fǫ���!�$�&�Y�h?	��0*R��:	/]?��R(�$�����#T�%1����߽{w��I��{e�po��f��I'�ɫ� [�]_���NRnM�ϕNPW�ǣ�.ΜBJ���]�Eql�c{�,�Yڮd%6_�����c[d="�Ou�0K�l�j���ND��ӟ��ף <Di�a~t�[y]�Ԅ2
��U.��-��J��UP�
�U��-��0��:e�fdm��\$��v-�����t�9�)�(�9t��2�_�FyB�0~�+�R~)Fo��R�l��/s���*�Q���������ŋi�����@���uU�vЗw,{�Y��B��>F/�Ti����^(�^��.\�0W�482��y��6�C�G�����!��u�t��1*������hR�
[L|��[����G�������� �h��G���\J;�לM���P>3�暓�	��"T��h�
��H$�(�_
E$ׁ��ߍ�n����F��j���-�q,&��$F���h,�d�Y�m��SWV_l-3�W��y9���1���
�}������(�O�Ӱ�q,�grA��	��^�JAZŋ�'w����Yq������	rK�_�pae�~;��h��k��OE"Ӑt/�S��K�l��F�ƚ��\�i�E��r�xso]��k%�l����������L�">��s�	�{&�^T&"aPI)�,�EM��'���M��Z�W7VB��)
�d�{�1ه��0��]�V�lW�1�đUMz\�[p��C�\V�������;&-i��
�/߸B��^��WI��Y�&�|A����i�v3�*,���;��m�D[�-D�Ƕol_Ό#l�A����Fچ�wD�J��P����dK�Ƚ��yz�2�
�@i�8v]ئO���~�*�i��<��
xs�T�V����eU	��2����Sk̄��P q��G]N:r�8�h:�6����vd��" �:�{�����A�'�f�6@n[����[����
t�sh�
8���"E�`�f����/��d�e���o��T�����������!݌�I�}��^���A�pa���50F�	�{U{G�)�lWk�^M�F��Ч �]��9I�q$�t�X��D3'!�l��t���0;Lg謠����d� e�E:p"Y�f�OYMʶ�ʸ��Ɗj��<�ou�9ت�Z*��f�T��dM�:�k�$�@�u-��(�$-�ʹ�j�N���� �$��W'�bF�m,�.>�fj�����;���(f��]{Vf��+�[�c�r�bR^u~K�:��prm�����=��l�8G��~
�yK��T���AGuN�<٢��N��Z�Z�qG�T�����$�H��fO�j���	D������G��LMp�8m�=9ҪVJ�R��/�ɦ6��nU
 �ۓ��0��5&�2���e�I��g3���eE�'�]y��9��$�7�--\�Y�b��$��	���,4`oL�Q�46��2����R�B��VE�`���k������<�w�,����9רĮ5U1�!i��Rا��pS�9(����"�V�+�z'�����W��AX	��4;ڎ�,7@p����_gT�-���.5G�Z���C]i5�Hv��������_!x��|�Ĉ��'ۤ<o�wWߢ����t�Ǥ�vww�3ߎx*�0��*T�,����3�\&�h kk?�eJe��K������e�9SP�1#ss}U (We���o�h(,ڌM�+��`�Ա��p����e��^w��loo.P�[`��Nd��ܘSV�~JXZ�G''{{{i�UM0�tC���$o������^���j�q��Pܻ�D4�}'GǨ_��	E?��;�ڰY�sC�8����8�x1)��#	��-�rZ'�sf�KE�#ln\Y]TqCf�lkh������:��q+&��H�^ƭ�b��BM�|����0;�]��S��K��;��<,q���'���EI	��؏d������n��s�
�G������@�{�Sjq%��dV��!IG�;B� G�t��w�U���c�g)R|�]������EP�	¯>ܙ��b���laFNl�ck&Dw
�Փ�=��[-j��c�T*(+�/��M>0ǝ��O�<�x�r��U!@���b��*!\~R����Nrx��qn�lh�?2��UeG�:U�0Yۓ���(e���.8{��x��qz����C�88�GY�-8�¯��gx�I��{����)T�-���kH���m�K�5�ط���Z#�e*�c�)ȊM줩� ��B0�W��Dv��r�?�y/�
����3���%B%�����,����	x�To@���t]�����}��&g��L��3W�N�U�*�<���%��[v��$���uKu��J^V�ԙZ�<	 bDȖ��JC��WXI��%�E�W�eR@G0b)��in{4v+O\�}�f��u�����B'�1Ȭn��EUwT�r������Z��:'�E�'��:z-�2�:|k��F"�VyJ�D����S�Ay��j�t�N��c�?�khnRe�+��-�9�ROj-.�>�!�ˑi��H6$�'ۣ^5m���s����3��.쪷�V���E�Τ�Y��n,��Z='�,����%L�͑p@&O��nh�L4E%���%Zo-��4HU,��i��]+{ƪ���A�@���C�"�iH3��pl����<G��,u(�*�3�q� t*"�����;̡�mˮ�Z�	.���~jr�]����V�*����Qe��0��ix���e�(���UW��pt( �2���;���~��G#��<mK�s�-*K����꾪,��>_���v�kr  G�[Bm��u
�K�s_���$����h��p�%]�$Sg�Ym�0<��r4�1��"�G����d#{���KUĦ2H��8{ae�ץ�-�,�3�_Ԉ_�}o�(d.������e`-U�^/��K��'��N/�jq�>{���j_�6��U�YFc���?Q��*�e���\�H�M"?�و����T%̊��OYԶ��'�s���;�_M�_����{[
�Dϳ����#��-�t�+���S6�����ܔ���t�A�3���`uS�����xA����Y\P�@�<ܶ��<�-�t񅖥=]ǭ�kTu�ན-�u��� e��.E�b��gш���U�OJ�|w�h �%�,K&�ZJ� ���w\G$���V��p����5�A�X9z %&��j�B>Ssׂ��S��ӗ��Gm���"昦#H���f�r��&c+7� !
���#\[�Y���ԡjd1̒]!l�³�+)��JFU�藎�v��(aq���mXK~^1$[}ES,�!�]�~�"�U�L�P���9�R�O��|��!�9�>�"�	t��Ϙ�ARY��U�X��ϪƦ�_�3��n�?�j�}}��x4Q�Op��ٿjߣ�*M��N�4[��<������A��תg�}�::��D�6jr��3MM���P
�?�<V=6Cq|V�eK��rZ_����3,��Q��K���y�0s��ڲL�ҴjJ�jz��gZ@d���J�~��M�}O���W�![�7kD~�!���ŔY��%��ݕr(����Y��ܯ`<��E�=/:`�S����5tXV������=[V-��d�$ZQ��+���H�n���E��e��-���/CA	���eK�㰋S�F��l��|������ݜ�7���me+gYZK?U�=��լפ��^�KP.��%����BU2��`:�f�Z�iH���2�����������m�[�6�
rU�v�3Y�)�=ϴ��X͚��F��h�\��l�W虜&�s�X�!��/(���g���ן �Ѧ�+	�z.G��!g=Z�GE�d��yB�\��s�(u�-��K|V�[Jʹ7g�~����n�T�o���>�(��ZAְ\���n�x� "�.V˶�5�b�$G�&4hprڦd���k�(]y�"�����L�*f�h��Ӕ*m!=����1�֑�c�vÅ%�<�j䙊(�K/�ʴ�z��*F��%�}��T�q��S�e=�	e���2�M����"%�y�`v���Ք+`�Qf����;����>#7mu^��[$�.Re8��U[��Rn�� ��@��)�F�j����?ᙝj�>�:ϼ��܏Uy�y��ڪ��������*�l5f��
M���la�+���s�ZQ|�e�ө��Ԫ�sH���Q<hV�SG�'����>_Ĕ�l}Sv����*��>w��Ҕk ��r�>K�f�����/qmR�ʇi�pl�̐�D�IV!0�=sZ�4�K�Cz���r��f}o������/R�~�g�{�)��:famL��e:��ϕo[����(ѳ�{F,��I}��%@?��O���_�J ���fEu�9ES2/�n�XN3������Cԧ;�z���;#��?E��0�}@U�^�/c$b��0\[[�\�t�Q��	o�t�������	G=1|�epޜ{y����֚�|�{{͇�."_kKa���8�?j,��A��z�.�?���ͧ��Y�#���LVU�����RU��\,�yj	Ͽ�O4Y�j����d�{�HKvL)?��9M�������~������x�V��:���P��W�K�6+�����^ lV<����]l,k�� [��(o(�;����S�@���/��𬮪����W�g8G��9�������'�w�e>A��<ڲ.�j��~����|��噿�B��g�QM?�ށ����ȶ���oi;w�=���l=���|?{�NK���I��$^u���(���r�`dY�    IEND�B`�PK
     uK\y�ݥ�  �  /   images/2db9ecad-5c51-4c64-ac4d-4ae785eb4e5c.png�PNG

   IHDR   c   �   ��   	pHYs     ��  ��IDATx����l�u'v�M����:��~9'D$ F�� R�xDZ3�?̲gͿ�/3�7��%{�f<#�3�(�@� 2������~�s��n:�{�[�J�rx�Wu�=������na��LKB�1���!�քq�(U�J�0^Ӕ1F(!~��Q���g�a�w�Hf^�(b�!.L� ������ �C���(�%������0>	/rM�> ׁ�񃷤��
����¿��B�~;��Q�?���%��*��?���T���Ns'l�8��z\h#2��8v|���1<�� I�@j���A�h������[��\�h_�����u�
��Eʔ0�p�cpy���S*NW�.B�N�#Af�X���­�� �$��ОZ�D%�R��U�z'W,���E�j�/�A:���l9����
�n\+��5��6$	� �?<�]�6>�Y�n��ԌJ�<QI"��@��5q�pPw�V�m���d�go�$=Q�v�[���zEev��M�B��@���I�:PX�@�� J��no ��󑝨�qM��q�x�B#턎B}WDTYϸ�;So�ѯ��S$~m�����F�W6����-@L���@�ɶ�2Q��VE��8e��'DD�o�z�I�S����CH�p	��PV�TÒ���j.A�����\_��o����¦�\�o����X�-������u�á1�h3�x�ŉ�����nY��2m����NJ��K�tR~X�<^�n�m܏je.�ϞX��6j���(���|Nk���{S�2c�`���2�V� ��P|c��ȁѰ&�R����v:���ވ���O(��z��к�/�,�(k��-�2ў�/�|ZK�294t�"TYmr��
>�*P_�w�$��A��;i�Hڮw���rN)��"����>�]����S{O��hRU������E�'�:�
���y����eci �{��91­8E�@hΐ�$�:�De�\����+���;�Ju/m�'D{֎O����@p?л�ψ���d�H'&r9�s�\��Q��@�J��sK�#zkn`��i2f�@������6���Ӈw��=6���z�~Py��Vmz.{~����(	
#w6�`/��96�X��.�@P����T�*���rQ�P��]�vE(���c�&"�ן�=�#�Zc�TBA1:ԝ�/4�G�����,�7֛���0O�B��y��H)ai��
�'���p7Z�a҃'��^�٧M�!I��D����������^u��`�P=Abڸ)�l�>^.GY���v���%��$5Z���+����w�thg�`5��Ae݈�R���Rp4�Y��TI&�ha�*F���v�U�^&�P�A5�T�P��������j0\WY,�ɢ�W�:Xڸ�Aq��*!�X���V&ʕ���s�Z��:��`�pIt�ZŪ!�+��`I�G��T7U(r�	��<5:0<(��_���2/O+��ݴ�� C�a���h��Ak��l?�^|�u���a���ڪ�EjD�hČܯo-�- 1��@��͢������X�~�jn�n�/�&����R��#�e.��i��I���A�$���Ǜ����1�]��e����H�0�(!�͠})hC�������B�P&�"��`>_��v������G�~���,9t��:3j�����@�Ch��U��(\��ʮ.s76�Î����*�P/�\�q��*׎�N[$�a�\���:�b�z��D=���W:>�Ա�++7��}1Y���%�G�A�N������ ��b�T��8�G&\ɭ?�E������둪q-Wk�O�;w��u�KP9�A�C��:&�|Y|i������Hn�:z}s7u����������&��6�K��_�}�p�u���GN�+�����Ԝ���[�)���V��Y��eS��VCߍ"��d�����)R�M\>?��r);=�x�2���Oo\��ۃ��^�D�%?����N���u}������K�]#�B��9M��������Ϝs3�+��O�����w��m:��}����Ź�nI��{=l@T�	��1C^ �D���d,a�IV������0`�Sw l�����ꠣ�[��v��{��>$��(!L|D ���Z�]6�����f��dad��>�i_��dV �)��ab�^����4R��_}�'����u�]��3�F�s�.]Z}��_��c�s�{���o�X���{T:$�#�'�xrwu������^N�@�$A{ɐ$1�bF��Ƹa��c�C�j(C�@8�W�J�I$I
�ܤI�ו��v�Y�SY��V��90n�#J����?�Nѡ� �sY>{�s�N��S���'{����>�u�t5(&�l7T�����׮݌�s1�#�����-�Z9ÞI�j�P���O�T��&���<��u�:
�{b�:81~��5v��.>=>��k�Y_� �t�S/AuB-��Q�DN�� �[ώa�.N�\$d�I���ns$RڋY�Ek��5W�'Fc_ Xf�Ӡ��5R�r3�S�R`DG߈�`�թ�����A�����N!����&E�4�\	1��ҙSG���'�ʚz<�A
�֞
��J�����N/�������sG��a����G���#٣�Dy����|�M��D�x`�TG�m�.KT+ǰ��D�A�t�դ������`�jp��l���@iQ�2ȥ���UR��r~~���f�(���GY~�	|�-�t'��H�5�KS��q�LK���ݻ����Ok
ς�S���A�Tx\��}�X?q@��	��Q)�A156?����du^ʐ �)�����cZ����.�[�O����{��i�<�l�)�ILbH����*�)�+^�Q'W4�ЀȖ[Fu�9H�a�!np�9:x&l!m�+��r^�x�ɪd��=�>1z�h��D���N(���[�ե���ho�Q@#,Q/Fa�t7���g�����y�����/e&�Q�[<�齏� ��b<.<���b��d��-q$ԶOL-|�v�:_]o�E�� g0�6 w�ؔu�����ZW޿����f�"�6�`�:r.!yԩ��d�-N\�:~�2�2t7��[ac-�o�p��kD��rR�� .|�ˈ
�y��	T))Rr8�(y���'��b7e�L�xv��[K/.��v��Cv!��A��=9u��ď�9�$��j�F-8s@/aW!��	��_0��T`y�)-%�	��Ӽ"�p�{�O�����$�fc1��^���ܕ�����8�xq|4tC��@	S�q{��ѣ�3�_^|�˧����:ԁ�H����m�\����҈"��־gP�5F} ��  �A٣���d�zO��~�����4�~�7���y|ᱱ\�|�Cս��&	�1%���'��`?���(��;�USP�(��qg"?2[���jM5@� p�nK�-�Lń(5��$0ŁI�Ax4&)	!Z���Z��TW�R*�� *��b���:ۯ���g���~��3�y�+%��b����7=R�:3>�i�C���瀰�ك�~�f����ѹ�^���?�0�h��(Y��[(�1�a�pa�ȷ��懝�tS�N&��4�޹��.i3�	�&\cn U!���LP���g_���ZX'2�c0W4C0�:��;$_(H(�<�� ��n�T� �]|1n���0��h�˒���3[�M8q រX�=<11�Kg���N�p��#:��6Kf11�_���e��)�At�l!7��i�x��@�e�]?~b�8�!1�������4��#Sǟ�;{sy��d
#�jʎ(�b��AB�$e
Q�O�6�S.���:�'�I��e�W�^#�X<�˴�B�E��:�B��U�	�����'�N\S}�6ٌ�/6eV,Jٯׁ1ɅBۨ=������8�\Ɋ��ұg�D�&F�����˒n =��ܹ���V7�JSLo�Z�J�ȡ0�5�ĩ�þ����2r�ш�.`�޹��w__K�}�d"E���_���~��O\~�2>q���Kwz�Z2�3�13�g&��zg�2ut���핏޽3{dB��}/z�c:җ��Ywe0锎,\��߽r��ؔ���IR�J�R}��s{�����S;����+�F�i�4%���#cӧǏd�b1.�Wf��������Xx��Ek�n��=��M�e��y�&+�Y���\>�;����؈W ��N�KD�^2Q����?9u�4\�[_�տ��?����3������o��h����/������a�ٟ�ɿ��?�>6۩�Ч|�NӅ��kǟ��o��;�8��O^�����>~�"Gi�X��iqj�|n���g�<��+?�����Q1�Ɯ�r��g(�Tn$�c�A���L�H�T�rsAH���j%P;j!&˙j�7��v�R"y ��q p|T ��K�ۍ��??u�,�& l9?��o�ƫ?{s���13C��P��9�����r0zE�෿��?����W$�`�nN����w���  6!���W�y���?��Z�o�f��1��o|gdt
��	�K_��{�V�g����#��΁��3�gBYj��}K˼�%�q�����BJI�4B�^�@��C~T�1Y��R�H�^�`�JT�ey)v��Vaa���J�������Lr{S#�#�ai�{��a"xύ�Xp�����]΅HJߠ:~�-�@��`.�g����,�� �#2�X�'��� Љ�;}N��g���	�8�'��f��:>���Ea���ѡNS�&d: ���IV%��1��j���h�"A<����b���^���!�t�}�����76ɓ-�Bw��A��>�a'���6\�3
����^��;6��2����	��~��Z� ߔ�%#�Kn5��I�s=[��;��[<!�oˌ�w�nW@]le����|���.Cd���p{Kr�d� I��E����Ό-��j����M�+˷��@��f��p����?���O���_�f��/��zg�����D��������[�����?E\p��+����w�`GF:�j�`r�ӻ�W���;_��/=��o^}���Yɏ0-��\��{�����!]��ꃿ���������=�<���V���:�#P,�W��*`� ZB��ڊ{-�h�Ԁ�GGA�P�|�[N��o׮<�^8;rZkn��f(2[Pk�*��k��?]���,l��L39sj�E�On��/����㗝�w�֭+�܊��\1�B��-���W�������~�_]�;z�ƍ���{�N<���@հ����jA���/Wnܜ��X�����뷒}yt���w��I|�������vuy���K;��O_��Rc�<1�qX�V2�bK�\y���l�Uh��M!H
s�X�l_�ݾ�4��N�*�ͮ�f;�MA)�4i�������*?61��zo1Df��ڲZ�l���/މ����)�) 764�t�ڗ�G�+W�
������� �\�뽚Ϗ����՟���#���C�z .u�՛1맦U��?�}w$7pS>�wOͶsX7�q�NR"���}���}�Ȯ?���+Ȕ�Od)l-��M��on�<|o�O=�7y�E��e}b��;��}����mFZ;x �0��m1x����T�X�'�[�{��?��ϟ����k�:6����~��;�����:uM����&ˣc���d�je��2rE}? ��t�pD��&�����2'�B��S. r������I�Ç0O��c��L���� �aUV�	g���<�S�;��5�IF���y%!x*t�Ip���_�����'�D5�ΙUHHrg��_�|��xg+"|��lNDil�U&���'���f�K����l?6s����ɠ��"��ڠ~e��;w���-!c��{uXo����Ξ=��8�g�l�=�$�4�-b�Ut����d^(j!ڑ�`R�j���%̃��I��4��N����9�����D,�b2N�����:�^�a]�R��\� &�jY6��֫7�+�̞?:67�灬���{׶����eY_��.`L��l1�"N1!h3t���!�b
(��t�GM�ye�����-�tWvM�c�l"��.�I���{��'�]T�`X���:��en��`�<GB�c=� ��Sh%�V�E�Ш�Y�hXP��4��ɹ�i[�!��)v�Y�
�iDU[E����NҼq�
����0�Wج0�iWp!T

��L���o|�w6W��G�M賈���"1��é-BXR{%@��g�z������L�88�
��A\����#<�
����J@�@�Yh�fEr�ې}Id%�O�^��6*���J�Ajao��h �)W"���ԗb��;��NP,�<w��I?��\���3�X&�\=�we%ރ#R�����j�|`ƌp�,�5S������ڕ�=��.K ����l��$�HA�*�%�\���� �a��p���Ѭ&����L�ռ�>83�'�[d�=2:��=�����С�r&ʐ %c�����U�kw?�y���K����0?��=���ڱ���a�Ag}9�\�ti5������r�8������
��� 6��	�2��Ŵ-��Rg}�������� 3��/LϕY�%� ��#a�i�4ӶZ���mj�[�Ɇ��8�ù�-PƂq��#N��O|�E�{��1 @��3�4���������1�+��6�(}���4U�ܼy����Vg��کg��:>��w��L����
e�1:]Q�����닏�/	@N�-S{m馌�^�\%���X`-���� ����m�@8�n��$��<��J��T�ub�����YעJ��X�ש-��$�HGmVkوEE���[ϱ%O�)�$K�w�}�P�ĸ�j֕��J�>_�9v��a�>\�ۢ<��vZ����z��Լh����K�D�5#�Qg�$tE2S��@`�-��i6��^:z���#���y��e"��tG�zc�������>p}gfj2�Gi��|�@��u �c,��ҙA>��[?~��w=���.H3lж��s��� �P�#z�J}2X~�$Yq��ѭ�t���-m�Nˉ�$D��$�l���`�,��X4�<�������>q���C�6ֿp���7����B@Ĭ�~���EKf�r� ���'�Z�0c:�����H45���--_8{�dKy�����|�	�ݘ?v���W~�rԋ�q`y�aO?z��ũ�C�u�/����kK�\��$�I�4F;W�0̹ 	̺�����&Gl�
i!����
�v��D���NK�6�I�y�@�C�hy�坱��������R�Y|�n�YYf��#�mo<v��s��_���]��:>�d2	���7�r�a�R{<�-&s`/#=�֝�`Gl}����㣿%����g�z6Y��0H���n-8&��ύ��'>x�M{�.�Աc�OK߿���sr$4����?x���a#r#�Į��y���䌰�T�ڮ,��p��B5�Bě̱��"xd�C�n��7�U�R�*A��(Fř��J>wk������Q�)$���w�۷�`I���vZ{O?v�o������Td�^�T�1��XIU�@�@�:i���m��ͽ���/~|���������n�\1��(�	Ǌ��\�Ǵ�p'��������$)A���T=�Wo����I'
��żW�N�f�;ĳ��5%l& ����r5�܅Cz2���N ��щ��J
?f�l0qe�
e�� $���nT�����S���}�[%���SR�S��fM㈁J$��΍O��n��|��G��k�b8�z�),0�!2r5qizq�b$w����GO3�vqtdjtj��m�$P=�a��[8�V:�~�ϥ+��#���p�Fpkr����d+�b��Z��B<QJ]�̕���0
k�VL�@�p��z^����:�-��<6H��Bz������Y��F;��� I��������fp�69]�j0R*��=����pr�z�ft�Ir7L��� v8��'���w���Vph�F�a-�� ��J�%��� t�^��Z�V�j?��ڙǧ��z�u��Gs�өs�ۯ~�����x��F�1^���~���'�/�^�Pn�>hM����;���{ot��8��|��]�7��vO��#�%>�������4�����a=]���B��P�(�0�e��0���0����z����[�o��ht�r������I$`*������ ƅ�b�Tr���cS���B��M�8�W�h���Y��<����*#���n}g�Q���G+��'O������I�m��d��DO%q�d&�|�tϰ���q��1��7E�V�����Ւ�Y��$<B -M��*�֠O��R�hLqq�ѽ���w�+>YTS% �+�q���~1�r�N~�G���ËSN�;N0����`�|l�T��1B�W���$I;T�='��;Q�ӻ7���1@M�g���a�h�z�?oۙ@��ȧ.\􏜝Ӆ�K���
��S%#�`��ދ�7���
	��Pn��p�&�UI�7B�6wV�R����Q�
n>�O���Ϻ��9��6Bb���~�[[b���./��6��\��f؅����p/jk�WXo�/|7���^��*N�#ɚ�펉�Р�D1���لA\�"p+L(�Nͽ;Wwr=@�B���DG�<�Fr�5�Nw�i$�+-���h�8�����ii;�BLJ���5��w�nl�}E% ����ى�B��Z l�0�cy��z��n]D��5��������Kg<�HplRQ����j���VP��M�x��mfj��@�����]d⦹��o��:�hT1V�ߤ�O�}�D1��Bɍ�s	(����'�J��b,����x��$�̏[Դ��������k�-ї�^]��l��#yi��9�]�aH
0&C��{،&)|��]j�a� cr;�ly�q.͎7��Bri71�kX�`C��h�Ĭ2s}C5���тRRdm��|� �V*B4+1ơG�t�8@#t��\�| ��ʬ��d�X�8��Ͱ����mt���f��ı#�c,��.B<l���'Y�����Z?�\��=Ic�sj��
&���	@OR#��r@}�ᤛ�]�-$L����Ҝ�\ő�@e��ȑZ=H��]5�����!$3�-�T��Z`�-ܿX�����
�Mf�AU۰�M�0#5(�����8�Z��#�5z $݁��FW��'����x�Vl<�Aa��Izo�A;Ą���f�laִ��B1��SyW'������ȝF�R�����ng�����:֨`��g��(�t1-4�ێE�:�[Ug�����F"�ڀP�`]ŝ�d	�;�t���&8�$�a�=�bh�Q�$�2��#UJ�,�.�RR��rm�ͥ���c�h'5�d������*ԇ?J��g�� �Uֲp���+}�0udj���׿��U&}��̩����>��6 E��#ؖge�w]llz�������/���\;�A��<�شBMĐ�pl�FS����a�e�e4�	*æi��Ѧ����	�����L$���LL�^���\'5.���T�X�h�xa��'�ot�Iq�yY�(�W`��h_��{T �M��k\��� 9��V�����R�O:����J���k��/|Ը�ű`�4Vi��Vvd|$�U�Ի�s~�RA+��kV��U���� ����4H@g��6�у�Vl�.�$�-;ncD�l���PY��D��\խ�H���ĩӕ���������@�{�E3j�l03�`{mqf���G�W�8l�}I�E�{1IF �J�\PAQ�QM)� ��i�h��G&;�>��Nl���!��4�d�����ݸ���_�(����x��wH��죂�ѧ��3�v:ѩ?��S�'����Mzx,IM�0`���8c�> �@�_�@��Pۧf�w��6م��,��М����B�V*<��
'��ka�� C+��W�4���$)�̜l��0��M.�x8_�z���/�}b�J��=��P6;��-���'c��������~����}t�:�ݳ+'�}��~���ߑd�w���_:��8��q~&7}��I����F�ŮǱg7���q���9�M��w?|�Z�9��ā����r��b7�.x��hlö96j�հG�f��������������a:���Bxw{�������?W�S1�b
Vt�N��r�����|�������)l+S� d�Ύ��#A�Gd�kY��*�T�����ß��`�����h�3�~[9;�ݷn<���ѣ'�&&��v[�1,��q�A+U��CF+�o��ퟭm�V��;)����h�_����BU,������n�&�?[�2d�Ҭ�L�
��T�i���t�rp���k��{������[W;�o�9�Y_&��^|<k:�> T��zMb�t�&���y��6�X�]�/�E[C'
>0OE�8r��O�ܻ�z�����k_}a�\�_� B���WW/�>�|g������<�P���Q)f�iB�m�`��NKŀ�\aF��7H9�I��|���x��82b{�7���m6�
Fa�]1_R��"�A�G鱂X���y~r�jm�w>��S�/�U'y�֫���d�����f��Bu2L�'/.]�z�+�p�i���ʊ
�v��D���G*�)t.u�T�X�6�7�-G�۵�^�u��d�Q�a�+���ų���Vko�a)M�L�cO lh�B������'��6s��PV.����*���*x����F$o�C*̕R@��Ħ0ŁZ�Bz��7>�،�Q�Q�������n>����\�[o���C�����?hȆ�>��xy��`2�����W�f��:]�_�� fϪ���h��ltv�d�H�a����^�#�'���k�EG�>7qjqm��8I�D�&s��;�����ޝ����MS�z�T���M�������tvO~���,��_
�)���0=
���+��Z�4�P��ʧ�92޳@ݖ4��B�'�HFs�֟s[������wK|	��7��o�)vu���*�)Lt=6�ġN��ׯ��vg9)��v�o�3�ݼ�:�P�$c�plP�7h} �Xղg�lO5�S�۫���;_���ٹw �y��Ϧf�X�:S�o~��?	�X�Q)�8g*�H �pS*���Fmc���K�&tŉ�}�a���(�2�f� e0�������,���"mf�ǖd��QRI�.�٥�%�)&&rtθs��ikZ1�p�︾[���+��pU����PQ�\i<c|��8��H[y�P~�T��E,l��0	pT<������f5u��l���/�<s��CS ǌDw�)�c��:����iZ>H"
O����c������~��yߜ�L��۰ɨ߶cQ��b&=�Ϫ�k^=,�@�ő���.RC���He)��%h�zl�C�`���ܙ����}}px��)���������..VJ����㳋l��^M��(�2,f����Jg��Q���h���p�ӥ$��;�v���F*��wmm�&�}<�	��R��~�$�(O	��BG8`sj��������ܻ�&^v���-��%��*�����@�V�e<^&,�P�����<;Yl,���F���yGМ�H@�[3�N��+��R"!�E�^5�9?u���1�L�����{�	G�*��xo�/��,���(-����K%��+���֚ �q@�0�(q��� :�x��������ʞ��k��>$���T@�Ҁ3uN�)�f���xL�}�4IIb�q,�=���b�(��ʚ7�Iu�h _1]iz�ظ�0��O<���x���i����n�ܨ? �W�I�~=�Z"��ڲQW]E��AHbu
u��d�Uvz��K)<G\Kb���dAbG%�e�G�J����G�*>����#�r�U�ƪ�\��j�Q[�UmM��r�r��L�;�ƾ�+����dG�/�N���z��ށŢGG�l��`����(�>Y#��×c��@;p'�/ܾ��F���ж�Hвl�D�;nw�$)�h��a��M���t{�OY$o����@�<��n�z�^��	�̖`���/0�g����g�� tҔI��(D���H����d=��a�%�RϞNyv���8�m�;���3}{?�6C���Y~h�1�n�\s���O����bZ�p�H���+���0UK�<	��S�Ţ�dF6���!��R� B�T*jI4P?�F��K�)�=b\ش���s��YHBb�D~�������ӏ����
��
 ��2�TL�<�p�*l�����t�nspyx9�AQJVRv�`��Jh2��A��]\��Ɖ0�+X�P��*
(��$x��E��p���a!�GB�̇k����� l$#�d'S	��S¥B&��䈓�r�J}�����%>�v�	��=�k�
<s4 =��^2�L�^��1I�V2�=�c�Pi��NFY�vJ�6pPc�=O�d�z G�O��a�
�~���/������5��C�+��9�`�� ������/�|��k��W~��hS��S�ɉb孇�kx�P�'~������}��A܇{N����/������� ��E��/��l��o~�Z�OR2ʊ�~�K���כ߻�����rX�gʱ�q<fc�A2�&M��hB��}S�P��,���[�|o�F��*������6M�d!�y���� v�C6K�Ѓ�!m���M��p��;&o�_y����~�B|a���t��ڽ[�/��p�0�/��r��L���*�/�?�ow���v��=�87�����K��c$���K�����̍!�'ZO��������%n@{�O�J���^���K�͕x�M�x�
��v��&/'ݸC�v�+�.L_<q�:>��`}��o�C���\-�l݊E?�'2�*c!�w���<�M��:��G͌�6{�O8`V-I D�����\/x����8'%����ڭ�8Ϣx���w���/�JMi@�� IW� �����s4�[�����q<��$г�\��]7e0B�$ ���5RQLe��vԣ+09pj��X���p�_P�vr���$��Ս�f=1u���������h,Y��Vb�E���?c�U4���ͳ�;���s< o'�Hۺ�b�*m'�c�3��]��T2R�P�K�ž/��
�y�P��;��Qh�����3�#��/U+�i<?����Bubr-�>p��I�X�_X�-A\E��'ϝ���,U�^VX	v-z��SX��5����M�{�카�y���v����=Z��$��h���,̳�$!��+��8<��Q1j��&MRl+�lY�`E��4c@�nܹ}���_�����Kq �+����KǦ���o�������|��\]3�N|�;��W?�����Z��i��o������8���[����������}c�\��^�y�����/���b���Qr����|���~��aC8����{�w��o/��ߍj;�q��3��*�xX�+��C�#��zw������x�R <��߫%$,����"��n}ֲ�#�ȁ�G�?�Y[tȜ9!��5�u`�s;E�ݬ=����0�3q��$�����;�����t���c�6Wq��X��t*�8�9I/�+[ok6IBi���q�pm�?(�:�˹����ҝ��� t*������ �:屮�r@>��,��R�W�kǫ#Gň�2��uo�4����VO�Y6���'7k�Z�	�i@�p�(esd�����_��$xКy�A�<Z펫m��;���*�ȱSp1JKcci�3g��d�u��*^p��n�?5Y��,y�@�[�?s�q[l�[�^��r9�4YN�֨�[��OTF5�bR	V'}��0x�Z{؊{#9֫5��N����:�zg{0َ+�V{����v�q�LR�?'����pb�;Ь�dg���tq*��o���ƾ���SO��������O�e����ƛ���u�b��xu�RiT��xv������ەJI�	&S�n�������8��[�(���W߬%��5BH:h�n�oĭA���ݗ���oĔ��B�X$�HDom,�Aɏ����rStp���n/G��r:5r��
��e�>#���T~�ԙi����Q:̏�l�AXP���sOTN��p�ܺ%��;����¥�����G��ݛ�.�p��6W޾��'u������ߨכ<�ٓi��;n�7~�W!�so�7�:�P�k��&�+wv�
PV�~��J��7V�o���𛋇�4���d��,#5�moF���l�����x�7����r�g�sFH�|���A6B?������� FG��3p�N�C����ar¸)�����ss:L�f?�`K���F:qA_�N���*l�#kǵ�o�a�N~_�UůЖd�,���v�R}�:EZ�i���fZ��ܛ���������46�NO�V��S`=���_��������'q�q�9�xZ����c�I{D�A�KpN��inQ��̔�A���A�E;�$�Z�u\�d�(M$ľ��3۠F씩,i5�����o��7�a���%K{x[��A󵾷����m�>[���_Jx"����0��X����2֭�Rj-�����[�qv<t�*6��ި�ʵ�=DG0�7~��kKn-��μ����+���7ND�m��D&�=0� $Qǘ� 6W�)η�^��@����>�(=��B�q]�"`� ���Iz0.�B�G�N2
��טMbC#&���	����t���Ώ��E�t^�8�`��믿��B]�c,)�7�6\;�@��L4���{������ƌ���-�,��q����|�~��q� r�{�W����aX�0\�m��n
ש���;&�J`ʋ1w4Wi�����t��|����vԮWJ�S��;u`�>ɛ�Rw���s�έ56n�w�n��f��G��2��Y.�DV��^�m�>/IN
�k-U�fV%�t8�OZ!iZ8�ն�Z���N-;B��S_�`gc��P?hf[�=*��Z3;�2�˪���s90��I�~K�}r���R-�HFF����7����������V4�����6621�����,��bW���t��4@*��&&�s<�Wä�(a��a[�gʦ�l�U�O�z��6����d5�-�����x��{�3�'���e?��
�vП��nl8��f��Ҏ�c6:#��ऱ�&C	 ϥN��mԛ�t����9|de�.i��	%����8�h�:Ã\���ڹ��#�~�G=㦭r�,Ϙ�ʚ�l�J+����@�	[��$+8@��m{36���!z���!��
�fH���.$E�TLp`�������G[�Kp�ىJ�Z�v��T��U�-= �֍RNt�P;�l�Z�������o�ܳ�����S��#�+W>���8�p����� ������cc��6>샃�R������'��#%v�ds�A��𴺵�A�/�I������>��^载~�J�R�ñ�U���"��P�m�Ȍζ����,�!z����2I
���C�����{*� CpX8�� G�x+��NC�ġ��a����&n�*,#A�d^�
թɥ�w_���<p���/}��$��|����>�c������y˸"��r~1%�^���9G'��,ǒ������̃�|3���4��TDq�����������vLc%��#r�1��^�'������`�&*�Ҟa��P��� Z�p �ƀ��\���ܞM�:o�M[!Y���<#�j�f��\;"�)��8��D���|ik}e ��3��F$U�`�᭝�gfΝ=sƫ��_�}��'	��2���/��DI1$U��6,�؊^���],y1�*�Ku�������M><��G��ݨ��ڃ6�(v�[˥CB���o�L���(�\����e����Q���$A8������G���켡���sdxf��O$&lw�F���}�F	IF��/�D	�^��7��h���Ο͕K^Kt�rē���"��'Q�:s����"Ì].��᨝&�����Zc�;xX�c�
����m��q��qy�}!����l�/;�Ze� ��p;�7�5����������}(�!M�����5�T0�	`R�\Z����;o�9d�ׯ��~��9��i'��N7�����:�e)�.������)>3.;��N��^�ڛ��bN�T��lX���W~�Kv�����zZ�sSͻ��bXm�~x�!w��U���tl��v�X��g��T�d�M�ѝ�)=H��my��sRlbV[n���Sc8 �ѱ�� uv�P������ɡFX��L�.6t�7FrLe�Kf+٨������i�`0�Q�"��sx�D�F���l2�5��lm�$��m�ٖ���������r�L@�W�V.��4K�炟w��n�/�S`���g���D��PXb#���N���Ͼ�퍝5ꑅ���^k���3��'�C�W�
<*%���!J�>��3̐�3�h7��g�<�!*3P
<U��dPo�2O'�ij�T��Y���] �ށ.�!R^�3��tGe�2�rp~#���� �#2��|����G�1?����Vs�?H2�v�Ps�!'i��w^:��rhq�8��ǯnl�~��/��ڨ5��-�چN��Rp�U�-N��c6~�3���dE�(�����ö�Q��t����M5Q�ǦM�?s~�8��ŀk�Y?a�d�K��|ty��__ r�Ƥ����M8\��mh�*I%q���-���0�vP���>�bk�Mc�  7��\�t��S�;xt:�|�s������������ �A�;R���=2��GDp}23m���;U�T�T��@ʹ��Xi��-,�`��<��'g_s�&N��0	�j̅џ�-{m�4�Jt���R{���; BK�0�5�����h�?/O/���i��Ϊ�V8±��R���S��e�N(:�ǂ�7P�|�˻Q��I��7�D{�'�NmO��a� A�M��;;�����ӑ��J�����{@v{U��f���hV�i��C֢;-��C���ٶu�',� �$UOٓ,leJb�LbpN�Xg^�`�#���Đ�u��-鈜æXv B�����\E�Ǐ�����v����}s��ON���^����PC�CRT���*�+a�G��ud�zmw����
B��-5x����{N������Ցۼ?�ä�rX!�q^|Vb�9ɰ��&�m��2g���+�����Y~��]ZN��q8|�N6M��h#$q �F�ܡs�G��>|h��ǖ�<������U=%9����݁+��f�B �\-�^�{��r�`'�����]��:���A��1�A�N �9ۣFf��߷���,��2�'�0�u�����Fx�_0�,@Yo1�_gg�0�K��p0@`�
��Md6�DJ��Ԣ��TN������{Q21V}��/^�&��c�Rۆ��Y2��ΨdJmg�b.H����F�g��4�r{����M�(����3^6���q��Iyj�k��l6̜��0��٩��V�y���Ln悴�8=�� >�C��ILEXL�����o���`$5��6��I"�w}�ڵ;�_[]{���4?w��4�~��8�W%<�gė�l�����J���q��������T�p ,a~��������L��k�Z��b�"�(�2`%� ���&2UD�h�7I:Щh�.�]�9���#��}�� =X�e'	p0��WP���T[�t|v�8^IV��"��g��O �sL��Q�eG�~���/�8�R�p�v�u�����QG�<�E�>*���f~�����f/0���nv� �̘0�I���ű��'�z��F���w^�V(��!]��+;[���i����DZ��_��>���w�"�ĭ��?��_���|�������k����B��������>$��_���A��O>��@a4U_��犹��W>��6�K��<��gg'&�_�Ѡ�[K��`��H�.� (��"ZYi�!-��L]�>�'�7[�v'���
�\�h'�R��ȅ\Ӱ�kF`A�	������!��0j��$�Y������S��^���z�Nnd����ϼ��]��8]�x���?���}�4z0�/��̅������wr3G=���-�7�h��=t��-�M�$����w���^��o]�]ݍF7�@l������z��a������pXa�4��B�c�FC���p	b ��zo�Rյ��g�|����ܗՠ�� 
ݹ�w�9�9�;�79s}����k D�5;?��Sww�ϭ�b&3�����y�����o�<�U�K�
�/ 	�L�͸�b����UGxU��z;����< ^�����^��]7}9��G�����fBYVI�>�Бdc"J6�(��� � Q������8/�H8Ιf��|���!U�b3�v����߱�p�����(����M����-�SS3�9}�?�(���C������f�{;��q_�O_���k���':Sn�����Ս{�m�k�!�b����@E�-��7u�0��#&rL=h6�����qIڱ��2k�6��ɁC|��P�%F�ǳ)G�Ό�a���(XRq!a^�������H����:���mϘ/�TK�ygKי��eݚ*��-���]80�����5>;1u~��C���B�D��ѹ��+q��R^.�N�/�.^Y�%��2�h�MϞy���ަ�A�yx����S�N�m���R	��X�0�������H��V-B�d�1(M3!m��~Ju�A$�;B��VDB*I@�\�>�%�e�AvLt�2ԗ1�Z4�X�TǞ?�¥kW�Pp���������͝��]>�S���?z=���q�#��B�K��K����N�&�^|��
�h�������3�J�x㕤���J>��s�s����:���<'���'�?���H_��\)�%�H�k�32`�h�bn�>c���ƫ:(�U�R�W�8��5���Ɇ�Ҭ���he�s��0�8쟥��{���?vEa���W�%)s�D��/Y���^�� ��P7u�;!�6F�M�a�N'J ��ap(�t�!6���U�Z��@��\,�Xβ�~_·I���q@U�?C�#�S
��h�QK�m�����}�w�i�>=8�e�A��3]E��ĩ����%�m|�l�a��Q?���!9��"�����a/"��ȑ \�@qx�4J��G�D���ʯ�I���ORɕ���o�6��x	ed�d�ڛo����6�Ib�x����'�N�Qař������V��ME�}]���-��ʑ@Z����{?���	Ku�~lv�}gg�Bv�E5��\m�k/}U�"7�:uWWF�xQr�}����va����fG��2)<$C��ha�C���7�Mq�/ͨ��~-��VL��P9䊦>H6N���EKX��,��4Uy�݋!bt$��~i��LP�a�^��4+�F"ѡ��u5]��	���i��7[�G^
���z�v���%1�3�����U��u=�f��E�*���[1�F+��o4�x⩟���g(�x�ӣvqe�4ݞ^8��l�Q�Y&5�\�ͺ��K�A�誺XMK^�a�!D�$y;0,E�.��S�ڕ�����~+`s��T|�zL4_DP�APO	dKP��)'���C K���Hv#�k*S"%+X�$��
3�J���q�~���U��c�D\·�P�q�8����]8�D�L�m�T��]/�K:e�B~�<�1�0a_ǉh�΅�ke��#غ���ں'��,յt��'K��4���}���Ά,a�|���G�P���GV�����\i�n�6�9�sFMSŸA�E�	�V���r��MӲLGG�5�I@����^�,��n0VЌ��I4���G�e�O4HX��T�+oY*
������9^��'�<1 ����G=Zo�[����������Tc]w#�63��A�G�����}�uG�7��S#
��-��1�̔2�փ6�l��܂e�\^��[��b*�E���O��y}��!QL�<�Hy5�������ӧn��&�4g�E�8}|�~��2EJ�&�i�'Ϝ�6cߍ��K��_xxi{�v��Fm��m��ӧv6���.䛦ۋU�ا�ݽ�f�ա�N�+��f��o�~vP��	��.-��x��s�l,(D3��7[��|ovj��KOl�����Ӏ<��������B>���w����؅��V��فC"�^iP��>��a��;(	�@C��13���ŷf��N�{��	'0��7n��+8ׅH��V7�ǧ�b��\[A��8]��j=��^j�{�WѲt�[oR�̒{p�2�]��������U`j�q����?zta3�%:V�d��5*q6?���p�I��9�������d7'�7!%���kw/�Q�~_�ӳK�P�*�k׃�����g�<�+������2 ����~sJ�:L���]����~AlE�>�1�n^�W5_���9Y�|q���0�o][�͛o)a���s���z�7��N����2P�X���_�ݿ�%qݎcu���֟���3q����*@A��u���釢��s��'Q@�_ݽ�;�%c ߻�����E�6r�b������𯍈�}G�Po�I� �����80|�J�<�K�[�g�vo����J�R��=oͫ���DP#Ipx��2�����σ����j�Ay�J�s++k_|��o�������i�����vH�z^�tQ����4*I���v�i�8��(��Z"�� F4m�}$mC�D<���k~[M5���S� aĲ@ԉQϾ�u�����|��&{Q�\h)B�@6� �Ʊ��<��sA{pШ��=z�1�7�#�u��n�}��ޭ��aP1
H�`	M��g�1��S ��*39�D2��Rs"[L�yI��o=r��sg���������Rm���͋���}�;q�R���E(
R��R' ��r��Ji�$�rKz7��(��xʥWufV���{��e[���9��+�^������O*T�GZb��t�3�B��	����;�Yz�㏇A�Ѯ�s�ʙ�O<����w<�W�z=���S4g�fC�}X6g�5�:�|�(�@�蒞#g�1��gO>�x�yW�����CS�S����to��:!`h�jE���Bm� 	K,5�	�k��T|D4BkU� |+�H�9� IϾ����]:~�{�?�Q���Ͼw��Ċ�BU&��)ɰ����J��ʹ޵���W�R�v��6|QV]: p��U�H(�?ḮG����m���)�UܰNV�O��F+� :�ئ��ƶ��fmr�g�߿�6*4��ȢC�����Kov�q}UIkVP2�X�b�B�5F.�q�MPq� t � @�UU��F#T��Ia3T����T�q�X;:1w����~��յ�o���=uti���X�h�m�N�C�!��~ ��4�O������,)�
#&�����	--��>=%�4j�!gqZ�ׇ��(��{r�����@EA��"�ra�������7���lH
�po��y��R�H�����Ɉ�~��V�"���,""��$�$�
N^>Q��{p�J���$�p�HɫH�{�\\��^��͛iNݯt��;�j���83=@�� ,|oi)�Н����w��訓ܓ?s�T�^5V���T��H�4R�◫�7ȁ����R;D�됳����CKL��e�*l�Oٍ����{������T%�������:C�UA|�5�1l��W�����Wn5�������%�5m�&[8�[w�V=���'�"��"��f�=�`�����k���K/��-���WUC7�w.�_�Ywi�C�N%�B��Fj�W�+n�����[�Iv{Q�Or:=>k������'s��%��K���x�I�����6��v��/���7$�d�3Q�s3NQM��)	Xr�����ʖ���7��O=��S@���Ն���F��;��"g#B�
�/S S�P�ssg����w��V\7U.`g z㚤���h�j�>��o�|-.�F��}ke����]g��p����چ)�������Ւ�Uń'��u�UTQ���i��N���~Zz,tfXi�8"~�1c���u���8/D!����B};�,�ǭ�L�J��=u��Đ`T��^�r-�q� YqĂ���'�B���	*^�Xb�*�݁�  /����;�1�`����q3?��y���G�(n���`5�K���у���ucG�%�޽t�2O�yk4�Fx�/��W�z��۔��r>�5�8�\-h��9TϙŹ���׾����o��/��9L�&Q�&r<���V�|��� �g�Ԫ�3�9 �����^�g�}2��ҤQ:rt�:�x`���b�+��2��ӥɥ�� q�Nv.�{~�l���^c���O��V"���z}�::�����'������>��:����\\�ѹ׌EK��	FϜ�X�%;A�U�8j�;0��y���S��hy��܍��z�>��h(�����<��|)�g�E"+�2W_����]�>��M츯z�;�w��{�{A�^� N��f�(y����{��T(��L�Dyd���&�����_߅SiI^a���L���G���r�[~|�Ύ��᝘ԖW������ƍ���H�b�軷~�P2�X��F����#ł::1>?3��p�g7��i�p�ч��R����w��N��_z�����bb$7@�%]�'�>|��CՑ�zc Ug�90 �����Bx��v;]k,�����o��<� _<�c������]:9}|~b�`u�w��!A�C5O%���s��}a�Qo���+���/ο�v�'��EM��^���r����ڭ�o������g>�ػ�J��.߼���Ji�_��N����
�1Q�VQ��Sgn\�ٽ_��׾Z�����K���?��3��ޑ�G�j�w�>����=q����}O�q/@P�x� ��uM���n�P��yxBxJ2?v��ur�3Uբ�"�p$��)�Z=15y?l�U�U���ʄ���$2>��dHNRH��<\�o����L�`p���O�z^Q�����:Z�Ҭ������G��ܺ{ʐ$u�>R�H���(��w�3��nw�ڽA/��?@��L�7�7�J7~��W/]��8��WZ��Sf(�1�w?{��C����xeeyc;�y��~E���ǝ^���ݍ����̘���D6�p�4��6��zn�/�9��H"ԎȼV!�z��QW��9f�?�ۼ�e`s�J�Z9��H�dq�♹{梼���Vڎ�p����`���$�2�Wo^?�x:?Zr�<�����(a- $���}�r�����n��}cb$̫]��2X��Q!gNTʞ��~E����'�s��5k�
z�������E!�G��ƅ|�W�_�o��pw� h��[�+�RQm��hf�'J#��]t��*���7�A���^3��{�m�v���:+�j��g�Nkm$a� ��BL
%�MB�l�4C�qF#�^=H�{���b}�^=��8h�!5#Ҍ[��/�ڻ��V>a�<�J��vCI6���@o�J�57H?5x-��o�L�-�������2��^�K��ZR��p0�/���4:?��ч��?X�����(N�v�K+��[[׾���z�F��INV�,��Y׭��xt�n��^~����%��@��ޏ�ŉ�N�+����d����hR	�8e���
��^���L�'Rs��7z��-
��#����B@R��M�杭�$n�kK'�S��{�;���	�l��W�Vݜ��fӲ�E_>ي�?���n�ݸE�jgw��H����A�i�Je;�\���}������"�4��&l�kG��A'���I҃��(*�5�a�k'�� ���ި���Z�l���VPJƔ59Jl%���ܮi�:��W�Ơ���r(�%ܔ|9�(�t;d�f�dɊ��~�t�T���O5f��8a��7�^�M�A�׬�F��b�:�?� �I�Vq�<15��v��a�}5�N"J)Ok��*W���@�N��� a���k7����V2��bx�bXLX�8�OOb�N0d�%	��)�~�~w�F�h� ���;iO�f���ԣ�&d���A��L��w���e���+7�=-�Ty��|dv�������;,�`0@�0$��?f1�}$()ċ��2U���}�G��q�M+���0yՌN���D6@@M��T�9���*�(G�@�8vZ
����P���Е��7�+�ЍzӅs�w����܈�)�
���H	:z�=M�콷�v��Qv]�O�\�NU��(�NG�9����0�`�$�!�琌A9zy��=� �.�u��Ẑ%�#y�"�� �k(����
���*4�|l�0�i�BM��9�+�|O^��X�������]�u[�����M5�;�����~��q^�vnqj��řso���4_Z|��/w�OB�Oe�F"��߼�$a�b�qr~n��r�|RLP5 �	2G�Օ����*1k(����2$�< ���}�)6���4�+�Zh���z�Ğ�¶�N�����W&"*h6(�m��j����_z}���т*
������I��9�x��Y����/���]͗J�V�q �D�y�؟{��#sww7�槞=��嫗ũ�������co����`ӔJ3R���@��
 )�����՛����w�n.�9(2�#���SOO�bQ��ϙ�Z)�'�=�`�)�h�G��?w]��\̦��;4(��'��f�Є/�h8�,b�S�49Y����6��,͍��;7�٪a���V��8d&�Ҥ��=�sY�h��(���1?�O���
il�M.�{��Y{��n�auB>[��F�s�[ ��j)g���'�$,����b
nE1��(�rN?��+/�I}jtnT���]%#n�������b�#t8J��ӡ"H�L L���L�,w���U�<��G{��>�i�_�'ܱTU���|��V{�/�Wr��D���>]HUTbN�jm��N^�z83H�9�Ʌt�Z\��-�S;Q�DK���vgkE4��ӟ|�����/<�)5P^����O�R2mԵ�Y���r���7��-��ؔ����!���SG^���\Z��ׯ� w�P���Lu�ʵ��_�3�o޹\��?�+�����6ae&��2��p�/p ")��ll�lli����m���*�/}������Z=��?����鳕B���G�-�n��lpzanwc�͓�S���+ٙǻ� 2(U,�ַ�~�R,�%�xw{���&�����Sc����vSS��Į�J=�%�0#��{n��s�1�7���2q�����
EXJ��;�����T� ��z�}g�=j�K+Ns����L5�B�*A
��NCڔ$IQI���|Ȓ�b���'}Ź�}K0P�Ҵ�ғ�N��#��l4��/BQ�փ��������UX�@U�*5'�mo�'''GF
i�vt�	5�V�`-��t&��?sF�>������6K��7���3-�ƭk7���X�v�.��#UQ��c�<�������J�|�gn�����4ץ�M]����bTC#�_�~��eBu$\��c���5==�ǤϜ~����mފ# l��}����G+%�O��U� �=��>�n��S�GgN?4=6��ݝ��䘭��h��� ����F1�^�J�*�����/��q'�<U-W	����U�j���t�*�4��Z��
�Πs�'�³)�F�e=��3�#�tt�y.V/]8���-��\0���@g�s���݊�׈2h���vz�e���@�\OԢ��#¤�1����1���A�鍝�4_Z<S-�PW�9��RLy�?P�Cz=����35.���)�k�#S��ݽ���F�y���h�,B)6�߇4�Ŋ!^�q�7sq�����f'�)Q�\��r��ƘIB����ה�;w҂��D)�Ľ�A])���#ܸ�2sb����[
�:��>�!��[N�B��w:����צ>3G��i��	I��������c�=r��Ν}lD ;���L
Qo��p��:qA���dzK2T6#<sxp��ѼSY�p�1�Cțg
pC	��al�o�R��sg��F���f�I��!^�(rZ6DA��6����唑�N�'q����+�@��t �Vp�zqp���o���+#�0ǶԾWb\K|����~��&�V�0�|���^;FL�$����������[��e��WG�"ݧ�v�^��b1U�J)�k�m=��gN�����rC�@}��B�'7���ދ�=��߾�܈�*c8����p���ZF^:M�� �0C�L"y��'K�G�_�|�\��M�������C�� ���;ՍIZ�uw�xp�i+�֑��)�+�ȳ\{m���A�3���	�Vn��XY�*%�U��͍�}t�S_]�4�,���;"L���z��^p�~r�כ+љ�ݢC�?�D��PĔ�T5D��g�pWW^)���r���3 ύT�8���qsij�'��P7���6i� U��r��Ԓ�JAW��Q��B��h��=����qz41�ݔ�DI��sB?�z��<��58��!�Ӝ")I#�a���3g���c��1��$L���y�D���Lk3h�~��Xu��On�]y���ln��~�0ivâ���t��Y��8�tW�7���!w�����RI��L���"�V�k��x�@m�rK���_PN=�i�j�rn�ԣ��P�:]ᕜ�(C�r8�"��|(G��bc(11+�u��$��&E�s�g��W�+;Q��7����(9 (���/�����KLU�$��SV�PU*�ŨjF:ڝ\�o�O/L���u�����۟���޾��k-�͌���G�Yx ��!N�y����m�08��z�62�����%�&%#5�B~�]߭�[���ۇ�uUްFGkz;���z�`se�0��R��]����!��2�j6ke�4����yQ(��ɺ�K�'y��8i����n����&��(d�"����Z%�Y���	�������JB�B��ya1����nQ�d�R�(ڹ�}-~s탷7�U��{�0�#cވ	EL�b����h�Pެ���W/A��h���=$�c��$���VjJ�(Ο�n�}���hͳ��&�o('{�o��v���d5��e��mjH�F�?����p���@o�BJf�g�����Q�Ǝ*��(/�iR��3)��1u(��*����w:^�/d^?���G��l�p�Q)����P}��g!��>M8�)VYTqy<Hb]K7&;��AU���x���.�8k�"ku�}����(хZ?G3ݔdFH�$ӕ��((�~��	�ԧ%�'��1I$	[�/�։�F��A�o�P�L��J�̤h���3"TĩrcC���&	�3��J7��M��V�p�������<��	��#ѡ�����a�4�3?��P	b�U�`�cnv`��E�Z(�뢳��I�ĎJ���`�9C�Ld�c-��`<C��L(�(�;�I��S�k$����G;l*$�0y{�O�c�T�� M`0G�:l7���TgҌ��	a
$g�7�"�~+�����	$���������&��.1n$4�&Ĉ/�v\�J&��&�p�2�E�B+�(c��M��a�H@����B��lc���Y�8�I��p P�TM�0�	����L�I�C��|C���GK�%��@��L�`�b@�D���8\j��ܞjO-�M���]T��=0\"d!�(���+ڬUm��=��6��1�����3���4�$Ox�4!��a�Oh0�w7��o+.sD+�j�p�b�yIT�M�|gl�q�M8���Z	[e�%�bN��i��O����$�II/�j:����Z�y�}���e�@"^�����.��iY�> S�e�H�*����r���V�A�~p��Ł�WCC�št��S�������˗�o�_�M�
I�r�J]9'�l�V��XL�`^aDJ.���H���H	�N�x(�X�E
�$��򀇛-���tJ4���r)ՍS_�qm��<��3?!S�~��8Dh/a�P��D"0Z9������q���.<^�t<��qij�I9-��&�+�9d蒈īe�a��N �� V�رRigQ8����6�L�G�9��K&�1�4݁�b��bOr�� ��8�\owݖ�� 6����=��v>Qh�E����V��w�E%8DqJC[a5f�Qw��C%_)p�o���Q��G+!5b����nO���|#�S��Fb��ȏF�k;!�k��U���M5���ZHa�����V�׉U����w~5=5-#^��TW���t�t�|=�ƙ�JK�$-�A��f�2��ɳ���{�׮]on��I[�#��蔑�5㥉Ź��~��w�O;����؀��r@�h���h�4y��b��~��Ŵ�6oY���4�G�1=��q���'��B��?w�j��I��]��EUce�TJ���=�����ݷn\Z_�_<RZ�j[%5�t�Vr[�x��=�z�.]HW�+'�kD%`h���J��ol๭��1��CE��Kɧù�u�`�B�¤��߯�16=��;o��y��f��^RS
�+��K�{�0*���������?hS����t��G�w?���?�y侊��G/����/���r]S����
U�~��s���M��sW��o�/�i^��ю��\G��C�����vP��w����ϼ��9�ZG9GX���X|���?,�*pD>����O��[+��Rn/D����P؋�}�����P���v��?�_��[�#'Ǎ�j*�A��wo[�#��ȑt�*�M�* �V/���c��xe����^�g,i�GZ[���s�񼗴­{�Ϝ}���������~���޿ri��~� �ՠbɏ}��_VUK`���?��g?u{���7R�"A��*3'��W��u�.yiq�Ǟ�§_�W?��鉰�I����7l�Jo�#K�w�;��]�wX�.o
�|�_/�&<E@_|��?��7��_�k� Q
B]Y7��������Qա�����+�����v��3r���X�
�p�0N�%�E�S#�m�DpY��sO������f9���k�ԇ6%�	3�Z��yV��~���V���)2�N��*:�<3��z�b���
�V0H���&''���	j(8�BKj>���E�8�㓓q�ÐOl}�r##�@�A�i:�0�z	������҂f��%i6�h!tnfV��h@!���Tiq3!Yx�XX,|�)��i���ma(�l�'g��b�
I���Z��#`V�h<�Oθ�AA7(�h%��]kjꑨ��׊���F䅪iI��w^�;$& �}Mu4����A���*�Ke�[�I�h�bg���A��+V��+�_P���:�^~��H��n�����C��P;����(�\�A�	'B�Z���߯��˲K�����;�8
sz�;����^�~��/�`wM����il���A:�̋
�fFE5��Y��k� � ��a��b!�W�tal�\sB-�<�������-$�LX�te<��q�Ə_��~�˚��"����Mjh�UN�L��
E��?��~�����;���߼J�Fy5Ԃ�uL�{�����\!i�¹�?��+���"Չ��M��?�����R.U�X\�t�?��*G���rCxfI��O������5�5��秿���4�U`���V�Sa����w����d�<R��u��׾�}6]�O���y+�3�N�t�C�〝�v�T�Nɰf�T��?�ko���|W���Wƫ�ɠs+���a��rz_������s�`^�;�����.�� �������7�����;s��F������yǄ��jN�A{�Tz���[7/�XX8�ٻ�v/5X�F�դu�Vܭ�L�u���?�o��,���[��;X�6-Oऱ؊ڵ���n_����W�>�d�q���"	ʁ���*�w�S����o�����Otڝۻ�k~}pv�~Y9��Ny2��� @��8�Z�]�:њ�L�q�sOp�i8w�+s�`�\_ul��n%�>��(x��W��-�ZC���N�9�����������ε��q���Z�>�#� �r�틫��cc�v���a��S`]��tX(xxM%��;>��
��O|?�����kŊ�t��v�^��GKq'����ݞC��#�̴�q_��+ۧ)�u�﮼�6Z�/L��"�9�h\�bs
�Y��.��ȸ'�Ȑ�� @eU	��N�Jb������P���Z�T:��?Ƒ��l�",c��k����La���(��@Um�0]q�*"G�%Ft8���UU��+��j���}D<�H�N����ZlO���ΦQ2��COʸD�n��h킽I=W�f�-R��y%^�e���YP�O���q�:��k�V5�p��Y��F9�*.�LD%�Q�ZQ5MΌ�j8��7�H�6����@�R��1�V���`wb��jy%y���8�[��$#��A��M�|��l��$+0#���!ZJ�î�[6�1"�H�&*Vi�ؕ�-y���n���Ƣ@x�S�˾���;HC�R��C	*���D�S��AU�I�E}�D�ɱѫ���T��(�a�J��g�T�����GB�.UT��T!�f#�Y�	HN�"*�h�VN��А'�5����~3��~ttjmwm��SJ�K?���m#�&B�ӹIU�^��RHm��X����CqL=>;�����}H9��?B��YI%�^\zr���ӱQ^L�u|L��s*o��9C�H���c��w���2dmm�α4���Kw�o��p���ؙ����?��G���dÞ�m8J�!�C6ӕL�CNS�L���XK}Q��%$�ĘY�Fz�-7��;0�j�)04�-3�a�[�4!��Mj�J�Ql��Y���N_��iCЎ!��B���Ze���!ى 7��nr�$�9"�cdr���D�����^�t<S��ڍ�<T��k�
 >���k�C_Mc�Lj6>��N��e��rUP{qx���x�M�J^O�c5��5�'5dź�̏���5Z>5�T����n*F*�����?$ǂ�Y�r�
OB�XR�*F
��FV$����0!㎎�'�r�D)�F�Y���!B֡��V��B��p�j�%U2Bu�	#+�s�*��N�f35���I��p��"Jj�c�O�Pr�(�ζ��d3I$S���l��F����	��TeA���N9�G*���i�}Y��MlA��<�NG�=���f�xdO�F��ag%r��!�R��|e�H��S���?hvܾ�`�7��{�QA6�)��Lge����~�I�z)1�6	�p����v��gf�.��]�w]�H�@/Z��A+*ŹȰ�"��h��\9d6�ZR�F��/I�|��}��lΨ�eba�v���|׃���+�<DYt�˹�>���f!lP�,M�oy�q��K��xЃ��$�Zk;��$L���(r=�b6xW$��{-����zdF:B�oL��QG�k̃,��##�w���=�%x5��r��D7R��ۑ/�k���8��)�}���Tf*�J�ʃ�"�/)R��yy\���B�I�}�<w�2��������Ϟ��W7�ֹk�4]E�8��&Ot��o���X82ek���u�4S=��(�r�����5Z�Չ��ܦPo�(�qc�v &��\����&˿ھ�?pb��4��gG�I�Zg���<�L��q��#'���m�1���������B�`��:>1�S������PȌ���������)�E*mqb�æ����dnY����"�U2PxQ/F[�E^��cgcgzv����ܕ��LD���H�4�	�[<;��vVȄ�4=JJ	t��?U�{&�Zi(vv���n�	�0aH
cj����Ǖ1m@%�����z��GI1/!#��Z� 8��~���w����t��~GW�"��)�������Nc�vdBC)4��L5�"Jg�2q:�"A�(h�Rl�+���"9�"��4��1Zi	>@#a��(D_�`՛(6ס��$�!H�(��22:Bu�5>1��dGoQ% �WZ���\F���u��Hഩb#�e���sl�F(�.)*���bh�0o��ؘn��S��ml{-��"
���1-bU�@#dm:���xM��B�j�����W����|��*&H9���371z(S|ȏ��^p4U�Y~�V�q"�ӣi�Gm$����3��';>��}�i�$S����9*`ʖ�jv�V���Ś�s�^�����$x��r5���Z�8W{�JR�h�P�C�P�Ŝ�Z�]g�+]#n �>0h�7*�3�v;�$�Jv���}�ld)��Lh[
��Fd����,sSVh6��2�F�^��U%����A������j�����T��J]C��x_&5�I_�}y���~�M�XǬ�*�u5F7�Ƞ��4�9,��g�%�T�BGV%� m������'G�&.2�J�4����r0��@Y%�hY����o�1��`��<�а�]%@�'\@Ù�������%���4�<��!(dh���搽���A��.�˃=�#N	7����`/����R�)� Mx:�0�C�j�B�@S���!S>s��ӎ9�!�2Rp�7T,	
^�#[jTW���'���rVd�m2k��d��,�3� �%H5./9a/4'�1R���J���@)�'� �[�3����1)^�(�e��th�+2����'=����
� �aC'<t�J�7a��%�̖]�ɗ�T}�~E��"Iɾ��DNE���gR�
�n�Ć�K�L�_��x��dJ�ٸg6J����m�b%k�a-�c��P33%�P	9p%+����`ͤ� ��R��#+¤���e�1���E�Pd���M�.G��B}���2p�D�)�����ө ��n(F2s��"�ʙX�g4�k3=�,��?�l;��@�Xoƶ'���	�ETe�f
��i��]F�R�Mj(YI��쐲�	�#g��b�ѿ�
��8�en*�C�	7<��tO�p�ま�9$�5���K�@Y�� .������������まJ�ǘ�ʡ�����i�+�2z? .}$�0��$CQ�CO����syԔ��dV���P�\u�����G�    IEND�B`�PK
     uK\�$<�ʏ  ʏ  /   images/cb669bd1-12cf-42eb-9243-39a8a80a0435.png�PNG

   IHDR  �  �   Ͱ��   	pHYs  �  ��+  �|IDATx����w$�y���{b��E�"Y\��&R�6S�%�ݞ�̙>3g~�n��3�m����m٭͢eӢ6��L�E�,�U(�	 s�'3/�L�2�@F���9qH�P���'nܥ   �"�  `��   �)(   f� 
  ��"�  `��   �)(   f� 
  ��"�  `��   �)(   f� 
  ��"�  `��   �)(   f� 
�0Ց��`��n�i�����R��+c�mOK���V*��j�ک�j�7n�����ϻ�ȣZ���j�����^���5��x���<��=;��v���΁c�w�G�}�< J� 
 iɖ�-sZ�ƒ�g��<e˒����noo�� �`�kÂeU�����A�k?�_v���l�Z��Vx���������^���jo�~3
g}������n>��X�1o��J�^_��@��r��o��5;�k:�wk�~�$��{����;������u󻻻گ���������u�n�Ɀk�z 
� 
��juZ��m�͖���m�����
^P+�-<.Zٶ����j@��כV�����Rg}(�*|*����KKK;�㎕�Z��ol��U��Za�f�k��n������m��-���-�A8���Q��ypƖ��E_�o�t(p���W��v���9�l�pێ�f<�#�'v<��:�766t�gC?PM��N����jG�������-�myǖ�my/��
��( (P��i��ϟ���6+/Y�w�
�����gmm�0(|�O�"fP����k8�w��-���������տQ娖�7�߱��膭�[��i�O����-���X������t\���;m�d7Iw�q��}�@<P�fÎ��M��t�e��c��NH���7o���+a���sJ�y���1�a�={�-����7��^���aNT9�(��������{�B�cV�=h��V���n�U���m����0�d�T�|?~����$��߷�7�3�yZ����m�������i��3[~h��l�`���7TSD�(&�l��)r��}��-��rA�@��X���M�^cPL�(��_�q7a
���A�3J��=�T�j/m�g���S�ǇmG߷sE��?�����������Ϻ!��3P��*.\P��e+螰�y{啕�����;m�#��PkyF%؃�h!:�da>�����2o�����C>a��-[^����}�W�s�����G�� �LMM��W�S��v=e�;^�ckŎ��n��z+񸍿{�S�� z��w�Cn�~6g����+��������|x������b��U��7�f�g���p� 
��+��B򉕕�g��777�B����[7>�r���}�ߙ����͂g�0��n�{�-(��B�a+�_�u�G�߲��k?{�>�:v���#g���.�1�H�^�^��cD!�^;f����[ǘ�z�����Z���G�w�qպŠ�s@__�~}�n/�:u��\O��?�������i��{�s��
@�@��hZ�\�B�=b������Vpޫ�Vϩ�U��F����P���-Z4�>�0ik?����}��^[��~H�����W-@�V�[�;���g{݂�7�w�a��pD�X�6r�hiqq�Ni�ڱ��Oڱ��#�T���s ����s�?<��\ͿΥn���=18�k;��O%��΃���ֹ�����혿�>��vv����3�r�����?����� ���+pϩ#�LOX��T�[���}��Uu&���Tت��!T���;�y,9�����M�&�R��q� ����z�/Y�|���҃��s߶Ϣ�q?�\7n�P�,/��cv<k����;6.޸q�ܨ�Il��ck�3ܤF;%�?���*t&��;y>�sA��>�[�9�w�5�{}�~�k׮�f7i߱�����	@�@�Ν;�d��=V�]�V�>���~�իW����;��Qa����+��L�H�qgښͣ���l��Cs\w}�R�w޹d�{���?ۿ�����_ڿ�g+���&G8k��1h�������'��s�h��~�������8���aA6y�����,~�lC�^�9���(����j@����s�s���h���sssf���~�A r� 
��8s���V�<j��z�
�� �x�M=�S�d��Xx�Њ����{��O��縎H��M�����%��>S˶�ŕ��j�h��ɟ���t����|�M����:�qp������;�9�^�٩c9�67�v
���L���U��ף�5�ɛ�h8�&)kZ���}}g��֓�?�s�ڇ"O��3����-`�ge�3V���B���~�3��M��kǙ,<GkG����~7�4��K6�mQ�����wضx�ڵk����M��'����������s�;^���z�޻+�X%�}�>�i��$��u�����:`�e7a���B#^�c��A��7��j���{��Y�"�>T����XA{�
�ǭ�U�'���,P���gr��X�s��ˬ�O#�~U!�w�	|���m�����ﷂX�f��B�������ԞB�5Z^Q��p�͗:�=aA�ۯ�666�y���:_oU{öjJ����[�t�ۢv�����U;��kג��y�0����z�9(�M+8�B�,?977�����=V��n�s��R����c��~t�71���>�T{�s�Eۆ�YX������h�߇��tT�7�g�JO���u{}���%;/Vl?/��,��w6*�q5����͵����f좝#�[}˶�w��_��[�Q��� ��vZ5�V���_j�Z��j���X�F�W�佶�$${4G�ġNX�.�����s�5����q:F����Y1if�Gl��-����)3���ڿ�H!�p�v���Q�n���5 ݤ�a;��<Ԗv-��&F���-߳��J�(�SKKKg�@}�
����Q��x�ڵk��<��=~_� :8<�����'*�&f�ѳ�%+��`_�V(�����5O-P�hzLM��[�|ޖG�^r<�䴗q�X�lҙ��N�B�(�~1��f_���Ն�[.����~�[�\�@�Z\\�M=۫��_XXx�
�q�_��B6>nO�xP�<�&Ho(�&�S�����q~{Ֆ�̹�d����;��P��`����e��Ӫ�����0??�΁��b��W�:��f�9ړ�KkD��$�!1R0�sDO� ߶m�g�뺽~�~|# '� 
�j>��x�
�g��@�7#3n��X��1S�����#>In��@�
9W,��ODw��];?ԄfJ#=��cvL���o����o���<�c[��ԕ�!�0p�PQ#7c���?o7k��rm��f/�8AP G.^����5�̗-�l��7nT��?�t�j�0��B�-����GWVVv� ޴m��kkk?	��,hV���v�_���e;���}��}gz��x8�|Ͷ����o�ұm������0��8P �gϞ��^�� ��*x�^����J||���M=6ɶ����i4������S���ڵk?�Й�s��Ϸ��/���,|^� Ԉ��etlۃ^���U;i}m۹j��i���v�///��m�1�<N
�^�
�˭V�%���IA���_��(��GQ�M��0>�]]]mY���������گ}��ůN����f�y���o�q�)5=Qw���K��I��@�C�~s��bס+�ƾ�͎�?�/�e��]�'�8FP [�s��=��V|qmm텫W����ĎzT�B� �G��b��j�Z�f�I�g��}{{�����oZ �0MtN:�ja��%[>g��%�+�yܓS�F�
�j��;h*��ׯ�������g5x�]�n�s��Q"�86P #KKK�좮�ѿb��[��Ʀ�K���v�7��a�/a��F��p �;m_���vww�4�߷� ���8N��:�\��&\��V��V�`\m���?������iv\�)9t��{
�v3|�n�^���k�F�_�^Z��c@ �q�ƍ��0K����>��ih����LS�>omܼ�z,iaS�����V�����x��k�zB�Ǌ-����m�t��z�+�Zi9�q{���p�Of�Mk=�΃����ö?��b�k�|ۖ� L� 
̞λ+���V���������9��/f'N��Z�[�{�~���A��?
���]� �_��7��X�L4����Zj�\���k���D�n�w횥PՄv0(0[:�4������Z��o붰��/H���N�GTAT��~�`���}��i�)�Ài���-_�岶�zc+�4ne����M��G���}s��ї�y��њ��s��kqdP`����q[^��y�z�&�V-�k�B���U}kk뱵��O[�]�O�	�S�ќ����n�^l6�W,�4��}����v4�[ ��yp��3������������Yx�d�g�"����XӠ���������Iv�P�l�ۚ�'|��s�V������%�3Isb>g�Onnn6U�c?ִ!;�F ���2�Y��~���F+�[�82(0��i!�Y�p��aPT����LB��Vr�+Q�a;�ʩS�40�f���}��k&`b+++w���=?k�S/T�n�G{7�Tl�1�ܮ]v?���}��]�~j���8(0.\��#\�h��z�B��ੋ�
�x�'|���#ȸ�t��l6_��tuss�����t�Ѱc�z�);�_������k��J���d���I4�Y��<��]�^� ����GjP��Y�\���Sv���-���y!�x&y>�M��������N�z���;�Z�õ�5��'A¶�)�~
�_�s��T��0=�%���l����n�K/ھ{ceee��M[KE*P�d�VWW���WC�����,��G�&|N�(!f�����j�z�~+x�����o�����t��>��+8_��ܼGcJ���O�i�h��j�z�ٳg�datuaaa�^u#�	�����i-..>h���Ɨ��}�.�u��]k��In�����ڵkU���>�����??��^��v��m;M��݀UԞP�lzB��?]�t���-�پ����ص���x#0]'&D N�������]������*x�c��`�ȷ8$�§^�(�n&t����߶B�]��[n$���'���v<����Vz���F+�4vHz��v����ӝN��>77����o`P����߱���I�(��3g�<g�m�q`��Գ2��ƶ�[[[�C�g䙷�Oد������\�Ѣ�'5���>��Mu������6LN�y��ae9��p}Hnk�x�����[z�c7��T�����&@ ���~Bc��ͽh�mC��8z!�$�
�߽Bq�,W���677�9fIz#�i��v�VÎ�q��}4�f�G�q�kV�zx3Ѷ����s��_��蘇[ �ǫf�%�8��n�����h�w
�b������}Vfcc�a�(�z(���<�m�h4�Q����@ƍ:l�~����v#�O��/� n� 
�%+h�XA��]�/{������C�����S�&���Oپ֣���M[��K�[>i����}�j;��hMZ�M�Oj*���^�勶�i��(C3�@P����^���/����.��y����/v���>V?go}=�;��m�s�=���r&��s ����B�<�4KX����S�z�y��}�~��0�!�"���]�<?m�;ua����_�l����L��4u������b_��A�f!j�^�s���d����pN��]�=�ڃ�Z-�_��^��y;� 
���d�gmy�
Z}h�ݼ��h�M���HC�
i_��c��\��1[�	���e���-�f��Sv�u&v�S�T8����gj�2�G͵q�$�T�������	[>��锇����X���i ����8�q����p>%>R�>����V������3���~�n(5�˖g���.mllT��s�qo9/|�\"�pGj�n��v{�v��vԂ�C ����b�����C
�*xU�Ʊ�P\���ߧO������I+��c߿�3͊-�U�U���vyy��E�D5��qmlJ�,.����M����E F@��5/���v:�sz#�|6�L�����Z��!�P�I������g� ������P|j{�΃��<��>=���M�~V�+��)����kᓶ��� 
LO/�?��^T�*��ځR�S\�5
[���e��=�v�i�Z� �@k��o��f�y>ހ��qP�aS���|��9���;��|�}�c[V�@ �SYZZ:oꃶ��#�豣$k}�*m����&kXc�WQ�CRH�����PԂ�bSY����c�T������0���f,�o�6tܓ��Ά������nڳR�zaa�6�	yľ�F �b�N����m��3g�ܮ �}���5Ay5�ƅ�dM�>S��jrZу�~��V�����j¢8<Ϩ^�GPI���9�/�	��
����y5��E}�l�C��h��B�Y�Ǩ�\HlJ��t(p���$$�7F�/J���9h�If��y�l6o�ϩ���H ��i��������
�j,pT0��ǌ�K���F�O��A�R��׋�[ I]w�<{�\��~̂����߲������{�����FlQo$���J2��c��xl�M����*y���y�����w�L�î�5��������	�	�(0� �d_���QI��y�d�,Tb MN'�l�kE�������k�ױ�3�����:-�|�VKӱ����m��>f�E[��$�_�7�Bb�}�gυx<'?y|ǧ j�GH�?�$������9pޮ���v8�E8��]`o���aw�3�*p�Aa\pР��P1|_U����e�������JWm]_��}i���y4b@3SF���R`�0r�}�ǭ��}_� j���v�<���tg��	�9���s4Hύ�+J�j�}͖M��XU�%X���x������),���.Z5�K������~Ǿ�@ �Gv�ܹ������ �G�'ۆ%_�n\��H�LϾ�Z�۳e�
]�m�3[��[l�ڢ�X�ۨ ��m˼-˶�f�㶍��N�{g�Kv����-`�h}&�����{�>��쭟��	�b��^{ՐS���YÙ�����t:�VWW�����0��GM,�y�@��U;=>P�\�`z������m��8e�}łhugg�j���ԙ;�ٵ�f����t��@ �Gf��JW�p�3�zk{��9�ӻ�U����VH�m���Ӣ�W��U�6T@<Y���:\��ځ���e�{�/ZV�X�>[.ض<5IǦ�9lv�~-�,St���Pگ��xؖ;�|h$�=�� �v^;ulj�)`jV+�u}�����k<VV�F��p�9�P��v�-wix"[�@��w�-�m��nX�FۚzoDT�kA��mǇ���F�G �F�����Q[����1��d���C�r�n�+aP��/����z��l�[�7�?�MՊ�vT5CgmQ��˝N�����wi.�d{��8l������� �,4��������������:�%�Ǜ/��HX��憎���[��h$���rc�?>��3����0�f)z4�3�a8s�e=HNp���)��jm_�>�?�A�/��d� 8=:S�����ow���X���Bb�
�7��?���ly-�WI���>\D��?
�B�1�Ѷ�@�l�[�ۦ�)�>����vB14-0=`AC��s�G��$C���uW`���K�lko�a�{�W�x�.�s@7$���i����m��h@�x#��§��K���O���?��������J� 
���?�6��r{|������R�k��)��-��p���B�U�f������7�p<�����]V�kǊBF!h�պhI�_��>	�tN���X�vCy���z�_�����{�ꤦ������/�r:8�����ب��m5�y̎���AM���'� 
�W���j'�,,,��i�üH3�����
�o�A �n<f���S��c[.�r��I��y�Ұ�'~�f�Z!|�ο����>�:�,--�GK��~�6GN �� �x��0���`y;��,��U�� i�۟�5�=y������V>sÿ�_zP =��rwlO_�?l�J����c�,��)��Ж����l˙�Tl]�Z�����P�6�E��0v�j�,`�%'&�>Ea����O�T�2|&���j	�.T�·���c���L][[���:'��u�T[h�@��N��]��Ǫ�^�q:�D���^�a��S5�[!;z<���9['��9[�Fg��ptl�t8-c�
��vâ�A`�,�e�seث���U=��d�}ߌ;L�>�9�W�坐m@ux�K[���e;�F�zͻx�k�{m�s��z��N�̊TrP =��VMV[!#�c;�Ѓ�������H�����Om��à�z�4��߄� �Z>cK5��գ���f�x<>,|j<H��|6�z�;vT3���K���7�Iρ�������q���VN�Q�6W���������A���ÑV����iK˶է�U3k��wt���H��'m���ZG�z�)�p���v��<�����1 �)Y��h];S�8f��c%�c�8�z���a0�R^h�'�ƪ��L�Ѹb�Z7�v^%k�����/Xa�-ݼ��RQ�;�X�&����CS�؏�6U+��0�ϼt�x��Y�=[��j�%r�^�9��5M;��k�J@�@�t�v1=eѳ
��0S�J����a����jU���`��<������AgQ��%�������
�8p�����}�M��7z=?m>�5�6��]Ì)|�'o�i���Eþ-ۢ�\tJ:�f����������H�������EDz���m��"��l�k�˲P���*x��HX�B��-�E��LlÚ�v��X����[F�vh�!�^��b�>�����(7��a�HC.�a���#d�K��˝v���E-h��;n�_��M�	�4�z@i@�tZ���^o�׊ǹ�U0X�Ta�����,o�>Iz�=[��������o�Zg���SうA�aPu�Ȳ��4�@[�k��T�s��};����Ga8m�'m\�Я��-�a0��K��m����F@�@�t4}�]�ͩ�W�0&�6/'�I�'*p@U��i��NA������KKKw�Yw�6��8Z�� ��V�S5@
^�Bt#@��7)�F�����P�S�����H���e��b�V{:�4$=_7 :~T�K -9(�B��<��t�P;P}���I�,�������Y�k�Ϩ_�AP��m?=�V��}���>��#���B�I�A��� 63H%vR�15���U�g�j��n�A���Q��BkZ׳q��� yg�J�g���n/nmm�PZP ��+�(�V�ߧ�ʲ���[�.T�6�W���j����q��wT<�O�uմ�����'u�Q�jq[1��F �]��f�nh4ެjA�ݘ�#zR��y߳����z��gUmY���kx������唅�v@�@�tt���/�<�O"�9�-�i����l�'�����Z���瘛����DՀ�X�z�ɴt���_�;��4#���9�Ьf;:*͡�sW�!;���S��ENhl�#��#�)X�[�װ����9�o�,����W-ʛ�\��C�
ߏ=2�8i�ǎv�hp}�>M�LTZC폩���8R��%I��Չpwkk��}� ��c?y�;�|3���@
v��Y��߹�=�uׅ?�zȿ9��/*x=��R��j���틐c���&D��
���OЇң�v�����G��M�j?]����Հ�;�&8��ݰٌ�!u�$��H���z�6�":qx�����k�޶(���^�R�����kv#�b6�ѠfǏj�րj��eGr8����ZO=�|Ҵ�W������15�I=&!Y�O+���@
;;;z|��J�Q(9Ϻ����>U��5�*<�6�N,t�<&hr��D��j@�	�k���Zr�V���G��^��j�ooo+�zk��WS���n6����3�y�Y�dd�4e���R#������.������^>k���Upyl�&J�
�]cO&��DHV�c�{���:+QT�d�k��{vު��[�$5E�B�;�����k�n�td4� 
LN�V���&�^J־��#�"����h�vm���z<�Ф�� �g�?N�^�T|~E!�+DZ��;����Ӏ��R"���4ӘǪ7��^/�7�*�<��Z��6�Aa���Խ$oNF��gz�i�s|���������~ �r0f=+�%E &׿`�A���������w��
`�*����z��{=���1�cB &UƵsB�����z�?�WE��*��sS��v��S����䪚FN���V �� �/�� 8[�)��~�s�;��"��@���k@���#���U�u�3��90H���}�M
�|b���@�tX��y��!�����>�r�ؤ9�����J8AP`
=�'����y�������Q�"�GD�gf(�0�C�y�Fw�q�@��U��wߤ��9����͊��Y��J�v�p� 
LnDz�g�(�&E��h�P� 
�F RЀ�N��<����}����"��8"(P.\�QvE9\|����h��bzP�z<v<�~nj���v���|���qL�������^���0������yW�"��_�������p�/�g8��!��}J���2�� 
��^�y/���?Pv�/�8P �>1-���B ����*�g ʌ��   �)(0�J�_��}� @ &��V�v�8��j��T�@@��)xV5��g�O �@J�j����#@���H��'>��ϵ.�A9@ ��G��(+�|�F �ᢏ��q���T�l����A R(�E�Ǐ7Ѧ�9`Jޏ��H��+[Ǽ�	��U��E�dE�� P<�)~
��@��Qh�ߎ���y�#���H��0�v�=��t H� ���]Z� �G &׿��z=[������,Ph(���1S.��A �n>?
�@�~� ��Px�Z�&���H��"|d��D���
�B &wӴ9̡�) f���Hg��i��D8��@  0SP �-j� �H�����f ���<�8�^�R��"��lU�o�z�#g8v�G �٢ PzP %s��_ N�\Qj���9��7Տ �#��R��	 �(�R�Z%�e������?��@ ҡ�Ei����7n �(��-{8*�L� 
�K�QcQ@QV$h cP   ��7�^�sP  |�&�@��q�80=�!@���p�q9@ ��e��B
�( �)([l cP   �  ��h@ ��y\J�Gʌ& �S!F Ȇ��K,()(   f� 
�/�u@��tP P ~�!�� �)1�u�h3��� �H��	�J��'�1�1( �l����#���ך�z�]  L� 
  ��"��+R��N   #P %z��ԊtC�# �  `����� C��i@��� J�$�"L� 
 H�u�(��r~j�H�B/$������(   f� 
�O� � sP @��[��0@@  0SP�|��� @�@xCx ����>  (0�J�Z  `:P @��4�   3E R�v��+�\���(5( o����}��ׯ��ժ���1sy�"o� 0{n�o� >q���z�O� �   3E  ��"t�C�@��q����P��PbP �P�bZE9���{_L� 
L�(PZ��1�P`r�AC� ����a�  S"���u������Q�5(�Nn��V�L!Թ�G�p��;�J��W�窦 �V����c�� 
�@%��/���� r� 
 (4�P 
�� �F ��}z�eP y�	(   f� 
  f��SL� 
 (P�x( �<�E+W�%F ���j� �   3E   �����#�  `�� �T��`ZP @*�D`ZP �P���Ԁ�� �wP�\����T����@J���g�����u� d� 
��|&��@1pH�BL�ce��&Ǆ 
 �G�2�P @*�ó��
� 
 ����#cU��v��^���� 0{�k�<�{Q�����lZ ��-0��M�Ps��2F �[ �܄�`jP �A��gz�^7p��(�"<B�Pͨ�-\�J� 
��Ee��s����gP �C�O�؁%G  �Ap 05( ̞���G� <#� ����ȳ��gA��<�ZTrP Ϩk    3E Pb�%	�x|��@JP�O �H��� p� 
�P�V  �H���  0(   f� 
��#x  �G ҡ�  S"�  `��   �)(0���7c @zP���Oڱ 2E  �����#PP�X�`�׫T\gPNR ����\C�N����( o� !(5(�R���G  �F �!|�쨽��!�G R`.x 9�M �#�  `��@��� �9(   f� 
  ��"� �Mi�(
/���^���_��0(  �p#	���G*z�? ʊ�	���G�O �cP   �  _z�� p� 
 �/��h��   3E R�v�  L� 
 H��_ �A  �I��3��� �4?8�D$���#� ���#�ROV��W�}��2(��A  xt�pU����c���XI�(�L�� ��@  0SP %f�  `:P`r��Y1�g�D#��#x��!���@��q���o�=�;�	H�6���
/@<_�<�;�	 0���>~� ���yAG��هO 9A �N�Z%� �cP   ��k��~a �H���#�	�#*�y�3�t�F �V�Ԁ��A�@x�_�I �)��pk!%G R�v�ٳ�Y��{�- ��7�� ; i!��L�%�1( �b (R*B�\#�p+9!tf�� �F ʥ05?�����(P>��?�P ���\W=3d�P �^��������P  |q}  P<���Y�@��q=���d��Lq\� �Ҡt:l=(����pdԀ�@ �	GF(�P�\(}�b�\�kP �P�f��`jP   �  _���{P �n�[��8��? �9(09���0�@  d$�yuH�@@ ��O2��PrP �Ph@@�t@�o<�r� 
�n���05( wzL�r���{P   �H�{����X��񕠙� H� 
����>�( �)9l�ag� 
��Ep�p�3
�aP>P �}��/|��L� fk+ � f��u����`_�5�B GC���J��2��GP>�@ �Y��/x0�� xG ����o �F ҡ�������� 0{� J� 
����������;� ��~cJP �Ph�p� 
 (�j�J�3�P`r�8  p���9�q�fe��P .�E��	��Q�ղ�yT7�P -�~��g�{�s�yݑ=j@�G P2�(�r�@�E f�@�@���@Vx�>( ���;9Q (5( �"f^���(  �"DkB(�1(  ���1( �t�P���}P �=υp�� f�s�#�� ���� '�@�P� �(j����&���	(P> @��@�P�=���M$�#��C�������A�@�to(3����( O*��5���p� 
��<�ZTrP �h�#jс ��G�U1�����: �� 0( ���� @�@x�����A�%(P>ġ��Ky�'�\#�����o�  �F�NH�c�=(   f� 
�j0-�! cP   ��\z^P� ��\Q�[Q>Pf��p� 
  ��"�)1M��8���!��3x_(�N���p��S_s��Dt� ��@:�g��W  ��eP�������'{� �F ����Y���ynڣ�*�P Bq$�
��P`r��jP �H�@@�r��8��@`�?3����܅�P(( o(|1! �� ��o�]	$S sP @	��((P>��  2E  ���@ �	 �#��Ј,[�O ( (��� �}���g2�< 2F ҡeGx05( �!@�@ �����H���� �)@  0SP @iT�>/x�TrP   �   3E   �L@`�h���� �4�8t+9(��oT�����^p������Ռki�@ (�2F   �L@`��PjP`&�op�0���=(0�  DP  0k�QrP @iTL@�X��� �� (x�����"� �"D�
 f�{.� �F ʇ�+#EJ��^/МSb|�#�����U����k %�υ@;��"� &��P��YI�P %��A  ������<!��H�����@�@��Q!�f�tHA(����۫�h�QzP�pJ>K�Q�H� �� \"��K���Vg�z[�����	"|b:R����GP(���8������k(�@
��W�(������L\�QP`r���SL���rs8��/9(  ��J ���;�� �S�ժv��z�^-���@�� d�2d��-5( o�h��G�8�@  L���p<�Y���N-9(  �C��=F����{��7|�c��� �T*���Yx�| ��l�d��9=B �	`*L	�   3E   �L@��hC �� ���A*�M��v�̂�� 
 �T��㑌*���^��7��a>�P  �>oFh�@���^py_d�{���R�π)@xD�"|� 
��(u���8�� P6���QZrP   �   3E ���ǧ��Hm��*��A �J��V�� 32�yj�A��� 0[�l��g$>	�()(  �"$	B(�1( o�!�(
��PfE���� �4� �F &6o�F �D���`Fn�%F &F��.�!��	� �)��� �wP�\��{�J���U ��;�n7 ���Y{���]y��~�E� p"�ٓ�Y($F(P8T9�Ĺ�!Ԟ�@ 
����� �V�@�� <�	���8:j@s�8�K� 
����V@֪�����h|�8"A�A�Oj@�| � &��Y�v�K�'��lݩ}r� 
 ��M�M5��Qt4&���� 
 H%�v����� 0{�k�5��6���[�b� �yz�ZQ�4��p� 
��E���I0�"tB*�u��~��@J�9
-L�(�Ϳ3�|PRP =
0�Y�y�#n`��YjP 8!�s�^u���;��$;��tT� H���\�T*�r8Bf� 
�S�0�!pEΊ�c��5(���;�dP	;.����Q��n�
4g>J� 
�����Z����ʫ́��?�D ��~����}�~�$��H�R
�F &W�Zq�,|��3�d3�&9��?F@`T ���1B��#�bH�u\TpH������}�q�@:އa*J3�DQ�>�Q|P �X�:
��L�r˟��T�(9( �^���x���8x_�9�8�J� 
Tl*��t.hT
�	)v�rt��YQ���@	$z`S���h(	���2ٳ�Y��w2(7(PP1t��"վI:R�Nj��%;'�������oV�ρ#"�k�b�,� �UD_�V���n�P�g�n��c�M�O�"��ׯgAl]�{{{��WÖjЌ��Z��⹹!���@A���&*xzvvvr;�{2|�}1\�n���W���e��������]�@��� 
�K��5�^��4�bMЊ����@~w+<�jѻ����G�3P`r��m\�[�
�J�����f��/|����4�F��H�����NMM ��OaT����~b�A ݫ�빾���}�)@�t�^�����0��5�ɰV)@h�� 5�^�,xv-xv����
� 
���j�"<�W��U폗 :�{/~W� ���tuܫ��c �}t��X�@����G�hG/�y�]4sss;�v�{_��=�K#��N.�LOy����� F;����+Z�R#���Y���]>:�N�CPj@c����� ��31���O.*z��0���e!SL9�w7j@ˌ 
�d{.����lܸq�?�L���������+nv?�T�kAojƑՍ�Q��Ę�ޏ!L� 
Ln���^�p���а�YS�_О�r� 3��t$χq�"mǬ���y��HA��T�n������f�������5�������Ji��b�U�_��"4A���FxC &���X���^C�v�@���Y`�jt �䏂�xv<?>��]��"�v��#�Z[[�z�f���?v|�ۜ�Z�8M��Z�p������{��f��y�ƍ����w�qǦ
ޫW��������k��d�f��bUs�j?زm���8XR8w�\϶���ӧWO�:u��w����7�Q�<'F�&ǎ����f'�ձ�О]��4�S�f@�4�IM�ߓ�3o�3J��h4T�n-,,����y.|5�RgnnnW����ځ&?k^J�dh�{��Yl�S�̎����R������P�E���u��+��@����5Q��V���j��ׯ_^����?���ǐv�geG���¿�#sq��c�j����=�:�F�<!�����0|���vUK|�C���0l���2���9��z12n�ʽF�nǽ���y�+&��?P %�g�,�ն�����Sc��=�1A���w8��@�nQ �ZЛ�/ףa3�����	�'!���E��z|�����QxP���Z��{��2�xh���a8R2�����'!0K��W7��Z5���xn�&���͚
_=���n���:�u�Ӆ��uW�)�;��V��4���
� ���y�T��� 
��54h�@��a'�������<�
���6v��glꎞ��q�UOx}��x�������tB�cP ��~^��*�F��	�Bp=���m�Jz7 3��&�SF9@�ɹ���]JԀL���z���]�&��wJ3gFk�+N]@���PO���J�����w=����\��6�����<mXg��s[a�D &����T5W�?2��u�]��2s���7���i���:��k��~CP�.O��N�x��.q�v%[w�h~S�dz�;_�Z8������8R�\5�0@�yW7�:ع0g/��<n��ZbP��t!U�rQ��[ۦd U`S U�e�2�$t��Qz�y�{������
u�B�'h,�3!I�B( P`r��v��n�1��d �
>e�^�w�0L�ᘜq�/������$f���t�l=����-��|ݱc���������b�e��|����_\���y+�Gk��ß�v,��o>�^~k@m{��72g���Cxy�.��q�3q=�u��D@�	Yx۵��j�:��nll�_`�����a��~���ģ���t�Լ�p��Ѹ)P���"t�q{� ���
=��fsw��~���#�d�g�fV�?�^�}ٵc��B��4�{{nû�1X=����)a������r����R������{9|�.1�k��O��n�w���7�F�{������V�lh�;�k�����h[:/zNnl�f��#��9�:J� 
Lhuu�R��k�j���7�P�*|ZHP���V�U��}1u���������n�S�l�|E����"(0!+p�T�o�3�7��rl`�j���tkk�����RMV�� ��<P�i�Xs8#Ҕ�g�@Y@�	)�Za;go#�X �(>rW���,��[pk.,,Ԃc���677[�e%>��(�q{�B-%�9���0LG��6�ߩ�3�FA�-���&��Ӳ@WKֶ�5\��R8���ݪ����4����Z#�������5l{/�Poz�b$=�}8C &����G��F���U��~��H�B���n������W+;�n����h �0�
�=n�������v��j����yS�S�	����QMTS��j�s�i�����ؾ������Άa���� vBr�g��v'ًЯ��!����� f�_�Z�U�8��7�@|� :i:���^u���v���bȎ���0v��ch�5�����9����+�l]���@����4�v�V����n������8 ����n :�����|�U v�
��=�Z�c U������J��QEz7M�������p�"@������T������q4�z����d0���1XG�/�B(�����n� 
LhccC��W��Oʰ@���!��i&�N��� ojs������(��Q+6�7ey���l�"���R�x��f�h�@:U��8���g���wDR'� �_�-������׮�0L����y���'F-�B̄�����*�q��ݭ�Gyq �d�����X�z����~:�55���JrPOAȎMb��y>��>(��Bh�⯞���$�c�˽\�S�&���f���{#��hc�'bH���ٶ�B��V�ul�k#�����z=��>�HI=8U�jQ!(fB������*=��u� �;��t���<�w���cB �Q��_<c��n~�\&Α^��z�өx������ 
��O�:c�t@]�lv�ou;�.�R������)h�
4�D R��ܻ<v/0r�!N,=sg;䗚@p#PrP`r=�=����\��'�Ԃz�'f�Q��j:рL�C�@ -5( ��d���?@�spУ���5;/T�-<G�H� 5�����1�>]}��a�g$���YrP 8�-��ȌM� J� 
���-��D(u�9�>6�f��d  2B ��>�]����i���(�4��rlb�i�����B ��⮪*�z�|�O�LS��y�k5���w�h�!t�����3�4+Ƚ�`�4z�gLGٕ�'��+�r.v�P@����7|T��n+��Pn�<��ْ���\�X�n �d��.;(P>�L�s���-@��5�*3���1x&����B�#(�P`rE��#_��h܎�8��U����Q�7Zo���yÏ.y1�s�����y?�&b�1���@
L���M[����繥��mbU�|^�� �V�=��(�����ގ��d&q�����Lx� ����
�f�����+8l[��)@(��3�H@�u��-�ly?�r�>˒����#x'��[�t�T��I�(�d0(�c�k�z����jA��s�k�8k��������o�������<W��.�缩�����1c����k��]���N��a��(0�v�]����E5s�V����v�y}?:g����ܻ����}��-��S��ݶ����p���F��^��}�Lyz��Cj��Zg�	9�`�|4�H/)�<Th�[�XN
��p�Byqq���ׯ?����}>j��<����^;�3\g���#�<�:ZrP .��[� ���xbo��:nnn�s�-w��z���{mQ���j���ռcm���D�Q����n?(09�g>lX!v�#xPuD��jq{;=���K�ă�<mˢ���N^j>Glۢ�s�����qb��� 
�ą3{������(��SSs�e[� �� ���b�e[�q��3�_b�&�|���
�R���7��T`�ƚ�(랷��2�	C?�:+���,�A��ǖ�ڹ<�d˃sss���>�j�U�l6��oog�꣣!$;i]m�C���q�%�J� 
�Հ��� �Ŋ�a_�����-χ�pL?��y����h����[b�b^���:$�ڱ��V�w�9@ �M|��nC���A(�"b0�Pt��/ؗo���|�C��}��P������:u*h�d��m��6�Z�F����1����;X0SP ި�x(�xԮ2Y3�gz[hk[8zjgg�?��g�N���{ŷ ���m�~jaa����jX[[��
uq{�ퟧ ���պ�Z-=vאW.�EG �a
�����F�$��|@,���?g����t44�B��BvC�my֖O�����ߣ�a���zj��4$�j>�}�&H�U����~;};@�\ ���9�!��ۈ5�y�~����Z9u���;;;-��v��;[~זo��ތWY����oZ[�;666Z��p�P��-|Fq�k[��j ��A ��gI[.�@�G�oX�ςۜ�\�Б��2�̎SZ*����ٿ�lˊ���-��N�׶z�?l��l��-/���3�N��n���VT����^����4@7��u�u�n���mݙ��(0!� �\�y�v��[�Smݜ�����{��0��BQ�ͪ����-g���b�0��Ol�~8��B5�3��{[~���+zԮ�yP��������9z9m��cC�ǖ�V�uնo�
%@ R�[-O�)�����,T�U���ׯ�b<�Q�z�X+j�E��+>��4���0 ^!����"_�P�'�ߖ���%�?��;�����+m�8^���0��c��@�	���A�1|���,\���h<{g{��P��Y�k��v�}��-h�k��1T_�1C���~hU+x��S�k�d������W�/�ߑr���Q�˻�՞��)\�9�E�@x�Z�����,\,��N����B�/>��cn��Yi��/����k����ۯ��f��MX���զQ���-5V�-�m�Ö;��?b�c�w�����8�ߡ�È��'*��Cm�Ֆ�H����± �����59���|߂�/,d<b�i���㼇)�����P}�ڻXi!�n˝�Y�z�޻j���>{����������߰�p^�`ٴ�Y��W�ߜ���h,����,��\�#jYXX�����Q��k۩]���]�o�[?�Y� � ȍ�$����4%�-h��^�S/rՂ�v��� �s�'�?,�%;�${����X�k��!��k�P�W����,��c�wݖ��-�[�7�5�?�����bg����0G{��{-�9�O�I��a��M�6�ĥ٦:@.@�t����_l��-�kH&�ܖ��b_���d�K�aM��ƶ��^�eX#�_j������}�^���Z��o�8���ɰ��NG	�y�e���#x��z���a��(�o�s-:NH�ͅ�$��[��h4� ڟ) ��؞����5�z�,�<ZF;^��7F�d��<ٶ3��<",|j����-�2oN�p�arP =�WO�럤t��}_���~��#�*���')𲨽;l��dP}o�5i\��ѿ�����@/gml��z�B�[v<|#����A�P�QP`B�>/�sq�wmy���K����t���I
��G�Y=B>���A�r�g��}�LQ^G
���ͭ�-����0��36n" "��N�����;;;�Xa�P��-TI�1�h��r�x��]���_��͂�Z�T��o��z��L&�5���� ��C[^� ����eނ�L[��>���$�Z��j�b[֣�k��t�����A�#����^;n�j����0s�XH�F����!��@(������d��B�}y��=���64&ۓ���W�IJ=�-|j�RՌ��"� ���Le�(��P����5��I�{��� ӄσxm��[�Li� 9�����j����<��!��[̜4B��Ė�����V���|��zz�}V�T(��q�K�3�o�|�n8t�ULպ0s�Q��@��2�)���v�X09ka��A�xP��5�tP��X��Ǽomoo����oZ }7��tG�A� �F�������c�)#�����f7߳������P|���E P47ly���_�����f�����0��r���5��s�����w~~^��rww������(:\#�(�_��-$�Z �`��Ը�3C��>G�?�}�g7q�� r� 
��4eտ��?vvv���j�F�����B������׾~%�_�e�2Q�F R�V�<��C�P��������u]�b'�#��p���|I�~�Ԁnt:�ٗ߱�P\��H�ycz�+o�����}�zش��9�W��K�����h,��ʃ�@/��Qb�B�-?��M[��� Z�����§��?��e����L� � 
xA}�Ql��m[�包�+j��T�� ����?�������������dǱ�4��}�m_~ז?��G�<����ǀ 
��~n˟�rngg�mL��H~��I�F����v߰�v��͖���W�+P �n�K��G���>�www���4 �ݶ4>[�������z���p4��]5�۶�>�k�X� �C ʥ�m��9EUt��n�˂��[[[=r����ag��-��3q�A��m)|�A�~j��N �@Y���?�ұ��������l>��t��alzPy��^r�%�7뛛�j��G��yt.#|N@����=�P՚]���ѳv]��
�KKK�B�zWd+Ym����v>��-j��z'|��uP %���S�|+zOW����i�󁽽�F�ӡ�{ƴ�5c���������m��6���A�^���(�RҘ>��'n-��/sss���ي�S4\��h�?��/à��	 (�J��W��Pb�{�v���zO�^������-s���i���B������US���j5�� 
� 
��ԎP�t����e{��f�y[�6��Ёi���Ӥ��0��c|�ѻf:"|B PvJ���rƖ�www_�0tj���r�����m��4��Hc}nmm��>�+�A�B#�@��[nք>Y�Ֆ�$m�|&��0�Uc}~#0�PHP P{�?	�ڥ����{��h��p��I�v�_�gKJ�zX��ƊZzXͧ6�j��Z͛w ���m��0�' 
� 
��ǃ���`ڹo��;o�򅝝�����P�P[j�5I4s�BSl+:���"�tP��Uh���n۵k�scuuU�T󩡖�.>�B#���|���v���x�^?�h4��4�Ф��c�Е���U�ɪ��S�.�5̒m_���0���~�r(jA�t�N/����~����;B_� uZ���D��j�GCg.��ۃj?��$n����k�M��K5�cˏmy? (( l5zȿ�����-7�������sz���<#�Ѩ�+f��qƅP�z*|����߷�f���د|3�>�!���鱼� �pkk�����o�׷[�������T��^9G̉�D����Dw7664��_����A��PF<�)9( LFAI�c:*5l��www����~����=�����~m_R����c�T�,��������g4kР�_��^��'PZP �)�Z����+�W��}��֣�F�j�Ƶ�^�kAG� h$�YRP�6Wà���t��0��0��T((0�����jxPz
N��\��oZ���-������ٙW��cyI�	�p�dX�tj�*M���f�W��à�Sc|�93M��I�Fi
T2��t�����R��\��Ȗ/��ϋ̚q�X���c�BH��H��F���;��5�^�k�� P�d��K����E~זOh.y{}��o�N�I���g��5=3;���Er�S�M��lK
��~��^��s8�ɶ²iK�HI).I�s��crwv���tO7n���
�=՘h u~?��@��h �x�W�YY�f��v�֝��}���k�io0ܱת�B������ZؿZ)�Z�@�rnn�L�G����	ՒM
^�Ƃ�?��XSݷ�����d��S��k�v�����}��sn�����z�P�?&���D` �n���zB���戾�ڇ�}��?����|��n?ϓ���b�=�����O�^j}δS�jH��qB}���ܳ�뵪�Sf�'X��
�,(_:Yj� 
T\�����MJl
�:��憪G���@����!�����5��
f�9��S����p���ٿ-/e��F���x��W����iyd���zupѣi�E�D^������PdCs���������M��54��x�^����{-k7��?�R���C�7���&��u�VzP;;;S�T:=�v�:%�n:�U�:���z9O� +!�[�;��N�r~h��n�&���uk�b���*0��@\e�"�(��~٤�}@����5M'P�T�T������7�����r�@�A��ZwP`k��}��p&q{��m7��;7�U{���Z8|�.���'Z����n�C��so�O�N���fWϦB�о>��ݵ��-��t����t0��?%5`=�#F �%p��"Q}7=��y�ڵ��?����3�`���D}O�;5��H4���>,���ѥ�j����7VaS��?s��ߎoW�d�NlEH�' ��n��C��Q�}�MC遵=k:��~|��� �7]��S]���T�ԒI�DS�T��g������( ��c?ni�(��l���zG��vG�J'f��@��: J� 
���v  �D   @��   �   �"� ���S�@�za!z E��5G �G���`G���   �   �"�   SP   d� 
  ��A�5G   Y�(��#�   SP  ʅ�k�  d�]sP  ʇ �R#� P.�� �  d� ]sP   d� 
  �L@  �)(   2E   @�������\E4�M  9 �K빊|d��Ɏ#� rR��)P;��� PRP���@�QPjP  �g�3	1Z��"� PU�O  ����X� � �   SP   d� 
��ax  �D VG `P`EA@� `P   d� 
  �L@  �)(�&� �&(��F��  �z�@�Ћ oԡ�#�K���&��  �!��a�@ިC(=(   2E �������   �   �"���^ �	�Қ#�   SP  ʥԽ�a���~X   �"�   SP`a2d ����
��  �!�+
�+��? %��8	5E  �\ʾɚ� �   [P`y� �P   d� 
  �L@  �)(  �Üt�XE �5@ @ء�1(   2E   @��   �   �"�   SP   d� 
�K�  rE   yj� 
��� ��@  �)(   2E �9W ��@  �)(  ��HJ� 
�/ @��   K�� 
  ���O@ @�H�5G   @��   �   �"�   SP`y�c�<  k#�   SP   d� 
  �Ɣ��#��C��� 8��
 �#������T�	�  �� 
  �L@�zb@��A5G VS��Y��  (1(P/�a � 
T��;�Y�
 �XM�[^���w�Y����   KO@�U:�Gy��� *� 
T� P4P���    �"�+h��cD(?6PzP` �+����Y�5D  �\J���(  �	P`E�� ���j��/D�Jۋ������>  wP`EL��3�J� 
,/t~ �Fdj� 
,/�L&P  �D VC/( �!��D�g�@�%�z���j�}(E@�|��X�Vq%����Q@e����H���JW4}�m��� 2�������ZgP`��D��
I�� OК#�5���O�ʭ
��*��� 
,OŲ�s�f�R�r+�gx�<!� 
���#�,}T�ýɒ\8�<�E�Q�j� 
,ioo/�FAP����O��jQQw��ܒ��_&n�!5E �װ�Yʂ��H@��S�u7/�!t�Q�j� 
,�̀5䫔5(�+� ���P[P`IV4�y)e�b��XV�=�5G ��h6�U(�Ux@ݝ�H�o4�x<�������Aە,�������t:c��禟��P6�n������h�l�8��P犮�j�b?W�!��j� ��؍[����U��EOtn�E�g���}o����u?+��`���-�]?==ue�yW�v[grj�kz�ڇmC𖽇#{M����I��v���M�Og�/�T��D�ƚ�H�0�ছn3�����C՟I��<z���{�Z�v۬����O׏��������}f[֢����8�,C ����s�f�i��nܸѵ�6�u��������|�Eߛ���ci���7
��nW5H���#���4D�+�
L��`]�r`�*�]+d#w��+��/2����ŷO�h�];.�����%�Ymd������~�_�yK~Ce��I{Ϳc7=e�=�mzmv9QՆ��_K����}��|�=����7yTt����}�3�ٗ�vl P\�#��O���)�a�n�ڡ����o^��~�k_S��3/l��&<F���#�뒳�X]�i;���g�]v]u*�M|�
͞�ޯ#{Ο֪"V�?����͛���j#�u<y��9�m��3�&��P�����_��f�=�'
�v�k���o�߆�@Qt���M+2����}�]޲µ�ʤ���M�A���)��{�s�'h���_E�oa��ړ*��>D13�^�¤6P����#ۈ���}��gG�k��}� �<�f��{|�~�����[��h��O }ݦ�ւ|�n�Z��s�F(m'���-t~��v���g)Z�-Q_"�I~G.���g&����	�a��v�T��y�Q���w��:�������ǭ�U�i��Ѣ=s�_.z��X�Ș��ƺ�����;�~]��E7��x�Z�!3P��\����ފ��NGUDai�lja��"ʚke��|��b�*f��O������k��w�u؆��{��>[��Fo#��(p>f�/�}�@QL�9{�����������;
�|.VY���wѥ���K��>�a��ЦZj��Z�۶�T�������i����~ϑ�2���S���ʑ���ejS����qT��w��^��O�?\�ZP��pX<�H M���8�=��m �����l=Q7��Ԟ�u��#� ��L�����EK�W�_��2RM�f5գ,�Z>ꛇ��7-�j��<Ž"�(:��x���@�V�7��i�
E>���F�A*�^%O�����f�%_�^��1�
����~*�e�-��)ٯ��h�vv�_�c&�����H2F E��]�{��Ҏ��J�"��+oP
2-TJP������,zm��Pl�ߨ��HB�Ĵ֭<�[�ܓ5=3sm����rP���<�}�BeJٲ�N��(
�Q��Kz�KJ��|f�:���B9�MG��%�!�h%E EYPd*(���r�"���.,ɑ��Yz~��[�g�K�9d� ��K.��i�Ң��u(P��!� ��˴|�"u'x��-���"(�b�C�hS�Qm���z��4���h���(�x�=�7�b_Z�O�At��l��g����[F ��P,�a��R��-P�¢�N��\��#�@Ei1S)��e� �2�P�η [�(͞�!x���(�x��K1ᡴ�c��$�/I����o������%�>A��`3�魞��(
o2�ltM�U���<W��{�(%(j����^`-��By@�(���?����6� �R�s ��l��Ơ2��DiPw�%����(ʀ�  @�@Q
�:T�� �D���	  �B   uFG�(<-D�J����
�N+(d~Wn�(
Dui��r ��19 ���� �8T�莣w	�G�.�ms@ E)0LRY����;���A��g� �L&c�g��R
��u�S�P4�E��i������(6jPE�t�9(�`����ݨWO�^s��W�l�b#�V=��!���Tz�Vk���]��t{{{nww�=x���F��.�Aj
���Y���_w4��;;;��hD���RX�}Y���c������<w��ա��������F�	5���>s����LUk��7��K��yS�����s���@Qt*C+N_��h���̺f'�W���޿�i��U§��ߨ���P�AP\�o�ox�����cQȬr]�5A�!t�U�x�~�?Ch~�(�(�ZA
U��,����Ӎc������=��]����}���ɓ �1��a��G��!x�
@�Z���]��j�>c��Yr�����=�5H�׿'�~��5ݮ�T�7�`�(:�3+@�����|��tAR���p8�_!i�}��1�����)��I����G��7 �=�F��~�z@����
��`7�[� ���*���P����SOT����!�W��D�@�AS��^�k�uv��aޏ�$o��}�P�e� ��Ӟ�~��R��X�ڱBҰ���E$f*}r^O\�����U+ja�Ƚ]��ܓ}ݶ���-+�;v[�H��9�!���pb������{c��[��Ƀ��<Y�)��Tt�iz��x�V���v�;��9�?�������]{��v�a��vø��a��}Lu�Rh�w/�kt_��<Y8j,�!����oܸ1��y�^sO��4���l��3m�B�O��$�tq���*����w�l��v�g� ��S��7T(���=,���$Y��m�~�0܄3��M�}_X{�ڳV�~�ڭ䓩\�g�r�!�u��������z��iA�{�k��D��O�=�#����n�~�v(ݴ�����XE�|�9���/Zzښ��U�&>�g���d����]�6_���uz���N��Y:p5`�S���o�����?swL�6o��d�L����F�z�1������;�e� ��S�W z�=<gxZ������E4>|d��V������;Tq^=
__��ޗ��7ݐ��uiC�7Ѥ��P\��׎����.�].��E�'��K}FT���d29l6���j@��t:����~��������+ι�`��`��}G��1]����#���qˊ��U���;Ƞj!4�s�K�|�§z{� .z#�ߥ��>l5�]�"�j��h4Ҏ��PyP ]�ֆ�������+��p��F�A�*���Y���V������צ�O�'����[#P`����]�/P`�
c5���A �����hT�e� R|Z��PQP`�����#~� �hѪ��KE� 
 2 '�[P�j� 
 �!�V�� 
��F�@��텏��u�D �Bh�@Dt�vG�
��i�k�V/����|u+��P$ArjvP�� Ϩ]�3(��M�P}&�I�9��czTN�O���/@������� K��§NW��+B+���(( ��L��cY�\WP I���Z��ک?5B �Q���!4�� (   2E ʮ����:~���+?� SP��6����C�@jBk0�3�  �j�A V���9  ��#� �"`ϾF� ���TB��N�G���6(0_j���� T5
�F   ��(��!��U��; UAݩ(0�#Ő�t "�����|�&�`��c/�&��6�p��h�Ʉ� s_?P �zA�2
 �\P`>b$  [@ �)|2 �@�tu�u}� �@��� `��|u�����*�e<G�(  H`��G �
 �P �@��Fe@  �)(   2E   E���!�   SP   d� 
���Q�����F  ���0|�/�����j�>	��(  ��0<*� 
  ���]P c] �=joM@  �)(  �E�xG�90	eE jJ�06]@��'�yG�+�7�Re0��ҕ��/@�\e8 �F� "�  ��@�tu� $|� 8�� 
 @1��SH�D�@x��@~�?5B �ծ� ��  �D ��
 oԠ� ��� �V�ѧ�"��խ@��[��O�@xP @&�@���>@����n���� "�F��G]?�u}ݵC �D���O�@D�/jP�@�K�aX�E�k�B �!��M����Z�H�,Tw|��׫�BM��,�O�@�tթ�%4 ���BSkQ��?j� 
�U�*�~^���ޕr�H�zΓfUz@�(3ԡ� ��5�d�{�@AE��V�%_[Pz� 
,��jE=�Ѩ�r���g{�%���K�_�C]4j� 
\B���l��dP[>���y�ե�����r�8\��|h���PQ2�s?��*I����C���;vu�PP �Rge�2!M&����(���U	��^�`0�9�g�@�t*�#W#��X�w� �>�j��	J~4|Zm�Z{�9��B ҩ�G{㳅���������@���g������7x���޽{�.>�ߡ�@:�<�m4+��� : i<_��U���ek��{:�_��P����z�ޛv�g�tY��@I�3�Kk��C�� H�iGx�.Y]��?�3�E'��X8�H��H�YP{ˊ�,�e*����g�o��u��#kw���C���~&_���G�s$O�y~ǒ�%=w������#����n���c�6�@�3k/X����g�z[��v[��=���@�K}���k���pۮ~���N�"x�ڷ�=g���v���~��lF�LuS=����Q-�kQ�.�Z����C-@��^��?���Xk�ak�O)���WWn�����ϭ�� �
����k�����k�����W.^�"���5hK%,m���'''Q=���������o��ܡ6��|oXS ��j��PQr!��eX�l�6��z
���M{Z�y �E�"�a�]V{���oX���7��<;��?O�O�R�=�P���u�;k�s���
�O��y5+��z���ҥ�}(�f�9��Kn�q����@�W��@�o����j�%�����P����j���X{ݡV��|��?��GV��7n������}M���⏎��P�i�j���������R��f�Y��Pd?��֞�������ݺQ�����y�'��4o���Q"?T���P�L�����C�@�����y���m��_���k>�y񑜑"�P?<�� ���v��6^/�ךW�_�tث� �Fc4Mf�jͮՠߵ�`ɟ�u�=+�^�ES�t ����;==�Q�z���NwB�@�˽m�+VL{:����z��*�:�.}���>�+��^?gUG��󭆓�D=)l�n:���	���m�#����}�ר�V��t:��<)�74��du��j�|�������g@��h�俶bߵv`��޽{w_{�ɵ��N���F@�[!�6X��������/��
�Z�!/�\�3����L?a��_v��Cr	�s��\�!���sSO�7Ύ���b_�����c�Z"�˻k��[֞��Ya��v}O=iD'�B��,|w:���iϧ�<!|���՝���a�l����,�.<QF�C�~���U]� ڱ���s�on>�;�X���J���
�V��	vM�2����Mi=�Y��S�l</L�h�Kv���aw��4\�����O[���p8����H�ӑl'X�>_���?�K-���C�@��i�����������?:���Y����)|j�d�X��Zn����� �Mcښϭ��O�����@���������ιV���k�K��yǡ����T�գ�œ��w�Z���P�ù���F�6�v���N���Ѧ�: U�:t
ݯ[{Ƃ�f�z��#:s0�;���_uӥ��9�P���;�oXa}����<S2��>c�=/�֪�A�����i�4�[�~�j�N����T��`��	ͪ&���M��������d
"P��t�����e+�����T��i$|J�6<:��>z�M{nTǙ�o[���a��q�v]�3yPZ���B�mG�K������@��h�oX��D��{�.�]����;�E�5?r �F�F�
x��]��Qo��A�y��3>	ƱPM�Q����zT�u�ο�B�Y��am7ߧ='�^�O�t��yށj��]�+u��=�������rqW��9�K�-z��vu�ͯ8N��P`}Z�N�`:������'���~Ԧ���i6�Z{:��~_�ټϷ�z�:����:Ј��vb���~����j�z�U-�uɟ:8y:��̞XC�GK�%��;;;a���Q�T�Tm��P`3�.���vd{��7o��+���H�� ���u��s�����m#��.-��7��ށ:ќt�8ꔻ�^�7����V'Z�ԟ1��U���{W��O	]k/������� 
l��:��{��������]�_��������ª��n���y���s�ߏ�§z^w �FG�������#����a��N����y�.��^|���n:�G#B
���TP`sTh����n:�7����g��m�q_�S*��V�����3ڀ���}{l�QD��*�립� �I�R���}|����첥�����ՏUFd��I�Ӊ�xV�F�i���?jJ �s@���C+����}�
���h���I+�Q�\5|��v���Qϧ}ݱ����S��َ^v �N!T=��C�����|�jюj�z2W��C��k�`���������`���o��;`(�yw�tّZ{ʊ�G[������'��!���7�� ��
�見;k�U��ԩ���y2��f���_��ٓ���_�~�Yɹ��<���#�#�����7�K ��1��N��Z�~�.?oE�i4�e�s�\��A����F*�:�z:V?� @���ZV3~�vb?`��=W]�cv	'�Io��Y�����V@ �O��
�C�\��ԛ02�K:��U�g*�w��b���x<�%���v���e����Ǐ}�+"�ۧd��}a�k�7a��uG���8 Xl�6t@�L@�c�1䎕@�l�N���ېv���p������ Ja�B�ɑ�(�}�x�H/
�i��)�>,C�bznN� ����n;a��	�<Q�peP ���2=�i�f���	!WD ��0|��_u� H�ZP���eC��Q��.(P3=���@�T�H��(�#z dd[G�S�p%P s�4!@8�B ��H��C�kO+�Ul#�R�p%P ;j  ���m����((P^lP ,-��Ds�b]P �G�&�~n`{@p��N(4^���e�c����qeP sτ�v��%��	�UL��M�(���(��m��� 
`�Q ]�ԋC(;¸2(�����{´�B�q`�jR �jƺ=���F���#G�@�l�H���}X�w�� ��=��q Վ5WB ������; �\@u��!��AHۘZ�� �9��Y�F��`9�;��Й���X�ƅIW��ţ�!} �;?�߰nM�)v�q%P �0�ɵK|( ,cbF[�gM&\	�F�Z[E{g��T�5��6n<G���j�H��;;;�}��at߸'��/ �P�X��Z-7��&�v;�+�/^�(�~NuH�S��O�ĕ@�l��1�+��q�Bgh�ٌ
��3���J(�e(���vtUOD�FaR�R���̆P� ���	�׎���(�U�n��Qhl�a0]F�~���A�3�C��}�׋ �cۈ��k����;'''������~H^uH;��N����çt�]ա����� 
d㎵X�Z�l5�Ͷ�g��5{߻������׮�.�;L;֎�����p9�7�=o��jˑՒ�՜�]o���>e��09(m��7��}ߴ��;v��tgX��Ϭ����t>�uk�e�_�a��z�p�zA	tNOO�i�_����{n����#��\��K������Z�iY۵뷬��բ��N��� I|iw޶�#��ck�Y�����tGXȆ��_��gN����,t����oY��S =88�zBBž���t�®~��}7�b����p�ѓ�X�Nuqjg�I�9����G} �(���t��������Mw|5����9�
�@v:���^��������
��&�H���}���|O ���-)�+�nww��il^��ek��P Ѳ(����8��ۋ�|��Q��+���=�O [auf��l��)gi��3�C 򣃋.���`���N���p��(��O
:�\5�����e�,� 
��<��{j< ��ev���F܀� ��:�~�g �Rښ�iws��`��@$��K��J�C �u��ے� ��rC/�#�b��@~|1R�=���k~X(�(��E �GQ�'j2G �ǤO @�@�|]8)��� @��C�((���u�R�'� P)P��� ��Z��!�   SP ?y
 �%(��F���{ؚ%j��N36� 
�p	 �(   2E   @��  �2���F@�����dnQ���ّ `;BG�D�@���l  �B �z$��#|(j6� 
�h��{q 
?�m�� sP ?�ѳa  T((��r  ���@A�4 ��"��G.�@�(� �Z!� Po�#sP���8  *� 
�`	��E��ѢSq&>
 lOt�#<"KP ?�G��[r��Ph�9(�/
? �v�@~� 
���ј���F �p �*"��!m(�et�`Hl�ׅ�ߘ��R�l�%�/�!l���2L ��灦h8j6� 
�!x @-@�����,�#8�6� 
��|!z �ɲu���"��!�(��2F �C �7�rA ��K�`�0d��6���@�|��  O�A�%�7q�+lȏ�y���l6�d2��_���j�^��������p8�o�7���Ij;;;����S˄T`il؀���\B��?7�����-�/���E
��v��!ݧ��� (��kw����nt���	�o;�� ۠��Z�ߠї��]7�ٙ���*���!P ?*�oY;m47>������ j����U��m ۡ��7��a�i�;Q���)��S��ݴ;`C�@~4��sk��3�w)���.�+�]k�; ���l��vym<��`�&�'4�������!P ?����ou�ݧ�0|o��k��f����dW�sP ۥ��oX�����~j8��ӌ;��j����@�1P _�y��x<~�M�䟶@h�S������1�vݳ�kߵ�yh����c;�o��oY���w�AP _�־�����|&�yМ,��"� l�0���?s�y��X���k�s�p�s�@���bM=_�֎oS
�a� �O;�_��mk�����n���aP��E@�N;��   �"�   SP   d� 
  �L@  �)(   2E   @��   �   ���-��^Iv�    IEND�B`�PK
     uK\�T�'}  }  /   images/1be29400-b52e-43b8-b531-83e2df2121b6.png�PNG

   IHDR   d   �   ���[   	pHYs  �  ��+  /IDATx��]{�W�{���e�ew!-�)Hy��Uch���F���E�J��I1�6�D��5�F"m(IQ�5���X5�G�B ]@ʣ-��
[^��}��w�9۳sg�Ν;sϙ��K枹3g������ǜ�;u����������I�&Y�T��f̘auvv��)S����\ضm�γ٬u���R0�
a�����˗����2�LN0D]]�u�ܹ1$hpp0�	��$���'G@:�΅922�stt�jll�.\��ڵk�kq�BZZZ�����0������%�\�7!]���8�H;Ka.Z�Ⱥp����Ur�#'t� 
�o���#�y8n���2��2�I�<z{{�8���ٳg�r���ŋ�ǎ{��1�v��4Ֆ����w3�t���5W���������\O�R�xW;��ր��$��.��g@�/����K�FB��ՙVB�`
�B������!
C©�*������~1s�̧�|�����S�u�]�~=W*@�CPS!�[�p�9I�9�9�m����n������,�i��F�6u6���� �W8n�H����gΜ����A��(��W�����|�r��ѣO@����0�}���_DX�n���?~<W���,Za�`"E��n���J�u�gW��A��e�C��n�-(�ŵ���P����;Yq��'N\AI{��ZaN&��$�E��%D
��?��d��w��r�JkϞ=���y��m�Y%�+5�5��Y�C��� ߥ�u�@!�U���#Hȝnz�OH�"Ka�w�ݻ�[~��gˬ���)�m�����Ĺ�ƶ��U�.]�e26�˅B��ۭիW�w���*X�E5����3�J+f�G�p��-(V��t�U5?槦�a��SzZ��)N?2�{7^��u<��V�	a%Na�ڵk)s���A�஁�øD�A ������$�g��r�8�｟ꑄ8K������{���`6��|�[Z�Ik�/��:.�V�Aa�ܴ	mt�Q2���k��_އ{� G���%����q����X)�p	��}G��#��#���25<ٛ���0�V�9����1�?L�K)����V��Î����@x�4ܿ	��P�[iܛ�/<�N���҇R��q�S����,ى�'�E����A��u!�,b.�QW5z���Ի�+���Q�{.�= �_��\�i@T�%�鐃t)��F�(��K4�����*s�4�ď{��Q�t�e�}�UL ��&%U�����	]��������`$!Q���'�bKˊ���HB}oE��U�p%��l��F1�7L%$�\���j��a����D� vT��r��SZ5*|�S���Z���T1aT�	�(&!�3o1oF�ʊ�#��oI@5����d��T#!�`J���q��؇0��H		-�8$��0�~U	�j$��d��!�u褆B$���F2���������k
&T	)�;�Ķ'�@n �JȻ��d�PTM'!%�@c=P����(IH%gV�SY�*�$��2`[�������D./G8�6,&L	I�:��`�qJ�YMxBg+�/!ai�=p�M��DFJ5��D�FȻ0���bL%$����e�S	��H����rdХ�D^c~���Y��k(�D"$e�W
&f�PNV��j�����J��'R�ؗ�0ݔT����F����@#���6�9f�����(K0!릪)!a*��m4�\%����c�A��6Py���zEXQ�$��q|�,��Hkb�	��}@g��;"�{��f�M���N���V_�)����<\nD��R���V���=�tÒ�-Pμ`�W����K���^-ev�8p3�L&c����n�����X+�� 2�{f�|�(�'������7*N-����e����n��(�h�$���$��4����l���&�<[ ta�[�y_���wŮz�+�Ax������S��va�`��{��	H-n��v�Z{۶m�nvEqUK��|ګc�l�L�r/u3/?N0wSpbۡ�&) � �w�}����]M�	�ϊ�|%y,N��p���ڈl�:���u�/ؒ�;�@�#��ݣ��U}pӮ���sw�a���L9Sߧ�t�ℐ���*tn���Ll�E#�i������TSi���ЛH%�B��zO�ꔛ�;�e����0�ztT42aUN�ǲ�u�"����IyU��B ��(��tK�m0�yF��#3֯��E��+f-��07l��"�����(�Ͳ������e�D�%��Nj��m���6�ܦJ�a�gˊ}�m�Z�]�
ʫ��w8��Ȇ��"�_E�2*����6�3��_��IRD���������|>�Ν�UYʨk��B�����~D�=��5z�_��Cܴ�?�{-n;�	����ڭ�h٥-��bst�B�ܹ�E^s��]8��I����V��3g�u���ғ�/���Z�B��p���]�R�|�/.P����vPU�J�F~�s�(�@���g�U� �����^�޼!�O��i@� 7������K8n�Rց��A���s�{`*!���j�C� ����f��p��b�,��.�Ӂ��p�������2Zv��c�'\
�����s箁����x��>���� ���RU�(S&8F�:����YX"X��:u���Ļw��R<�ח�	���w/�ܟJ�d<LD"U�
I�B�Qq�+���kr��ji���$�j�h��[��L%@J��SU��5n�epQT�� T;�L�3a��TԶ�0I\cX�0�RO&�𻁘���5B����:7�%d��F�a��������V�!�2��CU]����u�wvVaPp�	�a\�%��
�%~��Ɲ��"̜�X	a��-[f<xP�~ʭ�g=�O��Q�yQ@L%�[����l���Xr��b<��o��otvv�ŕ�$>㳦����1��ا@�<�Q��!��{}�Cb���G��ʯ�z��ݸ�!�@x��p��9�FB��R��>�����ϯG���\l�)�wi�����X	a�������$h��C	19��xn�:.Wk���+�T�x���,��O²dx��g��fu�
e	���#d��驳g��2�]]C���(y�F��jH���4��-;x{��:�g�L�N���(%|�U���X	!TYvB���#�WN���R?p� +ƴ�J	��&��\M��r��A|ͬ+���	9\QSY��CL�,X��B�$*�Y�ϖ� T����E�"�?�?�gJY�tŦ΄�;��i��������{�5~��� c�Xv��wϼ&��#:�/KA�����K�d3�M�
��"|y���/!�I��{��Y���q����������X��Ɋ��4���4S�?���uF�_�j���cY	�M�5�jEb�Iձq�]E�(�X+!��dB�w&u�L]����8:|�����)a�-������AM�15U�Yr��,}��u��TB��!�G4R����L�����,!��2�:�
���E<�"Nm^qű/��(����}O��Yg����466����k���#����N��bh�/����'�&�����]�sRu�a��H�9;E�ʒ6~�M���ʕ+�d2��\gp��y(#)nТ��Y� �M}@七��I��_Sz� �q}4��NC�>+��o�} �9�E�AhieI�H ����z�9%�5�_�\.�쏈�0
��%!�侎�E�L[��	��F��̳�T+]�� �	�/��F���$��1�߰��A��?��-k�g�l���褕Q�eI9�/�Q��(!���z��#UG����~��	���V�b��?�t)��7��{q�&�>�E8���&/�v���t��	ən��K�mL3����V�i%d��'���uP �Hj/!52�����%����T"n�K���@:��R��ٔ��B���7�p}�~�UU�@;!���q4&�t��ߍ������F;!"��a%��E898Zʺ���?W)!	۟��    IEND�B`�PK
     uK\�}���) �) /   images/146a6d58-0553-42c9-b8c7-03425202d69a.png�PNG

   IHDR  �  A   s���   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<    IDATx���y�e�?�Ϸ���{rL�쮞�8���D@DQ��\\����Sw�׽���o�kw]�]uՠ�r� �A#�1�LWu�a�=�g}�L6��]�OU���z�B���Lz�SϷ�GTDDDDDDDd�e: ��E:Q��E :Q��E :Q��E@�t ��U�V�4�g��Ed���S���e�Q�9"�c:#=���Dd���pPD�=���f�7.ܴaÆ��KT�t��ŋ����z	�� �� Kͦ"""""�4l��U�n����j�t�N��NG���ۯ�oUճ ��-�����:�U���ܞJ���f:PR���!�����{�l8E�/"?Wիj���ر��@IN(���}�OE��ƁDDDDD45�E�|�\.o2&	X�;������ϱ,�S ^d:Ŗ�F����R���t�8cA�@���? x��,DDDDD�
�Z��/�T*�1&�X�;H�X\��_�:�Y�����(� �\��>�gԧ���^�:�w�ޏ�[ Y�q������3TT�/<ϻ�t��`AO8�qN ��sMg!""""����j�z�Ν;��u,�	V(.�/�6�������:�oU�|��6$�X�h���s������Lg!"""""U�	�u�`:HT��'L�X\��78�t"""""�#����~XU[��Dz�������� V��BDDDDD4�k\��� Qb�@�(�%���s"""""��7�iժU=��D	W��X,�DUo0�t"""""�ixز���6$
X�c�X,�V՟8�t"""�NcYl�>�;�:[Uq�u�x��>�t_��xŶm��bz���yǲ��pLg!"""�T�t]]]�P�g*�~�7&����<8��&��4�<�{��6M1�=����q�e��9���0�E��?."��yc��������ؿ��u��?��DD�H"�l6�T*e:J,} ��r��oz��^����Y�cHDR�B� g��B�3�b;ٯ����'{��~�|����0�9E�n {�KU����"rPU� v�H����"r@U�m� ���e%�aU�����y�nذ��r�ʬ����HVUs�V+e��< h6�� �eY�T5 '"Y =�:ϲ���:ODzTu>�y�Ke.F��[K�L]]]�cP��=i0������ED��\.�������P�X�������b�eq&%s���h�n&�f��h�V��n9�� �� ���N١��Dd����}���I��{Dd����Ӂ�AD��K�kYֱ�T�8U=���_4��ǉ�  ��Mf&cYr�,�&��z�Z�t��j�Ꙟ���tX�c�X,�JUoB�ض��ol3-�S-Γ�7�<����a�Z-�Q(�|�o@e����eYe [���J�2d0cb���X�bI��X�`Y�U-���(���lR�"r��t�v�y93��u�2��X�c�X,.WՇ0�J�x�T
�܄S�D��9M�6 �l�YU7��&U��/_�u������}}}��j���+,�Z��+D��
����&���m�l����	)�  U��R���ӞGgA��b�x����t�vbI'��*�*:��	U��eY� lR�͍Fc3��I��+W.h6����٪�l����f�Q�uuu!�ɘ�A	��r>FD�W.��f:G;���D�X|��^k:�	,��.�f�Z-���Ь40�
���<����e=������7�3�����_�l6���}��| '�� ,7�����m�r9>RG�Kb9��s;iԝ=��|���ZDV��b
K:��V��^���A��xTD�}�a���|���q�f�q��"��|�?AD���yw:
�FAKp9 ��������.,�1�]�G��S|�G�Z�Fp�T�k � xTU�G:�.<�5�w�I"r�����<�Nth9���l$����E��r���� ���q+W�\�l6�-�%���!��:E#e� ���~ٲe�*NQ�8�B��O�,�U=EDN�, liȲ,d�Yضm:
�P�]���u��M�h�+
�&"2�#JX�i�x|Z����=���U��t:����@�t0��X�jUO��\����� ^�Xӹ�}2��c�ii4�V;�۞���y��s��=?��%�Fc  ��X�i�x|Z,��C������Ǟ��2�(L�bq���/�3D�_U׀�t���t��N,�~��+L�z�9��O >n:GT���t���Z��f�i:
Mn+�{�#"�������7�:��ŋ�f2�5"r&��bd���p,
�c��tp9 ������t�0��GToo�1���g:K����T4�MT�U��G�+"?�˲�ڲeˀ�@DQ�z����ݻ׈ș�����5Cbض�l6˲LG���r>�G��c:D�X�#�q�?�%�9�%�ƣ���jh4�OX�<	�'������!�=I9�s2�����1��>�p,��l6�t:m:E ��!���++�J�t����G��8�Xc:G\��ӑZ���*|�7��� ���Z��T*�'L"J�R��ޱc�i��RD���5n��T*�l6���:��ө�<����aaA��B��l���q��DiL�;E>�� �����˖-��ǝ��x���t�T˲�p6�~әh�,�BWWR���(�f,�G�[�u�c:DXX�#�X,~FU?i:G��w6��Q�Vy|��T�f˲n�}�6�Nm+V�X���kU�� �O��^�t�����r����a`A� �q� �5�#��ͫ3�����ܯ����R�<��?�(���|���ܲ�׏v�t&�� ���8����[���z�OU�r���u?j:DX�#&��?ײ��M�;����U�����"ru�\�j:����x��� "��Kp���d2���2�B0�rnYR�����' �*|�G��B�^�mYW��=�{��a`A��b��AU�w�9��%=��j��p��^_��n޹s�~Ӂ��}�Y���X�u����ә�Y��\.���d&�|6{4���Xn�+"�$.��GL�X\����˲�� 8T�Z�Vh�%=�x|Z�Tu��|_UP�T�W��}�&�����ͯ�j��VU}-x�[dtuu!�ɘ�A�4�r�ｪ�^��^���ux���m:D�X�#DD�P(l��t� �R�R�l۞�$>j�<��di�Z�y�\kY���r�g|���!��w[���,k����Z�� 9Ɋ�1 �������f,�:����sEd�Q�a �џ� p @������.��j�v�}��ڵm۶��O���+Wf����e�AU��%�3u�T*���.����t˹eY�f���E�l61<<���W\׽�t����GHoo�|��`:�l���V��Z��3�,��P���xw7�6�ڲ��>h:����bG��±���wU�� �)�=�b�DUU���U��˲|��T*[;y�DDR�B�ly������M�l6�t����t˹����;��11+�]�}��AcA��B�p��|�t��rgѱ栾FY���j�Z�����*����߫T*�C�!"�dɒE]]]�|�_$"�Tu��.�������=��M#+��x�y��]���r��l��|�hY?#7d��x�3)��lvFϛ��� ?�J��EةbA��b��W����s̔m���r�~3�.^*�B6��7��P�C�Ѭ�p���Woݺ�FU��dٲe�R��R Y��KG��h��K ,���6k����eY�����<�nl��f�q����g۶�U} >$�F�(r4;3)��ڽhh('��	�r9�ȇcA��q�	�ݦs̄eY�������w&U���p,�9DT�"����6n�Ȼ	���7�^�; ��Z�e �"�@�R  K ��hixLU)"��"�p�K{oo�1��+"��� �M�M��M3���;wn[~/U�}�v�u`:D�X�#�q���1�c�Ds��	�â^����J����{=
�O�1��"�t:}ͦM���D3�z������-�"r<��c��X`�ٔ��� �GUf�������6*,�����"r!���<��ǱE�L�y�V����l���fBU?�y�gL�z�8����9�+�˵e|*�Q���QUT���3��A _O�R_�b:�N�P�UD^i:�$���Ƚ�V�����&mFD�|>�2˲ޫ�o�X��ZM'sf3:gΜ��d�Æq"�r���s�="Fw@�ݡζm���=���Z-��,���l6Q�V�j>uU �cY�������U�
���ȿ��A�� �(��}߿=��ܓ���/^<7�ɼMD.p&8۶��f��n�l
��`�ܹ'�������Q�6��u�7�$�}6�)�9��]��c�ذ�%ݼj��F#v��Ly�U���g�R���0��K�.N�� ��D�_��=������}wRV����� .��p�����B&�}��e���W<�St�r]�e�C�="���cYV�t��j�Fc�:�!�N#��iA���Ӧl��~���=b:��X,^���Z����CI*�W���۷�-�� /W��	<�LAL	��V��s�"��r��o:G�X�#��������jCw���Q�%��j�����Q���[�u����n�a�}�y���A�6$"����|߿'��q�gx�����,1�'Ix[�����}\]�}��AbA��q���t��h�N�c����k�����}T�U�6���}��r�R��t2c��ՙ�{�np��,� �#"���-q�%~��ՙ={��ID>�e��$	�c^��Ҙq��y��\�Mԩ&,�Q,_��?5�c:L=�t���P7�`IO���%�& W���5>[N �8ο����L��ݲ��������n���q� �] ڳcm�Y��l6۶MG������,s�����l��u݅�C�="XЧ.�������R�����W*���;�X,�Q��M砎��0Fw�_�l�]�ׯ��Ν��,�Ȧr��p�D05%�A��1���)Ǭ���ǂ���ñ�#�oR1W��g]����0]��<
��9�� p'��}߿�R��b[��/_�r˲>���r�����	�݋c19e'q��AЌ��y���9��Ē>3��j���E�m���{�պ�c�4E�p���q�8�9�e�q��Y]�!������G��np���� �F>��chh�ǱMC؋�F�m���5��@Dx����q\A�?jc�f��O_�����0W���C �#�J]�[��b��\U� ��EQ1�Ǫz�y��4�e˖-J�R��~Ǚ�W�m#��²,�Q"�]��l�t:�� �;m'�ˡ�j�ډ[AgA�Sݶm��?��v}H�1��$K�Ԩ*��:�O� n�O���e:ŗ�87x��D�x���e�P.���^�|�۶�T�c V��W�v>�'"����fI�����P௛��J��.�,�S}�H����h�6��۳qjXSŒ>�V��j�ʑ%�p���]�\^o:�_�X|��~�t�ɨ�v���j�[w��q�t�#�>��z˲.p��<q�J���fy�({�ض�\.��A;����,R����Y�'Ƃ&z6�����Q���(��Ȓ�L�z�S��T�_��C��8N�� zLg!����ܧ����m�Ry�t�#�������� ^n(7-G�Ner�s˲���hI�M�Hww��6dA�zD�.��H���J��9sB����Y��W� � |ݶ�˶l���0�L�B�k"��s�¯�Ȳ��6
?z������aZ�&1;q5=
G��r�\ ;�7�MT���WΏ��}b,���������i�T�qoL��@��}�X�y|�m"��z�~Ŷm��C�����J��o5��( � ܨ��7�����|���ٶ�I �'MY�%1.�P���d��dft��>j�Z�;�O��<��X�#"*�VI����:����4� �/���R����:��X�B� o:Q�����F���m۶�0h�ʕ+���� \�6%"rh5=�~m�N�'�Y��h�Zh6���snYr�ܸٱ�O�="�TЁ��� u�C�:��w��y��T�+<*�L(
�OD��t��D��z����T*�d�B�P��� ���,q���آ\�'"�m�Й�"U�����P�t��.�,�cA����1���3Z)M���d23��n4���y��SJz�Z�.k� �����F��2%V�P8ID2���M��"��f�y�֭[7d�ҥ����� ���>%]]]�d2�c*.�ܤ�V�ǰ�O�="�ZЁ��t`�(��Q��F�}�G��@�ٌM1?\&�I�XW��Ą�����r_۸qc4v(���8ί �6��Ȁ� n�,�����{L���E˲>�" <|IZMg9��tueA�zDD�����Z�u�C��Q�$|&����1���Y _��y>�wL�R�
�O��gL� 2IU���u�e]].��m��X�|y�m��}�frtuu!�������Mw*􉱠GD�:��#�S����9�w ��e2�ܴi�^�aƳbŊe�V�r �X��Lg��]� �%)�`���DY_�b��V�u)�?�g�P\�cc9��m����֯aA���Ӕe���=O�(��>��z���vR9�YU]��Q-�"�r�#�V�	 ����R)��4m�J��n�9�"�����w�P(����덷l�2��%�e�PU�k���Q�����P�N�a9��m���b�X�iZ���G��Z�ǎ׋c�j �@���y�.Ӂ�S,�,
�<�������m��qC�Ȝo�@Q������M�yޛT�4 m������8�k�r>�T*���4������+c�a�[Io48x�`��nD���:y�뺗��[1h<+V�X�8�U�z'��LD��q�ڛ�L�d2�02�ADOw��M==����y/�6 �1�#��Vӣz��r>�t:͕���ӌd2��8Zl6�P��t7; ���K�����ry��0�9�8�D��3�{G}�F�9��FUo�@u]���V����3E���G�6�e9�\*��B]�X�i�:���وrIo6��{lʪ�^��N-�ˑ~~�q��
����q��pԽ�p̝��m�j:�Um��{����p)�H�ob���V�ahh(�ް�O.�� ��q�=d,�4+c#.��:�z��j�j:��T�Uwª�n ��R��x�wU����q:�s�x�t=G�;K*��	��':�788���G�T*C��^��� |@4�j�Z2���r>����)|,�4ku�\�шDIo�Z8x�`'�� pe��x�뺗��?""�B�B�<�x1&g�G�;���@UD~h:Q��b:�D<����G|�_�.�y�fl5�������hk{��S �Y��L��z��1����\׽d۶m;L����8'
����7 �K��cǎ?�u(T���3E��Ff�}"�J�!�u_���0�'j��&<ض��Z���$�9t���S`x���L�t��144�g�""����u�s\��h:�D��|��8� ��ڪ��u���� �7��ڤ��!�������<�G�3�'JƎ}{۱�z�W6��e�6W�'�h4�V���z�O�,s��ŢE�n�<��y&����`Y�c �#c�A� ����ɧ�M��t�X�y�.�!�kÆu�u�`��sU�k ?�6a�r>�l6�rn:ζm̙3�+�{w�NY5�f�X�p����yg�q�<ә��8N�q��[�u�ސ��$��w���g�}<[�ly����>�~��<Q���_ϰ�O.��"��}~SX�)�eq�}a��F�����D����i,\�===�m{����d��)�Ji�q.�[ ok����_����z?2��x�s����f�R�����U�� b7��&Y�'���X�cA�а�O.Ȓޮg�L�J�    IDAT�?.<�7��@�q�����o��s ����o�QիD$����6RU_Uי�AdоE�%f�YU}��J��/�� $���M��86������J��4t
�eY�3g,�_j�	����֮]OM���±�;�/)�J�mW��nw�eY �7��B��1��Om`Y�ܩ�ݱ~��ĝ�y����r��"�R �2�'Jj�������r>1A6�=|*�bk�ЍݑcI�lJ�L�Qŉm�8�c�`���~�0�Lq�u���}@������˟g:��\.?  �'�EDn3�!L�r�n��Nw{�V���ј�����D�\�+���Dm��>����U�z���9sp��Nwы�:묶�9���8�sF�a{���m�?E���c������DT��� <����DI�Z���>�󉍕s��G/بm�J:?�7���������'�D�t:��;s�Ν�K�����0r��P(��h46 xO;�wN+
2������Mg 2�7�ry����n�u�7���Fps�CƎc;�1�V����aC������łNm������qWœ~|�eY�6���׈��e��������m"��q�x�Y�����x�!([�n}��9��IDn2���J�r}*�:�W�M� <s�ܱr����fkl#gN�FW�>�2�Z����>v|ZRWͧ�	ܔ��^��. �x��r�#��?��g��>����W��*$��p�8�4Y�````��[�u��>n:OT�]+������Fg�nH1��������V�,X�7�L:�~wP/v�|>r�P�����{����D�(:
��|\M��1��w�a����=K�.}!�K$wS�i�}?��KA;]��꣍����rG=ϚF�j�D����[5?���b�|��X,~.G�͊��s�X\n:oppp3�L� j�������_����� J 4���ɶmtww��� :��fY�'�Ļ��ea���?~�#V/X�f�� ^(�Ͽز��T�����i��@U�4�B�}��ڤc�����<�;#���ܬ�fĲ,�r9��`A�H`I����8������{�v��|>��8�e�e�����/��A�K�RW�c��n6 �F�d�\U_��y�<۶9�3,��lv��]S����ϛ7���$.(�J�3���b�%�e=�H�g��~���_b:k```�_��A������t�(�<���J��Ͷ�#�%⭫��%=�D��c�=��v���GU�:�_0�j��w�'V$[�׿`:OU`:Q�8�>c�� � x�tj�T*�g�c��"����-����T��r�|��y�YD��Y\�X|�eY�!���G����M�`��C��cA��u�f���@�t
_*���y�%���)�� �͚�A�s+�z�� ���~ `��/+�J�&�	}}}�ǹBUo�ۦ\�����r���sPp\���Q�9�BR�}���C��ƍk��~����K�Ӽ��9t�,~���0��z���u+c?x�����<����b���j���ţ?��,k4�1��1wJ�;+�ʐ�q��}�l� O�H��.���:EZ:���r�]����|8���L p�y�����V�Z�3�j~ �P�H�K���KL��X��1wJ*����ƍ���{���f&�(�L���&:E^*��Jz�)�/����9�κ<���03z[شi��c��8�k��z'���Rկ�\���bpp�1U}�t����\.����i:��y���S,p���R��"�Z�u?�aÆI�r���!�3X�uQ__��b��u 7(��a�n4�2��UtJ�M�{,P@*���y��|<�-���r�Sl��Q��Tuu�\�e��Ʋ�� �B�uT�z���Z�U�y�N'"�����M���9tJ���D����~������t�:O�L,�+�ms%=� >Z�T�\�T~?�_x�}��R�B�uT��ݻӪ����C)˲�{�JQ�y�# ~c:QPD�=D����j�~ �6��&��fY���bǶm��������m7��,��jᩧ����1è�hM>��c�!(0�c: Q@ڶ���B�cǎ��{t���<tt�l�t�t
	:���J:Kz�}UD�GW�f��㏿�P��Ʈ]��h4�|�D�O���o:͞�p̝�ⶁ�������,�z��Lg����r,�	ǂN�ŕ������p]wx�/�nݺ�o�>�3���={�`߾}\5��n���"��{�ry=�ͦs���m688�k % _4�� Aww7R���(2t�5˲�����r�~�E��~5�m�Z_���l��V�صkj���A�D/����6�q�� D����jF��;��GT�B L��T"�l6��1����b�%=<���j�Zr]7��z衍 �	�T����޽{��~/I D�sK�.]l:͎�r̝bMDr]�b:G'�<���t�N#"��r\9� l4�c^���&�K=ϻ`�Ν��zU��پF�^Ǯ]�0<<��{z�c����L��٩T*�(��A4S��s�=*�� ֪��Mg��e�����Sb�C,0����u���~�f�y5�}3����={�j�LEGxg�X|��4s��-��t�Y��t ���y�@�t�$��S�bA�D�٬��$��~ю7{�GX7�_�l6�k�.��&���E��3��f����Mg ����J�~�!��\׽RD���,I��7;�)qX�gD\�y�9��>��7�,kZg�㩧�B��+=S1��~�t��e˖�`��D�%"7�*7��r�|w��|!��Β$c����w.��S"�(�i9��绮{���}V�������<U�޽{y|�9.
��A3�~�����j:�t���h{��'wz��j �?�	,�9sx�p�cA�D��rH�ӦcD�& �{�w���:�*��H{�ZmW$z&KD�,�J�S��1w��F:���t���6]׽�� ��W�m�����X�)���,Wҏ� k]���� �t�* ������!�ڵ��E�	۷o���4c7b����g``��fĄ����/0h:K�ض�\.�rN XЩC�r9d2�1��Jϛ�����vU����}{��������F3�7+W�\a8����{M� �*�x{�x��p��\০���9��:FWW�݁ay�뺗�j�V�,�:t&��H{�V3��nN�����43"�1w��V�u��4}O>���l6�*��t��K�Rk�g`A����f���e:�)OxY�\��� G3w��xrxx�v��s��{M�Px��4}����).6W*�ߘA3�q��Z�\~/F�K�Ԃ@T�R)�r9�1(�XЩ�d2�N,鏶Z��\׍�Y�[�lI�޽�����3��@D��r���s�����; �5��h
8� �祟��4,�4t�H�L�l�t�v��V��x�֭�ݴ�q��f�y�^?�t����f�L����n��e���(�˷�Z��l4�%
��t']����S���/z���;v0d<�b� ��r?*
��A����)�g2n2� [�n}�� �2�Ť�kO>sNaA���N��:b�����U����"b��ό>�Q�x�D��E��ƈ�y� �e:�xD��7r�Єq]��l6�j �2�ń�ޤY`A����瀞��r��旅�g���s���U�� x9�Nr�#�C�ԩj�ͦs�GU�5��±q�ƚ�y��Mgi'۶;q�#�!t"$������_���'��;�l�. o1������bŊ��s��q̝"�iY֍�CPxTU=��K�@�t�vh�Zh6��=M:ѨT*۶Mǘ�GE�J��� ����/�,k���b:���j���4u�t�f u�9��⧃���M����寫�k�!;�W�U���,�D��Z���3���e�ٗ��[1�e<��|���Xl:�ⵎ��t��M�6�p��DG����y��e� �'�EUQ�qk�:b�����J�u7n���"b
�p%���<�/����7���c�9�m����ڶ�� <d:K��G�iR,�D������_U#�i�z��L�P������,��j�ʳ�c²,!��G�l�2`:�ߖ-[���jg��t������ڄ�:^L�f6\���g���s���{�w��Bm�G�B�T�!hr����<f:�U��t2gǎzzz� "�Lg	Ş6�XЩ���C� �7��{�� �Y�r��ѝ�_m:��%"W�l�xPU�F���?4���ڰaC�u�w��Mg	SL��MXЩ��p�h����v]7���bqU�ټ�;�w�����A��,+����[�&�d����<����N	!�נ�&,�Աbx�r����R���t����ժz/�g��Bf���9��7��&f��] �M� �Ce[�ø�{���#��%NL�8�XЩ#��CQU� 8��GLg���˟����Ǩшy���L���T���(,���j��r�k"�v$�Fb��XЩ#�l��1 /q]w�� �)
/�m�� ���B�!"�(
/7��&&"s'��Λ7�.�!(���� ^`��,a��5)�:u��ݭ|����z��2�B�p����8�Y(zD�K�R)m:M������M6l���A���]"�
 O����MuR�XЩ���C�'�j��J�����'�ϟ""w������۷�t_�\�  �7)�,���j4�r��������t���l�BƂN%FcD�f����ܹ3��\���ȍ ��B����0.�T�v��c5D$�'�P�T*�_H�Jz��Q)d,��1btw��K�,9w�ƍ�]������Dd��,s�a\��52ED��m:E�I'��/�J�X�dɵ�w�B۶MG
Ț<)D)���!.z���J��n�u#{'aٲe�R�ԭ zMg���0�+����tz�z�~G:�V b:uU���4��������7�0�J�� �m�c���ݻ�j�̆P��@*�B*Ŋ�ɸ�N!cC"�J��.U�l9��뛟N�o�\�Y(~�a\tm۶mFN� j�T*u��=���'�J�/���l��9-�cl��Wf�p�J�J�W4�Q�d�����^���� �q'�z ���B�5�a�gM���	��A塁��-�CP4�z����;D�By�T~�eY�V�cp�7%cS��l�t2�+�hqm�+<ϋt9#w��4��b��E�OL�����	����k֬���ln�+ L���+�IZI����$9_�DG�1!U���y�(�P(>���2���0��A����7�MD���3P�����j�ڻ������ڵk���>������^%q%�Z�bΜ9�� ��߄)��~�QD>�yއ�^�ǹ���A�1�a��M砧s]�) L砎��r�̯�0<<�!U�O�q��f͚W�J�u��|���'i+骊j�j:��N����������CL�X,��ӦsP"�+7��$��S[��զ3P�V�Z�cY�_����ݻ�V ���?i%��lFz�����N�����}�<��X,���� ?'("���(BD���BU`:�笳�ʖJ�sm�~XU�����0����5Z�Jzįi)��ĉ�h��|��DyC8 ���}���@��,�h�0.bl۾@r���T*�A�����/�J_ؿ���u�juő?�V�a������.��J�mۓ���{�Iƭ%�Qm����z9_�t��T*�#9�tJ����� �a:���8� /4�����	r��'/�,�<�?"r�؏�߿ܕ�F��ݻwc����h˲�p��Dl76ꞔ� �W�)Q"<t��y�j��C�J�t:�^'"+Lg�� "�søh����@������T*��f͚+lۮ��v��7��IL��&�z�P˳eYX�`,+��'�׸������h�M�l��Q/� �}���R�9��pø�}����z����43'�tR�T*}���#��U�b �G��L�L���ݻw��h��v�m�X�pa�K:G�;�$("<�~k6�}�ƍ#�p��|��M��s؆q�5����N���G}�Tz�իWg���^-"�I�Ro�$���hL�l��/X� �Lf�q�ʶ�C礇��{�8���}+�hTD�~��jo�I9-x���W+V�Xf:����N�9(�Z���c�T*=�T*]��f]�#ǣM����?��RU�޽;�ŖT*�@DB{�v��5/��_(�":ھ��v��q�t�����>�w��S��y�f�� �g:H�SU-
?�7��B��m�֭�Ј�3�8c^�V{���������������݋y��!����5&�N��`��Џz�ب{X��y\A�X��h�&۶_��S��Lfٲe�|߿�|�Y�D佽����s��)4WG�$�N���߿f͚+���VU��L�90���l�*��ۇ���Y��D2�zzzB{�vu�d�
:�Z�|�Z���-[�<i:�dD�.
��k:�(���/�ȋ���q,���G�ڵk���>�?�f��;44�V�H�}����}̙3'��;RWWzzz�w��P^���*�̙��}z&t�����Q��n6d*������t�#��8��y��}�˲Z�/����c:D�k͚5/�}�b o�	����R���?w��@_wL6����3zf>
ƦH�٬�(0��S,Ep�}���s<�{�t��(����L� :U��ҥK�Y6�)�T*C��[�9(9D�Ufy��m�ڵ���h�}߿#�v��B�����������V��!��U ��S,El��aY֛]���� S�8Ή �b:�
�t�� ��� �LD�<�9(�{{����u����QU/�W e��jahh(��02:��~hύϝ;����{�8�<\A�؉��BU��f:�T���� �]L��˗/��f=b: %Ʈ�[��i:D�X�v�J��e=== �F7|���vc���V�سgOh�?o�<?����B��R�%��S�D�CHU���o��1"b�n
��t�)�ٶ�� �i:H���#4�D��CU�̝�$*�J=�z��\��v�o��@�Zm�{�j5�޽;��= �N�RW���m n�^�]�R�R)V�$��"�J�Fۿ�y�gL���|>�� ^g:�4��P(|��<�(n@�^(��U�lo��X������{ �[D�۝�����u�޽�s�lJz�u���U�VݸnݺC{#�Z���z�. /"o;q�=9X�)6"6�~��y4b����D�/L� �&�ω�i<v���m۶�P(l�%��P������t�$9�S�[������ Xe��Z���h��}��z�)s�1��i=����|���_��;��6mڴ�P(�#"� �"o�pW��`A�X��h��Z�vA\�����s,��B|��(D/����Xg:H'�(�զsP|��u6l���w�w��e˖�|߿ز�� ���x�|<�f{����&+��D仪�����O�?��b��U�@8;Ӆ������=�������s\�5�]i-Z4/��^��}�!:��\���w�ƍ#s����
,�4;o��5k�<GU/p�Ŧ�B�e�ԼF�qh��(%�AU���l~��G����ry��8 �1�Ku��X}�Qg��h��U�5�7o�n:�T��
���|�Y�fie�V�0�1�Ө�&^��,�����t��9���s�z����G�)U����h6����m�ކ�]���l��k��{��8��'m���:EZ�F��z��y�5d�������t� ��_
�ox���t�Nb��&��MǠ��'_�����߲��U� �zs������B��®]�vڶ}����A�����8γ |$��G���S�Eh���<����S�8�kT��L� 
�1�e}�t���t �/U���Qw�'���q�TzXD֫�� ��5�V����!�1�AU5������s�~m�����~ݰE�����"+B�헻�{��SU(
 �	����Q���dP����A ���fb[�R��tr��7    IDAT�(k�ڵg�J�u�Lf��\�����cզ)oY�O�91�UU�;���-BS�4M���H�Ї�=ϋ��d"�� Ǚ�B���|�t�N��- e�9(��7��C�N=��B�T�D�&��op.���\SU�բrm6�� ~����䋺�;,"o���a��bM:ERD�r��j��s�B�3"r��DaQշ
��L��0s���x;�����R�tn�m�f��2 +ǚ6U5z��4������E���VU}#�h�7E���i`A�ȉ�ݾm��qǎ��n�8�� ���D! �d:D'QUt��͞��j8h��r��K��e===Fv?ۍ}:��j�ͦc�[�.��=�B �i��J�)bA�H�ȇHUU�R�Tb3Ɣ�� �@���M����8�kL���e��Ӵ��w���J�R��o�X��k �@9�����zBIw]��� _3lY��)bA�H�������_1"��m�ϝS��\D�=�Tu�t�U�������߿f͚+ TF7|{��LA�ڱj�4V�_䋺��W�z]���(\c���p<������l�\��ss�|�2UM�� ���8ι �g:H�j: Ň�>�yޯL�[�TZ��Q���ȳ�Z|��f$�U�� �8��j�u��U�_�x񻺺�~`u���)�l6k:
M��	m�#N;�@�Px�����D&��?�J���I��>:M��\e:CX�;�<{�x4��np�D�����+遭��ر�@*�z����a��bM��"!c7��f�U�ͧV>�wD�ϝS'�۾}���t˖-� ���V����6"h/zы�]*�.ۼys���?��cզ#�>00�EU� 6׏��I���q��7���[�|�ɝ&CLG�TJ[��] ǚ�Bd�����n�!�l����h����3N�N䬳�ʎ��j���ȆoKL�j�o7� �
�S�zA���PՏ�za���*M������|�R�<d4�4�ر�r ���A�m�����I�(�D䛦3�V�T�����+H��h35<<lz�$L="rs�%�� b����1� :ez�FD>W.��n,���7��GM� �
U�d__�|�9�ϡ�d������1'�|������ �/���s���8x��a��7��uP�6���4>t2&w��t]��M���+W�Pկ���M�������p,�4�k6mڴ�t��k�ڵg���_e������N2�+
����cզ�GDw߶m�A���`��(L��ѱ���?Tu�m��Ӧp"�j6����Y��FD�tѢE�L�H*U�;M(.��'�tR�T*}����w���&"��3�+*Z��ժ��4_Dnqgm/V�T������t��(X���c5- �ڲeK�.8��{ ���AQ�f�Y>�˲b�yI��]׽�t�����u�J�sK����Tj#ǣ�4�+����׉c����8ΉA�X�\�VU?�k�Gݣ���.w�����^H��8/U�X����ŋ�5"�Tu��iߎ�DZ��J��e===.�u �`�Y�Z�z�tS�}������*��' �4��
��Vz&tj�|��y�?�0]���� �
�� ��q�l�b�!�HU�2��"�*�Ɯz��׬Ysa�m"��ٻ�8��2���TU/� 4�{�Ӊq��BwD�Q�q���2,.q��5㨃3��':��+QY5q7�%aIW'D[ۤSu�v6�$�RU�����L:��UunU}ޯW�B���!�^���<�ۣ�:Wԩ������!P!��b�;���M�B�ZH$�F�wD`�������4���U�f:���Xko �r������/z��ȓ�3Pd�2��mq����sٲe�
�U�il{4_QU��p׮]�P�ٮE@�Z�n���S�жm�v�GXZy��,Щj?��[k�AM�y�� ��ATCڌ1��:D��:���ru��N;����늮��_�HZU/0�U�����|~AOO�9{�����!�X,vgGGG�T/�= >9�H��Y�4&�: 5�|ӿ?�\���f%55�(">���q]C�"�$����ȭռ���e˖��Z{9� $�y�6�vc̪������RU�<�w�"iI�P��������N.��O���pv��UL>�G<G<��%��SU8�6� ����������&�d,(
�QO� 7�D��^&�y�7:�S�,[�����~k� ���y)zTuEKK���t�7�=�8O�R�S��\����t�[x�-����ʒ��8��=>��s<�=`���OV�P�~1��|@D����5�� ��CP�|����_ݲw���T��X,v��J%�WG��5��/�����H-Y��YU��f��g���?kkk{�Ν;�O�"A���_�' "�u|p�kKǈ\a�N�xj�pq��;�}�� �5�Լ���S�A�ȓ`�N�-���[�wvvv��% .0O$��LTXU�[DV�����������|�������+����,Yr^__ߤ��A�3��>'"�+g�J�Tw���N�x���5���y.�ՙ��z9���N�,U�����)��2�s���SDN)�u@�����W7o޼�ԓ�ɤo��p�b�9gxx�;"�\U'=-���m�]�^�e�W��Ø>}:����X�S�
gS�EdC5�5� 1�����Y���k���)anv�N�QT0��4Ջ�����<CD.��b������5|+�1����D]�y޷E�M�:�����t����"k�& ��֎S��a�N��v�@��X,v�T�p�������]� �'Ƙ���u�:Q�f`}"�l6;0��_��'���E����XĆT%{�� ��N�'�p,�J��ʖ�����y_�wNvI&������|���ʎS���6U�˩�"�����Nn>I��흪�1�9������G�0\�u���: �ůM���K�6577�ND.���o ߃�jPD��������S��ҥK�T��rk`�'��= >:�A�-����7�1WEp�{��#��˩�zC�vr�Ijkk��H$�nCT		c̻�t�։�^�(2%�v���z1���������Ū;=���P(|k˖-���|�����r]�Q�ȿ{���\.���^#�H�s�P8@���ʎSݫ�:����}���OV"���%�sձ�:::����w�é��^NE& _:���3�<s��������k��� p��~������X#�/�u�����y�\n�d����:�L��s"����W����Nm�"��ݻw�sq��J�R��'�9���1�|�� ��Ԫ��*G�iHU�?ҋ����Ƙ�U�- fpJlI���NDV͜9��֭��Dc�gUuF��߀��ܒJ���f�wL�a�M�Rר��Wn��^=,Щl\Nm�l6{���OF[[��x<~�U���,Ч�#��۹\�9���8�y###� "����5R�� �>����C���<�{��,��}P��~/�L�*�M��@ss������ 8���ʊSݫ�:�������\�|2DD<����]g!j��R��l6�v�VYk��bc����i�-[�k�� .�P)�0�ۦ�=�dtuu%D�ոW��i��I{{�+3�̶�����7����km@��_Nu��: ��S�"ri��-�}�] �u����Xk��:C-c����`[[ۮ���wvvn���	`9��= �ljjJ���7nܸ�Z�9 �ܹ� N���T����N8�ɜ��d~�?ʜ�"\���(���ѐJ��R���}�D"1�*�BCCCeJ41"��l6��Nn>I,xI,K��:Q�RU��St�4�d�c̤�pR�9sf�i�^��7����Ed��|e�ƍ��
��� �@�������s���F&z�����pV�c��T뇑�����+�SA�+�Ţ�#�4%����̟?�Ӯn>]]]�X,vX���j�y������e���iӖ����XU]+"�655-���^�8 U�2X�W�YCCC7�$���U�� ����|>��T�����\��1���鼋�O��ݻ���u�F����Ϫ�u���$���|M�ȥ2�6�ϔ�"��X,v��?��:�A��_$"���hD��d�7 >>�ss��oR���U�3�VV��^9A�Is��LU?2�^�fx�w��~�u����}�a������7 Ak+`c�U}��E�����ʈ�� ����JD>�yފɜ�� <T�Hew��;�G�iRS>�ᵮn>�dr�1�& 1�Y�� ��!j������y
Nsn(���0��9�x�M���7mڴ�u�q|�|�!��|��\.w�D�S�b2�|�1f3"�<�]�+�?qiRNm5ƼCU�.n>YƘOx��D���mmm|�:Ac���Շj�� ��U �J��'��髣\��R�� ��uBBD֌5ꛐ0� ��
d*;vu/?�4a.����'kpj�� ��Qt4555]�:D���--ijZZZ�5�įU]���tww�H���]:��K�6��W��.Q1OU�dɒY=1��}FD6T"T9q�{�q>M��o�_͚5�jW7��ŋ����_�D�������Vs/�:1`��TӧOw��� V��׺��{]�������<�y����M"��iP��6�L^66�}j{"W���G�iBNc)�������W���~@�u"�/�}�L�!j��r�A4777қ��p!�T:����s��� X�:���}l�'�a�����J*7Nu/�T2�]�?�F'7��T*u>��]� �#��u�Z#"Ϻ�@�� k��D� �����N���������D|������y�'z����G+���8ս|X�SI\~ө����ѫ��|�N8�㬵׹�ADG��������QKD�#����	MMM�cT�0�5Ƙszzz^���}U:�κ5U��_
�l�9h\""�X�`�K&rRoo行�@䇧]���T��V�e�w���������r�l�W" ���]��%���f̘�:B%� ����)�N�/ܸq��z�A�y�1��i�9�$3c�ؚd29�)*�l�~ _�P���T��k��E4y���}+�����擕�d�pR{{{���R op��XD����ˮCԐ!�������H$\�(��Ed5��vwwov�R�1�U��\砒��s-&�̪��郣���8�2����ۖ���,��Ӹ�'y&�}����!���A��ٳg/�־^D� ���mD�HUO�<�e�s���׹:=� 6��
 �����\������~7����Mh�ϭ[��@����Ot��i*"�r���;�ܼ�z{{G�0�-��^h�9�
�nGD�qO��I\}������Ƙ%�t�̞��U�t���^�,Y��{��(��DףAp+��T(RYq���@�#r��+�*W7��L&�T�� �2�,p���r���Q��E]]]5[�T��rP��}�G��3g.L��+7nܸ�u�j�(���A�6=�}���։�T,�`�2���Ot:,��TEc�;U��*@�d2�_A�������8�T�����"f��ݻ��u�Z����3Pe�X�������~:�>/�N�Y�n]Cͧ�<�e"�a�9h�N��>�U����9�}rX��a9����L&�Pӿ��t>�Apn,���[׹���r�{	D�#�u�F����-Ƙs���K����[�l��:�"7�\�3ꀪ�������9s��� OT(RYq��ı@�?��i�����wr�ؾ}�� ��`�1��*��T&�w^2�<�u��������U]1<<����璍7�u�5��>�����Aec �0���;4����
f*Nu�8�����D�}���O;1c]�W455%���3թ&c�D?
��קvn�	�Z '��鮞��U����\����O�o�sP�u477��DN�f�w��+��8�}bX��s8�ھ!��}���#n�֭�A��f�gc^
�j �s����\�:@`�^g����ҹݪ�Z H���+����\����@d�;Д����WM�X,�����/9սt,��?ݲ �T~�U&�y4���x��� ��7����}�$�!�LD�$��D`�< p��vQOO�9�tzM:�惠��}%�N�9�b�o�����"��lS��T0Sٸ��[K�P4�����e�ٴ� 5����� n�<�"�v op��dD5�" �|\�^_Z[[�;y+8��ƘU���w����-X��%�X��]砊[�H$���RO��OU/���
U.�|��Ϝ��t�|��3�X�*W7��\�7A�lii�U�BY��M�?�7נ����2�%���7n\����D$��n��:Uŕ�����|����ixx�Z�1"��0���v��U���;��#}}}# � X�L&_d�y�w `wj��$=�;����p�~���"�U�V�"�]U�.�No����y���u��8����+T��J6��{�w���S�lS��(��cDG	��bx�io����ھ�2@�
����Qu���D����z}�J�=� 6��
 ���W�8��d2y* Nmo<�y������ŮP��9qf|��hH�Rg��}�s8�7A��u�FqȨ�e �q��(��jii9alF
���� ���45ӧO�T�> � _K��[+q�F����R(� ^�:9��B���;v�)���W��
f���� ��:D9q�\���yuU��[<�8Q��+�!�*AD0mڴr^�xp{��3g����,�ˣP(|,�ټX,v�DN����L��P��@'W
�ڒ;TRyA0���n
��k� V��:Q�p��a���ո�ӧØ���{��|>����h�֭��鵵 �L���]� �D����g�z�Ν;w�HMl�FG���Pկ�a����a�9�MMMI +T�1י�\S��/^�x���ֻ5�3���C �c����yI:��z˖-����ttt�1�|���BΉ��"RrGGU�_ �
f�
c�N.�K$��:=�֭[� X��Rk�9"� �lR�j��u����r��͜9s����ꊖ���=Z�
�/H��A��r���Z��A���*��*�:��?�V-�TՆa�6��^("/p5�']�"�6�4�?Ţ�F��q��Lh�Dd�����t����g�����V*�J���ͮsP�|��+�	[�� HW0Ut�����ßu�J��f�A�2�{�z)�G\g"���;::�\���A�]%��ۃ߆��ۺ��WlڴiK��ј���E���9(��ZZZJ�nol��*��*�:U��~|Ϟ=|_c����s���A�b���rîsUX�P(��u��a�^�������4�!9 W��������V)���JXk�	��/�H����%��� n�`��TMO�a��!hj2�LO+��B +�F$T�8���X�נ#�y>`���~ѢE����͛7o�n2:h׮]��+\�Hk�	����g�a�NU#"+U�[�ԉm۶�
����?���F ��DT�MdĢ�@�1���H$�~�Qx����{zzn[�z5�:�J�^���sPM�����sJ=8�_�N�P�]�� "������A�N�� VX����i�����Ջ7��8��ͻk���VmPD���������s�-Z��xU��R�Jd�������%�����Uu9��Q�H�:U����=4�����b��@���]g"*��]�V�5���u�1fE>�Ovww�`q-"bFGGo�f�4/�}���(�lv��~�����X�S5ܕ��ֹAճ}��� V�����@�:�� �Ju�,�k���\��ӳj˖-�]�?���GD����D��'�.]:n��C�����l#Q�@���O��@n���=�5��bU��î3M���ֲ@����ܹ��yD������W��A5k����?�z����w �B�P�@�J�i6���ur+�N�s�ܚ N7Ɯ%"k �)�U}���\� �5@D6�a�-�9��:::ex�C    IDATZko��)4]�xq������O�}�P��@�JRc��]��h�d2��� ^�Zp�Ն���\�pMD�]Om���RT]�����8�u�yǎ��|�ԃ������V2�t����d2=�CP4A�� �(
\`��DD��7��A�8U�.g�E��|EUOu��ꃈ���<��㇇���
F�2`�N�bU�k��v�ر'�O���v �x�u&�#�����ѷ�a�mÉDb��tx��_�����Au�UDJ���{��}"rM%�Ա@��P�չ\n��T;����� �Z.�;�Z�z ݮ3=�1�v�:�u�D�z���g������A���W���T�ޚJ��zpss��Z�Hc�N�`c���A�IUm��Ap�XC���3b�� ��@�(U����|����|��� }UF��J=�����|���@����g2�G]��7�P�c�Y n�r��{��{0��1���{�uz�d2y,��8�u�_�zQ2�|q��'�k<U�H4,Щ�D�O�2��� γ�v� v'&W���uW�zd=�M�C�s���j���\g��3Ɣ<��u��A�I�"�:�����N��� �cNp��:�����Y�G���OU��0BD� ��鮳P�x���'�zpSS���Q�Hb�Nee����T�2�̣A\b�y�Q�j��F��lٲ͜9�b�9�O� �˭s�������uj(FD>Z��c��_�`�$�TNw�a��uj�L��A\""/�5��Uǜ������~�g�vuu-���SU��b��D�1
�۪E����/�sP�Q���l�\`_����@�r��� Ԙ��lo6��PDNf�Nՠ�u=ͽ���sٲe׍����ZD^@T��1�A��:�Q*�z �&$WDD�*�� ~/"_�`�����T*u����:�<�+\� �T*�LU?�a�yQ�=={���{{{G])��O>yn"�X."�p����!<��GĞ���%c�T)���ϱ����ujh*"��f�K9��<OD��ե[OA0�u�r�:���@tP6����lk�9 6��Cui����k]��*1��v�k���V755���p�✢EU?��<:�������9�'���R��r9�v%�İ@�r���r?w����0\���:U�B []��R���O?�t����Ý��[��w�@g����p�]d�2ï�Ax��rc�O Lw��h̹���Y���O�w#�:M�����]E��j.�[s��ǿ�
U��:������/Y�����kyWW�m�Ba;��]x�㭵(
������0��|�����PՂ�x��B ?0�u���D��a������a�t\�5�}`�������ے%Kf}\D� �:�6U=7��E�Mͩ��z�1� � p, ��?|Xka�}���� �n��]�  �L��1�H��Bt8"��l���bl���
G���[�w�j޵,Ω����=���_�� ��q$�aƘ� "W�wuu�.��h��'k����<��"
�
�ְg����:mmm���`qN6���~)A<�J�6��++���:M�>c�*�!�&clk��M&��c>`��LT{T��%K�4��������~����������b���p$���g�Y�!]2�<6�H��E���پ�*�{J9�X,^m��q�3�Qp:M��|-��<�:�T�ax��ٳ_�J {]硚3ghh�j�4�L���K=�����[Tu�1fC>������b����������C4:��1Ƭ�R�Y�JT�NK�x��Y�,�i��"�E�!�ʡ��w4�k���I8�쇨dc��+�;�R��o�}���8�g��"�tr�
�35]GG��9�!Ֆ�|�U)�5}�Re��ѰI\D�Z�8U�N.�{��D��y�%"�9 u�t�*f�����rOs
��kT�l9�J��T�ǹ\�|�9���� ���B4Q�zg.���R�M&�ӌ1j�=P�5��:M�1泮3UJ.��9�H���Y�&�>{�Y�p�	�����_
�] �?6B�⼱���\�hd�/���j����y�+J96�gU��
G�q�@��x(��v�ATI۶m��%���]��{�dN���X����T��b���� �K 5��:U��~z��%9�x��٣��,Ω�ȇJ=�Z{-�b��8X��dp�95�0o���K��5At$�HI;��R������-�B���U����*��`Y`P(���M�C���\g!*��S���R� `7wGX��D�iii���D�����t+T�� v��C�t��yg�Ŏ��������f \���ţr���OU߷s���U�)�Cq��8��!���	MŒиX�ӄ��W�E�U.���P(,UU>U��y�4w�T*����P(��� �Gʩ4w�r9>w���}�������BTfoJ�R�K90�{<R�<t,�i"
80͗�a�رcO.�;_U/��-:�ߋ�̟?F*��g��zU�^ o0�u8�) W�ш����Zk9rN�*���,"�V0t*��� ���\� ��\.w���@��,I��olnnΨ���:�&�B�r���,Z��xk�`C8�c��V���%� ��p$z�4_r�(J�0|<�˝�`�S����v���R�]�D��s4�����|>��\g!��fU}_)A0n9[u,ЩT���~�!��FUA\%"��u���jއ�n�:�:D#I&��B�p?����BT"��N8��c��_w��*�TU��:�_��Vd������N��ND4Y�ax������c�1� /p�����b�)��0p_���!X�S)���w\� ���[��r�q��Ө�<DTS,�+�0�z���
��z ��U������cN���It�@��R�����?�:Q-PU��y%�m��Q��R]�h��l��@IͲ����B��Β�=�{ vW8�a�NG��_w����d��tKK�)"��u"�6U�k��O�9E*�Z�. �]g!r�_��䴣���;
����!�:���AT������f�XNy'�#��Ƙ���-w���y��jU�����E�|c�;J9�s,š
c�N���q=��A��s����Qd�HDV��w2�<�u�z�J�^/"?0�u��`WWW�he2�mc���X��xF��<�>$*�L&��ǻ ��:Eګ�1ݾ�߼p��\����_�����:Q���w���R�+����ơ�?ܱc��9��E�ӹ\�� V(��CD�e \\,�|�����\�e���M ⮳E��~XD�h���� `��
c�NG��pD�7���j�[ O��CD�6��<�K{�w��0��������h</K&��9�A���� VW!OC�+:�����ݮCիl6�k�) v���"��"����/.^�x��0�@D$�J}��\g!�"�R�S�+��@��R�o�*;5UP�AKK�_cnv���"/�ݣ���y�W�z�F��Օ�<�fU�W�Y�j��|�?�h�r�<^�<�:��~�u�F���7��d.�>}z���_DD'�ȚT*���c\���d29m׮]��"�Y�j����K9PU9�PA,��p6�a�'cDU4cƌ��͛�X������Tu���&���\g�������X� �:Q-Rշ$�I�hǉ��`�ۊa�N�íՈ�lѢE?�����y�����:Ն6c̏|߿n���3\�q)�J-��ޫ��t����%�1�r��� ��B�����/_(��:Q�Y�zu�7�1�3g�O��:�pyss����3]�q����DU}�Q���Q�(����T�0��:=����{��Q,o �"�3f`����t"*�"k�=��_%"�����Ӭ��8�\"*ɬ|>�OG;�X,���*�i8��J���D�l޼����oii�ܹs�.��J���ݱhѢ�]��4���������U�r�ҥ㮷��Y �U)RCa�N����A��T��C��H$0o�<$	W����������<���E� ���BT��O?���v������hX�ӡ�A0�:Q#+
k <s��1�7oZ[[�"��Yk����A���2��}dl�+�\U��|�h?;�Ν� OU)R�`�N`�Y�:Q�۲e�~ ��^�5kfΜ�u�DT�8�O{���z��."�T*�U�oh�GD�s����w@oo�(�T)O�`�N�.�ͮs�� c�Gzmڴi�;w.��o"*����ttt,t�c���ڦ{��CU]�:Q�P�-�Ns/3��# ��|_U�s�q�� <v���Kg�8"���
�B����:�D-Z���D"q�s]g!j0�koo?q��0\`�Jyt Xk׸�@D$"7��z,üy����\�DDT���T*�V�AJ�J�����t��BԀ�Z{�x���*�i,�	 ��ax��D�G�X�& ��1�`��٘6�M���dͪz������~�睮�X�:Q�8�L�����~�ZaA�0Supz;Q�<��C� ��hǉfΜ�Y�fU!Ցz�������A���7��� �s������b�q{?�a��\���=����D%"Gl�|����7o���D�_(~�dɒH=��}�
�2˽%�"@Uߵt�Ҧq^W ?�b���wr�'��\� �?5cƌ� �Q��lGD���������""���� >�G%������w����Za��58���EӺu�
"�͉���p�1Ǡ�������3�H<���\X�dIs2��6���@DG&"�n�6����*ũk,���r:
Q�YkK��~��`Μ9hm��P"*�" ���R�o�������;E�վ7�FUOM�Rg��zAU\�L��zc���׹ADG����<8��D�f��̙3+���� �$��S�uÅv � ��o��(Tu�QtNs/������îC��&3�~дi�0{�l�H9#Q��g��;�JU|��T*��P(<�ŕ�����Tj�^�6m� �V1O]b���8��6���|��ɞ��҂�s��;�j���Y�"��sUu��_�{Q� �9ҋ}}}#"�*�K|�ָ
(a�e"r���wl94i��ND4GU�hoo�,��=�{������6U���m���3�9����N�@o\�s�;-Ո�Ls?�މh��Zk�������6jW��W �i!Qm����rɑ^����@ M����D�eӦM�x|��9��}ڴieHED�X k���։���M�<� ��<���k�{��m2��S &�ܖ��z���]g ��Q�[�q�̙3�ᝈJu�1��d2���ɩTjA"����ED.��K���k�9��h��zcz4�>�!�hb���M �����DD%��1?�}�DN�}�dU}@Ż�Q��ȿ���O���@o@���D5�G	����lii��y��ᝈJ�R ?I&�%���}���`R#�Di�-\���p/A�+ �*�|Gրb�XY��Q���������x�ܗ&��s�1�["2n�7��� p;�YՉEDUf���?�űfq4	,�ϐ�v��D49CCC��S���b1̝;�މ�x���ý "q�������L�zwY[[ۑ�K�:�I���sOC�C��������7+qmc�Ν����J\�����T���~�㎛�yޏ ��Q&"����D�͇{att�. �U�SX�7No'�qƘ�Os?ԬY�0}�������<�o`�---�Ǳ����8�'w�ܹ��U�RX�7k-׃ո���^U��=f̘��Dt4FDn�}��b��0�]"��{���'�Y[�0��zQ��a>�:M���P�{���`�ܹ��ND��f ǹBDUe�."�A���`-�I໮b���v��q+�g+}���&̙3�E:�G\ �����X,.��l6�>ҁanA��;��j ����N���A ?�ƽ�Q�Vկ���Ap����cG;A����	��aU�>�!��|T�����m؈���~ �xA.�{W����,"wU$Uc�� D�\.���DT>�6mZ`k��g���9s���|�cT�Zq����r��6�� �+� 's�x<~g�s�=��Z{��DT^z�����̞=---���&¥�DDD5�w >a�i�������S��؈{Y�5�c�� DT~�x�z �j�s�H��1��C�DDD�/ p���=��2��Se�6��O ��Plnn��u"*��z(�����{l "oWՂ����mp�X�k�0,�1\�>1l��6mݺu�u"��AU���}����|����� ,������h�Q�υa�-U��L�x<~O>���-�
G���ձ�������j;+��,Ή��j��l�־>�Sr��͕.�`۶m� �U�>��zc��u "�����QU�N����Q,/��}���hB,�����f���jP��վg�b�^�
����� �_���T�<� �m;Q4��R,�Ap^�
b�a?��@����ٳ�u"�����_�\���۷�{�E�~ �ZkAp����a�F�&����z�{�u "���q���Q<�lٛ����p���ApE���@A�`����z��]g ��hjj���J�g�^N�!""��~��|a���rO�t\�,��\�X�:Q�x��~/"?��=���ϩ�DDD����^���*��y�q�{	�z}���"�<k�"��J\�X,b�����4�HD6�ū]tc�
k���p|�h�/T�D��H�̦M����ĵ���U�ĥ���h|��"r���Ҧj```�}�sD�:f���v����M����0FFF�}Y"""�>����y�l��u��R�"��9��z�D�X,^�O���Z��pDDDյ�' ��^��qlt �X�ׯ�ٳg?�:U��͛���\�{��gam��}""":�� ��0��� ���@太5;�Z�$�~m���u���P�D�5S����{�Uރ >���~4�\�.%�n�3>��ׯ�� D�Nss��<=���۷��ለ�*��{�zFgA��z.�������r�#�X��)Ue�����T�Q(0<<\�DDDD4f/�U�zb�s�܃�U��p��8X�שX,������S9���DDDe��'�1�A���r�q�������l6�}�u"r���{cWW� /�蹣���V����<zT��0oUU.�f'�q�@�O[��OD  "7��g'z޾}�*����QX ?��^��Z�a�DU�E�u��������D 0��`BCᣣ����JDDDT��Xe�=1��X���\.�$��u��b�^�D�: ~��'U������s""�	{���0��t|[\�*Nq�C��ND�k�����s""�҉Ȧ�i�\_>��ED�u�#�X�ן�\.���D�-���m� �ю}��g���������Z��0p�Fq�8ŽΈ�c|zGD�Z�zu�7�v\>�g�v""�#pm<A�Y�O��<�:CT�@�?��Q��� ��������������l��Z� �+�����T�r��V lzs,�댪��u"��͛7����Gz�P(p������"��Z{N�A�*C�+U����aqz��:�����ýƵ�DDD������_
Ð[�U��lQ��]��u�Z����P(�I$� �u�筵v����(z �J$7����bu�Q�a�@�/��I���`�!�j0퐿�9�;m����EUg�H�h�U�� ����Q)���! �aj��"2������!��{���"����) ��bO
��bO��Zk�1�P(<�ǋ�l�U-�����b�lٲ���k5������0T�]�NDDT�FD������r�]�i@\�{,��K���.�2 =ы�w驼��Da "G��D����U�Cރ�����<�� {�s�<��"2���Ed�����"�WUEd������bO��}"����S| @�b��-��s    IDAT�Z��}hh�U"""v XU(��cǎ=��4���������5������-M��f��9��/,��y��?���BD`�}΃  <ੱ����O���?�I�m��S(v�a����_R�ڸq�]]]�x	 ����P�ΌDDT�Dd����0�m��۹s�n���p��,Q����:M���)�Rf�}�?������}?`��� {Tu�1f @�X,�Xl{;ǺiR�U�j��ለ����o��3��TG��<���t�#JX��c�c%��Ƒ �`��e��b��(��i����=�E$ �]DU� �M,{b���;\�P��b��
��'�����Q�q����NU�� |-����u:<U} �C�@�#�|�7%���/!",p֡}��������xBD�(��ijjz��Nk�C=���������9Ցa��X,�
�p��0T�'\���cdǎ����)�4Q� t�}@Ua�A�P(����(�U�u,{4��>Zb�BrDDn:�u""�2x����� �t�Jg�}��:F��@��-u�����9�$� ,�8�`�;���}�� ~%"���=a��Y�c׮]!��Q���Uwq`�6cw�!jX�׏R��CD8ŝ*m�?����{���}�@�cLOSSSw__߈ۨ�-�M��lp��ܚ�d�r���&��m�<o@��,Q��~�vǲ@' N���Z����g}�� �a A0��e��{��f�9���J�4������0��:���}��-����,��GI#�"b<��*��i ^1��/ �����t��km�1fC�ZF���%�6�9����aE�AU��Z��0�/h��m��}���W�A,��9E�lU}-�׎5���?�#�Zk7�a��JS���ه����HU��ȍ�b�Ɓ����<Ty���:C��@��X��tct�5�ұ�wc���n T�~c�� 6�]iD$�y�ߺ�ADDt�A ?���̆o�GU�9p�G,����L&�����xS��:�j�| o�7�*<�۟J�Q����---�mݺu�u�(�}���z��DD��Fܡ�kT�{��޸Tu+�?b�^����qtt4���MW�Wx�1���E��� �^U���{v�ر�u�(�֞�_�DD�P�[
�­��L ���9i�X�ׇ������%m�NT�b�/"���q���� �12�̯�FtCD�s������lR�5ƘՙLf��<-�bq�1Fp,�낈dK=�P(p�բ������}?�~��X,�k��s�Tj)�%�sQCx�U�5��z%Qc
��Y��v���D�:`�-�@��b	N!! x ެ�o6���]Ƙ�Tum����: յG�� J�a�8�� �`�^&2�^,9�Nt"r��.�|l�}��\���z���Z�W\NDDe�,�u"�b���0K~OJ�<� ��u�(`�^�1%ƘD%�Ց�X�9k�U���\.�8߄$��iƘ�\� "����NU];::��ݻw�s�j��d9�� �u�P(�\�[k9�N49X�."�����ݹ\�I������T�&�9�����p���-�?m��-T}�:�:CT�@�}������t��Y�r��M�R�Xk׉��###�EmDAU_�:Մ�- �Zk�N�6�����ס�D���j�ԃE���G��Ψ�"r*��777}�conN8�{��t�qF�DDt8E٢�w�+��߿s����CQ�a�>�z��	����&�$���b :tc>�k׮}�Tꡱ�k3�LO5�w�q3[ZZN��=��(���oP��"rW6����P��X��a�^�&�^��mֈ�o����k��!>�ݶ}�����LFss���"�ƴ_DQ���ڵƘA�Et�\.���"r44�5NUwN�xkm�#�D���C|�X�����p��ܝ���ʽ�OD�*����(ҶxPD*��RU��C�GU������u�X��8�5��11��E���KDV?����"r������p��2\�����Y٬�=������m۶M�!Q��`����Mt�"��i ^��� ��w�Ƚ���E�� &�NPD��S*�������1UMc��b�����E�Z����zJ��,Љj�|U]."�X��7c��S�T��v^u�Q� ���Z��X,>���T�Tu�KqY�׼X,6��R��'�]�����= n���<���O(���eGDy��=c���Y����v�!
X��8k턦�����:Qݘ�\ �c���� �BU>gΜ�{{{GE��qF""z��� ��w�3E���D�ڦ�g��3�s8ŝ�~��$����೩T� )ס��X?�GDd�����i�D�'"{�̚z��}oo��DN0�~�5�ic{�Q������y�\e�6��{NU�I:YH�S�T�,]	����:���QFq����������8#��Ό8�˼��Ό��D �����6�t�S�NHwg��|tC�R�9�T�s�+�$9��\Iw��<�y�033�xO�3�De)�OY�Y�[��� �A'"""�ƈ�<>{��&۶ojj����7i:Q#~��F���T������4�y^<�J=>00��t(��bAz����!"""z��<�q ��%�_���fc%Gkk���Ą�Ʊ�7�Jf�-��NDDD	5�w8�YqΊՇ���I�u��k:�I,荭��M∈�(���>+���>n���\�ת�GDG�XЩQ�j%K�9}NDDDqR�S ���� ��ܹ�OU��QyDd��v��az�,�r�QU>�NDDDqbOLL|`xxx�� DTUM��c���V�wp����b���%�3nDq!"c�3�Ƃ��XЉ��(�Dd��DT=Π��7� F+��;�Q��j��DT=Π��74�_�=�(�����Mg ��q��э�{C,�DDD+�e�`:UODX�M�ʉȁ
�aA'""�X�:Q<�*���@��,������:Qp��74�h��7r'"��ض P�g��t�x�`,�]������s���"#"hnnFKKR�,���o���"���0==���	v2BD8�N��Ƃ޸�[�n�*�&)���eYhooG[[�q��m���hmm�ܹs1>>����#�$%z�B�U�D̶�ɤ�`Ao\eϞ\�NDD���ֆ9s�<o��"���6���bll���ڱW�X1��� DT9U�4��4nנT����%�DDt$"���̝;��r~���͛W�XD�R�V���:,�,荬�� t"":���磥�%�1[[[YҩfXЉ:zê�t`f�{�Y����͛7MMM����҂9s�D26ѡT���&Q]���t ���T�`gЉ��P���hm�vⱭ�-� ��t��N�Y�M��T�K):j�ܹ5y.u���*��58Π��7���6���A����m�&�e�6g�)R"�쳙�b����U�M�3�DDtP؛�O�K�)��t "�NKK˴����7(UeA'"���H�g����k�z�,�b�3�D��X�T�E�X,��R�T�^��3�D��X�W��W��;�K��=��ץ�t�gYV����7�*��Wt~:Q=�&qD,���g�Uu<�,DD�xT�LR;E�����qU4����A'""�ڒ�[�PT������:###\�n: UL*��X,r���P(j>�m�5)9����d:Q�X���T����0gЉ� 01Q�}Ck�z�,"�u��qB"jh,�JU�� �95�j��-:EŲ,������W��BD��i,����Y\�NDD(��ͷ������s������DT����j:N,��7(U��//�� `�޽�?^,���H_��M�٭y޵jժf�Y��r���M�3�Ƃ޸8�NDDUSU���Fv욪bϞ=Ǝu�d��g�������fqD*�J���@���Y�A'"�gMMMadd$�}��si;E퐂 \�NԠ,�J�
���t""
����y�LOO�2^�P��O?�xD�b��ټ�-g�q�|SY��r�B�3�P��:��P(`Ϟ=ؿų骊}���g���9��a3�-�T���Q�,�bA7�*������:�����SOa߾}%����i�۷���U|�JV��b9��:,���Y�U��t"":� ��~�߿�m���	�mCD`Y� @(�����l9u�w�깧�~z磏>�7��*P,����[���7(i��vΠQ�jy^:Q%����J�R�_�!�
�7�3�*�&��Y&ΠQlLOO�
��N�`D$�K�Y���8NK%7�:�������122����e�̵kמj:�NU��`z���e�:v""""�T�����ݻ122����+�-[��t6"*�eYsMg0�Ϡ70Um�T��T�:������MNN�����N�up�eY�6�FDG��,�P���tE3�e���"""J@�� >�n?��A�?������6���f��ܤ�.qo`�3��7v"""����eݾk׮�L&�C�q.9餓:L#J:Πs��USйĝ���U�"�hjj���dR�� �q>��L�#JU������� ��&t"""��I��+ �²��������eݔ���פ��%���� T9YX�}MMM{
�B�q������� ^�g��ǹɲ�l۾����t8���g:�i,荭���Ϡ������G��x&��_U7��m:Q�$~���5��ܴcǎ1 A�Y������UU��E۶�p]w��Wuvv^����b:Q�K�:z��
�� �9Q��a˲n,
�d2��]��lgg�M#j@�M0�K�[�K�`�����(Lg�ϳ,닮�n�!�����n���4���-2�4��VMA�Z
"""":�������8��dP՛���OL�#�'����1��4��V�w P��<j�����f�ή۶��u��EUo�?��[�n�2�Ȥ����OX�]�3�"�t""""sVX-"�=8������\n3�]�J��v���UU��u�����.<;��ٝ�d�V�Aܒ��=��j�,�nA6�M���N�{��r�����>-QՋ \dY����UUo�ۧ����o: Q�,�Z�	D�Fg�޽{1��ro�:QC /�� �t:�.���3��o�,�~���g$
g�����D�DTP�+�������J��cY�g<��������ܨA�������e��g۶W(CDDDD����>11��u����=,����� 8�����7<����رc��8 ZB�DDDDD�8���eattt�u��03�~*��o```��D�#"�Mg�,�nv�{�TU]��� �HDDDDT?���;� (���[ �������|>�3�� :M�,�NU�Vq{,�DDDDIbx1��ȇE����� �pGGǣ\Op,�qP�w P��� """J���x/ ���\�}���mo��rO(� �����8N5������*]�>{/�3��R8d�=8�3��� 6�bY֣�\������8�2̬�H<���t ^hA����VD~��"�Ϧ�Q�Y�ͳ?0[���yLD� xTDU��y.{r�Hj�ҥm�^�`���>*!"'�,��KU�
��]�i��^�EdCwX�uG.�<���~ �j�و�(��9 ��قUp�OD~�OD��''''��m2,������������eu X��s��߇��"�q:f������[�K:��op,药�u�e �{�aR��ox:Ql��Uu�eYr���c,;�,�DD��������Ү�H��p]w@�'1S޽ vȧ��;v���ꈈd2���Ba��T*�^(ضݮ��"2?��"�`��,P� ��W��� ,˪4J___�d�s��Y,�1P,W������?�� BEDQ+ ؂�sm7�x�w���N�rc�Z���h�=�| kf@Uqp��B� �q
����W�!˲����U�,���V�۶�l��_,�r��^U��'Ie2���B�N�R� �,��PU)��g�Y0���� f��������"ݮ�� ����q�� �-����������a������� X�ͫg��ǀm� Tx�o �<�8D� �# �W��&''><<�������o]�}�KCMHDDT�f������#�<��S����u] ���� E c���_D�}&ZU�"r���X�*�)��#"����^3�6̜E?�q�g��������C�v+���HwTAz�jW��,�D��p���*"wz��LX��u�ʂNDDqs� /<�o^j�,�u^�kJU�*� X�g���@��7�!�j����%>G^���[�,�#"""
z�X�c@D*.��k>�Ad�v Tu����-�w��W���r�\׽�kk�zDDD���o/�b�u[,�0OCaA��j
�t��zFD6 �5��|��M�o�*:��	U-�zq�X\a�6�,�x�����y�uݝ N1�^���`���͛7�G���� ��BDDD�P��msy�!X��aβe˖��fU�("o;Q�����j��{L:��[�Ne2���'Mg!""��({wn��{,�1���|2��
�eYU���:O XoY�M�\��7wU�X�ʲ,t"""
��>^��At���cA�	U]�
o8�,D	q �� �����<���q]���q�DDD۶-�z���\,���m�~�P((x���l�̳�7�������7i:PH�,�DDDT��;v�,�D��A��Ǆ��\����#����x���p���,����?i:P�.]z�]��@�t"""j\�Z���8N��qĂՖ�{B�(��;� �)�N����?b:P�z{{�3�̿��?��BDDD�KD��s}&�YAkTyz|�@D,U*��. 3QyTUopS>���Gk||�������0�����VY=�F�Q���G���� �Jn�m��b�r$��U�Uu���$�K��1<<��u�o �s�Y����1�H�K�_� ��z���
��;v���[ ����n����t:}����w�To� ��eY�H��BDDDgrɒ%�-�Ue�8z�ض}2���/"w�	��3"rG7MMM�x����L�g�|�s]�Z �5�������<���;]�m\�~�	�`u���%"	+�!� ~�G��߫�|v��e�C�Lg!""��Q��X�Â#"RUA/
�H��<��'"?*���2����e``�	�u���Lg!""��R�q��.�$�,�=^^R��CCC�]������E)৖e]����W�0�+ �!�=����JW��/�,.�;�D�e��8N5����
C�m ��5��uy�w����},���<�w �m:5�,�rn�m��Q�id����e�~C��_��(y ?�LymA�e�@��,DDDT�v�)��#�z�T���� <R�J�pMo�}g�k/��� |�t"""j�ʽAUO�"H�cA��j7�Sբ��V�2���uA����c��y������Z0,�D��0������^Y]D��eih\�?U�Y� �(�q��gZD~�5"rS.�7�~/����{%�/��BDDD�˲��
��+Uu^Tyz̨�EĮ��g۶o)
<n����������o߾�t:�T���
�A����>
�Gʹ^U���Qp�{��d2�V3@��������xTu��|YUO�<�T��d9������DDDT����Se���Ϗ�=���bO�c��ad�ěp���[�l����>��~Ygd�y����/L� ""��T�q��G�%�1$"= ��fU�AD��)UDU��"r��y>�A�    IDAT< T�S"��6�����ꇪ����3�14[Ы2;˹=�8�S����>�ϟ���WX�����GE�Ǯ�s��A\ww�| +#���X�cHU���WG�ȍa���py�Ppr�ܺ|>����S�i�9����~LOOo.�� ր�Q���S[&�9���2��'ÉD13-"?	��|>y2�ȫ 4��ADDDu#�s���rnPյQ������(���������<��pRQ��?A�s>�ϙC�����R(��	�Y������}򓪮�"H\p�{L����E��0�PcS� .O�R��.c9O��˗��P(<�s""":����bA?Π�T}�O �?����<��������E�a��ǹĶ��n:՟rwpw���Q���R��E$���j�inn�����(����Q�S 7A��|��a��N:餎�����w��BD�OU!�����(�N��A�eYYn]tl\�_��^� }}}�"rC�����9��XΓ�uݵSSS�YΉ(,,�D�;�o߾��{Ί*O\��ǘ���8׆1�/� �\.��\.��t�=�u/px6)߃���Ϗ�=�T��a��t������ci���,�˽��M�!3V�\��q�[ |@�t"""j�s��X �e���Pf�{{{��4���n<dY�+g�yY_\)^2�����ӏx��,DDD�PʚA���|	���q���[�q'��,��2�xȩ��}�����}�Ð9�V�jv]���z�e��QC�J�ӏ�s���2�0q�̢�r�;�c,2�̜c~���W+��L4�uWMLL��g��DDDT�G���'ʹAU_U�8����,+���U�("?c,��) _K�R'y�we�_H)~\�};���a:5��7�����k'�ٱ��ƣ�]�J�>��߿�t2oժU�_�	�Y����ᕵ�pww�
 nA�3��wFggg[����0ƢH�VD��y�E,�<���A��Ql��e9�
�s��7,������ ~�X� �wtt�4���j:��u߁�O�O7���b�N���fv�ر������t,��pnXA����O �����S<ϻr�֭S��y���-��~3��7����KUo�}�|���,D=U-��sU��%bAO 	��> ` ��jU���]244�]�	 �8�ɅB�Kډ(r��k۶�PU������|�t&"��C�\��B /�(K찠'��ŋ�c ��e����I��_��~ٟbR|���Ny�i��Q��N�Ro�̼GX�dɇ �b8E����炽�d��J�Tkkkh������� �)
�x����}��n��� p=��y�(�&T�m�?����;��D�~S��(RAkkko97���
G,�	���-s�}#�ma�G%{\D^�y�%;w�6��Ggg�) ~	����Q"������G��9����B O�8E�񾾾�rn�2��'Gh]U�w���k�ZZZzr�ܽ��P}q]���e��Kډ�v>����|�:�7��(�FY矻��	�䈲�zr��jժya�J��������R�ԋ=ϻ���o�t����~�9��Q2��U���c)���y�y ��)QL�jY�E"�����zr����C;ޠ�������KUw��:��.���&zVgg���Fp�v"�!U��󼏕s��y}"� �"�ED5�J��)�z>^>����kB� ��u������Lg����d.�,�A �Mg!�D�������Z,��\.�QU/��`D��?|c����mR��'������Z�<M����r�u�|�)�a���H�u�/��O�]ډ���J�RV���wx��>Ս_�sqWWש :��_,��rʊ+�����oLUok�S _���xa.���t�?'�x�b�qn�Y b:%�����OT;��y?������(ky{��*H���'�쎪����/�����<ϻtxxx��0T2��+S�� �&GD��+ o
��S.�� �xDT;A�U���ݤ`AOU}C������0�L���MOO����]��P}r]�êz�Mg!���2==}��yτ=��y�W�{\"������'K��u�V ��.N|��'�y�V�jk0U-����/!��=ϻlhhh��0T�,Y2'��\�* i�y�(q�,�ܡ��ȎG����_Q�OD��_�j9G,��-�<qƂ�<����g�9�eY��x16�ʎ��5�\n��0T�:;;Oinn~PUי�BD�toKK���D�"����_*"<���1����"I� ,�	$"�.s��r[l	s�z�X,��y��[�n�2��S&�y�eY8�t"J�_LNN�A__�X-^LU����{/�[j�zDT9U���5�Lo
{@��Gv ���jpp�צ�P}�jDTnN�Roڽ{��Z��֭[�� x�{k��DT�g|��ԋ�/_�" 'E�'�XГ����+�0�J}3�����4��TU��JG��d������FDTs"��K��=���*���455] "�M�>�=��zq*�zs�a�=�
��[�o��� ��� �O����y�3��W&�y�����+Lg!�DR _�<�����&�l۶mtzz�� ~c2=_���U5�պI�P"rac�Lt�۶W{���2w��q]�2U� �FDf |��+����Ν;�U�����t"�=۶K.�V������zB��N:�P�u�m� ���� &0��kw���o:կU�V�s�z _�P#"3�x��y_7�p���"�z C�� `,��=Z�����o �a��cAO�����P���>���0�l������9��/���x �;Lg!����U�����鳏����~�OTO�+��-��T�=�� }�;�oD0f�*`�\s��y���o�<B���y@D����GL9��~� ���B�pw�z�U��E��W�=�D�M�W�u	��y���u�	y9�5��}��� n0�t"J��wtt����M)U>�@U/0i:QR�jɛ@����`^�q�=�:�����U��
{�:� ���\.��"�
˖-kw� �~�%"3&|��K�e����w�G���T>��ԋE��Q�I
�aL�(��7773G���쮲��<��|>�����N7�N��]��Qb� ^�y�7M�F.�����	���a&�P�Z���"b� �<���No�P�l۶mTD�s�:p����K=���� T�\�}�eY� zLg!�ĺ�P(��y�C������k |�t�$��^��+ ,�0Nb��Sg&�9;�qc��]Uw�ȅ��]2<<��t���|��7)"2�������;w�6&L��}MU?m:QRAPrAWU��tB��3����7a�[K"r�Ss�܍��P�����OD��6�'�T�t"�� x����c?}��2�+L� J�����e\��Ȓ$:���^�>�[�Yc ޗ��������0T�\�]�8�m >f:K҉��DF��u�T��|>��,Q�<���w�sř��^굙Lf���$
:����2�A���� L�=n�~iY���}�tj��� ��BD��WU/��r����GL����?���b:Q\�s���D$�X�	 ���/s߾}�. 7�=nD
 ����+��C�!�ɼADp��,D�<"�����f7PK�|>�� ��t�ڟJ�~Qʅ"bE�#���  "r�����A�D��eY/�<>�G�s�S�z3����Q�����w���o:�)����\D��t��������gW�vF�'QX��ŝ���
{�|>�|��DE�?� ��d:5�l6�v]�"�/�fpDT{7��j��������)�o��B#%���wG$�X��Y�e��<EU����a��ay[.��h>�?`:5�%K��ٵk� >h:%���R��{�wA�;+���L�G|�t�P���E$����ǂN�R�wf��t�~@=-�MDN��iT�L&�����^ o2����("�)"/�}�j�aꕪ}߿DU�5������r��R.t�< K"Γ8,�t�v��z������>����O����R����/U��n:%�� ���r�<��aꝪ�-[�>U��D�+gy;wo� :=���/�q��b�2lp��y_�3{T�L&s>�{���Qb���}���y��Hz{{�[[[���t�FdY�M�\���ݢ�F�'�X��ptuu-{�|>�3 a�[𵖖���y�x}j`��~pv��y��Q"L�����}߿�(W���o���i:Q��r���R.,
o�q�DbA��5ApQ؃�j "�{��T��<ϻl��5QIDD\��fv��A"�é�թT���.�k:O��<o<� �m:Q�P�����G�%�X��y�Z�n��7LG1�ܖJ�z|���T����Ϙ�BDɡ������0�#N��������x�t�q})�\�r)�7D�%�X��yD��L椰�����>�q3�ٍ�f_��d�V�jv�Z ���,T_��4D�t�1˲�u'}}}c�T�"RҲ]����|If
����'���NG"���H�r��ߨ�˸Ubɒ%s&''o�N�Y����ϟ������t��7g2��C�Q��mۯ��t�z%"ח��YU/�:O����ѼO"�.�<�v }a���������F06��ʕ+�677ߣ���B�����e!�J����-bQ�(��zČfJz*�:3G��a��bI��3�� /�8N����ќ��9a:����8��?�<���!�K	��ݽbzz�^ g��B�����9??X�/^���vX��Rh>Ň�4���Ĳ�7�5�����,�BU}�a���*�X>Š�B�1�x�H�R�y���Ƣ���zq�Px �*�Y�>577#�:�F��eaΜ9X�h�̙۶k��b�$�q^e:D��ijj:�8��P�S��x�^��	�� O����Q��EQ���s��a ?�b�K���;�R��/_�� 6 8�t�_���ǽƲ,���cѢE�?>���j��b���El۶m�MMMo PҌ!Q\S�E###8!�,�ǂN���E4��Ux_^U_�y�e����:��b�q��l۾,�t�m������E���X�`N8�.�J�+���fK���N���_�r��| �0ĂN���(�<�!����T*���]Qd�dp�t� `��,T����mcΜ9X�x1:::8�N�hU�w��۶m���>�ݦ��""�.������#�C`A��{��n���/���/��>�6�jtvv�9[ι<��ɲ����������Yu>�N�PU.s������---op��,DLA��R.�m�R �V,�t\��,zss�� �2ϲ�s=ϻ���+���uݵ�e�`��,T�����fڶm���'�p-Z�����n@G�����ɓ%j���o,�7�����z���>�E"�R�?�A:��=�/���}}}� ��h�/"�U�������~mJ�q^�6 �Mg��������T���.\���vά�sX��'�3$I>�?�N��
�f�Y�jED�Y�u���o�<�84��J1���%�#���(�� _�<�m�|�Gt,�Ϝ���tjMMM5-��ts��98�>����d*�z 7�L��uvvV�����b�ҥop��,D5��y��r�eY�F�~��J��( p�!��S�WqI;��uݗ�>s���da={^�g \'"�3g�����7�������ԴXUש� p����,��C$Moo����.u�,�F��_VU=�u��@U_W�L4��Q�z�y�����`�� ?�,�O�D��0��p+��9���,�����D�� n�����m۶��n����V��sD� ���Z%�.�]�!�FU�"򁮮��b��.�y�"��P(�t�9fNt
wS:&)���L&�JU��t�����y���."�8�Ş��M����3cY�= �Lg����ގ9s�D1���U�aӦM�U;��8���ZD^	`������bFD^��嶚ΑD"b�Z�����q�_Bqs��y��իW7���z �� S��x���t�0q������?�����5,�
�q˲��9�ID�^�^� ���b�Ǐ<�H_�����c�k�w �ͦ���N�,�U=CU��� ���'Վ�~�'L�H"U���Z������7�(,� J:�xtt�"�w9�%t*GS�P�0��5��H�-[�$�J�`��,�xB�� �;Uu}�P��-[v��$������?����8'��� V�� ���h�,[��/����(��̙3�-��޽{M�!����$���J���o�T��d��8��D&uww�O��?�"�Y�1��U�a�S�z�������ٖ-[�H�n��7��9��lz׮]+ �$"˂ X."KUu��,�̬�rp޴�t:� %�D�z�G���즶��˲0::j:Q��T�E���g[��6�0�|,�T�w��� ךBtPggg�eY78�tjL�m����Ƿ��ɲ�����뮻
E����G,����n	��3�!��j��.�<�V>tcD仪�������(��5���r��R.�m�2�=7�����:ՉիW7Y��c g��B�����'D� �oڴiSԙ�E��	 Ϟ����y�eY,�sz&�Y���6��D�� ��nnnƂ022� �i��X,���R�s]� �y4��\�l"r��8���A$"����w ��tjlG9Z� �~ �,
Noo�7n�"I��h,��o5����ΐT���;U���?O��X�`�5�;�+�B��t�y�(8�N�,� ��tJ�����CU/2��[kk�o���KD�S�z{{�����Dx,n�]��������=ǿ�"�] ��I*���g��E���J��W�u���p�q���UDU/���tM��r��|�tj|���{T�U}��������6n�x5��щg�k�5����T�t�� ��5۶�p�B�Ӝh������w�x�{,�2:U*mY��2���uݏ��tj|"���c�-ڴi�%�6mZ�u��)ә�����#|��1 7��ea��G{L��^��R.������q��S5>r�I'u�A���{|�t�U�'�6�e�f�i +M�H"y��8�2�#��w�_ttt�����y�J����[J��q�7 xI�y�8XЩ�&''��tJ�L&s!���$
������p���ܹs%�y�I�,ΐ����x�h�?g�̛7\�@�DU�����w�a�$,�T���l
Q�\�=KU�nnI�z����L�h4�m�b:C½s�ʕKM�H��G`~|�kZ[[�����N��N���(��L&������S��ݻw��t�7�u_ `=���&*��\e:C#RUt�����?`:D�w�Mss3.\�c��8U�\�r��N�+UMU��t��+V����Xl:��ݹ\n���ݼ���m:Dmڴ�n ��K�RX�h���j����T�F��Yʵ]]]+�=�HT"t
C��8\C�[�x��b�x���0���ED��t�F�����8���C$�� ~Pʵ�ea����<�LP �/���s~�W'X�)�e���/�W�njii�	�3Lg���=o޼��ѨD��>p�8CD���%E����j���?Zʅ˖-[���D�JǂN�P��:;;�6���ADdll� ^g:���<�2]]]��M��[�/_�e:Dmܸ� ��sOkk+�K�Z�F��MMM��]*�JPh,���(��?ͥ����6��Q�EΞ�۶mujNI���N��p�B�R<��"�u���J�p���sU�#Q��S������c:5�L&�Q n:�ֽ����6����ח�^����`Y��0�oYl�ƢE����CI({����)�����Xa� :�JU?k:5.�uߡ���t�/U����̲,��r����;M�H��~x;��*��ܹ</�B����}��]�\�l��X�    IDATٲv�dԙ�|,�*U}g&�Ym:5���W�_�(:��z����;��U���	V�fqG����%����~�ԋ�����=E��Sج٣�J��ݽ�X,��g�P��������X����3���!�(� (T3F*�����R*J*U��R��-[����"�DbA�(\��*�!�1�Z�j^�P�QD���B������D�p��tD3 �6o�<,"�GD�����ب����kJ�8�N���PX�)
6��M�����f�����x��,{��|��!Y&�Y��|uHU߽r�J~�iFU��u�(6۶��BD>��A)��Ξ�Yđ�
,���wvvr)$��ݻ�&"�7��⏛�U/~M�_ͅBღC$���ԏ�k��G�577�5$���r��m�^����p�����STl˲>g:�/�q��goR��omm�������7U��l6�6�#i�lٲ_Dn
sL˲0�|̛7�����LA��R/���nQՒ�'3X�)Jwuu�j:��q.����$���\���7f:G��kuo�����L�H�Ж����w��N��|>��R/.��<�<t���L�����dֈȷ��?T#A|�t�8�z��f�����(�>��{[[[�SS�]MMM_��K�,�Ó�� S����_�+Vt��M �N�je ���m:DL�l: �+�9�t�����V��_D0w�\tttp�;�o۶m�ԋ���?>{�X�)j���7��s]wa�X���@���Rw��������"�eY<�� U�d���ZZZp�	' ��V�_�s�Zgg�	 >a
:��y��dƺu��5kּ&�Jm�%�TK*"%����K��+p���{\��4�#iy�{��u,��w
D�����`��_�a&
:Մ��_��v�>��֞��֬Ys����GGG�*
]�sQ�ܝ�嶙"r��T�4OȨ=���Z��ܹs�`�X��'��r��R/���tU��Q�p�_5��k3��L���d��֬YsI6�����԰�ܨ�޷oߒ��q��(�D��Åg�� T:������j���PMMM�����uɨ�T*�7��`Y���D��"��N5��_������:�;��^���s;����m h���	�߿�hFJ�����?2".T���,L�R�5"i6o޼��Z���`�' ��}�|m2�o����J��u�U �a� V�Zzigg�� pV���]��TU�HU���w������hɛ��JU8<<��t�aAo0"�i�7I�-U����]�_v�ҥKG�z꩗��� 8�ƯO���ҥK���D���j��=˲`�6���MG�+�ͤ��������&dݺuv6�='��~5���Al�ݙ��h��E����0%�sqy{�X��Ɏ��t��Q��(y�]�cǎ~��_� �2P�D�ӽ��%7Y�u�RՋ��TAKK�<t��N˲>n:�i������sAOO��۷o�� >�;A�={� 8iC������q1�h�
�9�|"�#�jl�����K/�g�u�"U-x�w���VUw�A��q.����T��Pǧo455��m�1�:�p��8�L���:��3�n�>�N?#"7��� t�3���(�E~pO��w�9~��m����f�9�|�z��8��Α@5�,nVS�Px����r�{&''_
��03�O��m��˹�q�u"rNT��e�6���LǨ[,�d�|˲>g:k׮]��f/�f��Y��kv��� ���޽{155nH�2ٶ���Ĳ,.ool���4�ǭ���Z��П��<�Ry�|��Ph��cǎ�w�_�zu��}����M叅��P�?u]��s$��X====k֬�"���:�m ���rԁp���PrUa�����Cĉ���70�8��,7�#I6o�<�v/�����e�Ῐ��nU��T�Z��:A|�����>�n�c777ò~_A����X�ɔ��t/.�=�ܖ�kמ��f�����H��&o/�5����oOw!�f7h�A���ؚU���5V�3�gY�B��G�����}�ݪ���5�E����|ɳ��,Rտ�2S5R�������Q�u���t�8:��f�ًzzz�޻w�� n��&o'��Z�B###���A "?4"n8����o:D�
���̹��7}߿.�N���7�*U�g�\�rn�+ ����fngR
��z<��+"�-Cp�gv���|8�ͮ������M��F������Q�s�<��s��cAo|�
�¥�C$ɖ-[�Xo��X�v�Ǻ`���|߿PU�`o�rQy�R���sCgg�) ���yKK�s�����O)AT�7e8����C4��kמ��f?;��[��\��M��Q���bdd�B!�"*	��G�$��z������{g���#�#.s?���W�ŗ �+�HT&�������cY�?���*�J��N�e��Ă� "R��@D��y�Zi֭[gg��s������Al�E���[��c;ՙ���沖��-^�x.�L����B��^�9�DDn𔁗�XJ\29888����03�?�XT�_-Y��k�ܐ�d���M��cNr��'�� u��d���������n���`͚5Wm߾=�^ ���T���q����zy��Q��m�6j:G�477s�<^>#"u� �z{{�\g�W�q�/+�bUU��^,� �a.:�@U/���S�իW7��F�����|Ķ�5�_��7i���/1�^�u�Y�֬YsI6������n�QU?`��lSSS3��9L-%�;n;';��6�!���&˲�S�=�����}�l ��9T�*��Y�=###��"U�����A>��cR �l:�Ig�uVw6�������b�8���p�9��T,1:�IJ�;#,��t���z�\n:@�lڴ�~ ;����=��T�7�j��+d<~,:U�e�vYG�9���_D���[�NGǂ�`�������u�L�B�!ji�ڵ��Y��l6�[,�cfW��0�E]	� ###��t��P՟nݺ��=P�n�(tk\�}��I�3Ӄ?0�ҋ���Ϋ�f��~�J�^�J ��b��X������=e��O����C���r�z�ꪝQ��������e˖����C6y�j6��� ت���c:۱�*��Ƹc;�%1�g"�g��.g��*�k��1�D?����	��.�,�5 ~J":"U�=��}��{�����uQe�FSSl��S�����X�β�z[�I�ӟ3"L�l����炞����o��4f6y� �p���۷����c�HGG��!bl�� �7��{��I�y��' ��֯+"�8�Ӫ����K����L���˹AD� �5>���e���gٟ�=a��)U9�r�ȟuuu�j:D5�<��ų�������(���w�arTe���oU�e&7n�vUO&q%��L����
(
Y]����\o����sUXQ�uUv�"  w��P � Xu$�骆I�:������c�1��L�tu�S]��y��'�>��L��[�=�� ��֬b���{���!Ĥ���}&�irT�m�Q�#@�fq�,�
��-�uG]�=����D�)��
�?4�۶?��&Z�ɺs�A))�cf��TD�ۮ�j���F���őG������������2���I ���6�\.˦pBk���>��� �J�l6ۯ:D�\@�&.-�����y.\��p�N�A�c*��r3/�f�K |�MyZ�H$t��$)�c��S*�4�*҉�X�qޣ:�T��X�jժ�Mޞ�}�I 8�5�Z�bǎ�c1ioo�J��U�A�3Zu����ry �=.�i͚5���\�<���j"��{�3���ZC���;2u�%�L
�����D�Vwf�(���:Ǿ�?����GyB�%�V��(7���+Tg3ˎ�B{Dt����3K�����8�vm�LE�{������Ʈ��v��GAf�g����<�gͼ�q�S��M�Z"G�G
����k\�#4㋪Cv�a������jժ�w�޽����`|��Ū�����.���}ioo#)�c����s���%�������}_��t"Z`]���@ϔJ�O6�����pi��$�N�vts��W2f�ۈA������d�{Е+W��Z�����;��� 7Nl�67�,aA�XTC����o��~�:D'3C6��f>-�ͮP�#~��_?��a��̯9�#��s�|>���1>�.ǾL��>4<<���פ�����' ���D"�:FG�=f�O$�,+�41ø�����}3Gy�����Nl�6HD�a|���|�J%�����!D#����bf)���`��T��"R��N�e���lf�L�M_���/�����74�?Ц<36�]�_Lvq))�c�ы �J�ԪrH�\|#��kך�������_������7� ��[�*�
v��!�"��N�b@
��xG&�y��q�̷أ`ܶ������<�x g���/����j�Dd��>EMЬ^���2C�Vw":/��l�>��U�V��z���6m�T �+ �8��V�N�s"���1У:��IDZ��ir��^"�M�ЯZ�zuhK��w]�r�0p_X�ꎙ�-
n3�q�#̼�]�fʲ,imo)�E]�e��� pUӟk֬9p���g����X*����|���ǌ��;w�Z���!D�~944�]u�N�bŊ$��s���Z۶W�#&�W4�;�phhh��y�����;4�B�py3/�m�`f��
4SA������KI�3�^���x��-[>��_\�fMo�9�V��I�Zf� �`v{#FϞ={06&����`fioo��{n1�!n���Cu�8�={��l	{\f~)8����u��M�<@SǊu�������_KD}@Ws�H*�
��'�N�҆��S�pW��/Y�d�3Ǐ<��CW�^}~�Z�np1� @�6 ��E�ND�@u�Ng���ov�8�!:�}��W!��������85�7o�<�f~�gU�P�s�B�ͼ���xm���X"���]f�_J
1���r��:
 �L��&���6mz5�g�����Y�\Ʈ]�T��Y���;�:D�#�Ū35��? �Fu�NGD�1s�rOl�@���3>�zٲe?*��_p��,!zl�_i�K�.��]GK;&�H���t��vi<�C�ͦM����&o��M�};w�DE��)�㋈��f�oP��ӭ[��7 �v&��mӦM[\�=��O�ԦiS1�s�\ó\DD��_�e����[��^������ނ�"###k���<�9�J6�Q����!�}_
�c�/�X�'��D�b�����D�N����� .�����hhhh}3/p���|B��T"�h���R����a�i"�L��`�b޵k�\�3�k�.�J%�1����O=��C�CĄ�A��U�m�Mu�N����*��L�F�r]���_�	�y4 ��ؗ,Y����)ό���ey�RR��L��N��R	����cD���|�D������"Z�:�P�:�Bw���������+Vh�>](~�p���� ���03��u݆o���,˺��6暑v����d�K�Qi��qquu�s���ݻQ�TTǈ�ND�Tu��t���������:�����:Y�����re�u/$�~ ��3SDt��yM�βm�C:��'�I���:F�H�3A<�jg��LH�9=���}�vy�!"�Z����\�@ ��d2�������w�`�nm�/���7z�w4���V��IC����h�Gk��n��V��q!�������e�ٳGuU<@D���3Ϭgf9VQD�S�B���C�Y T�Cha?"jj�hΣ�>Z`�_)���zի(�a�̮�^ND� �Mu�1��m۶�*�e��U �iQ����q"�����.m6vػw�.紫6
�.f>۲�L.�;vxxx)3�RL�V�OTg�����!�b��8�_����T��[�D��
�mZ>��u�S�y-����L���|�Gͼ�q��Xݦ<3�ӾSq#_��	r#"�]���,3_`m�X\���N^�~��>��۶��>��h�����<$�Je��B+&��U��d�r�&��M�6��<�&��p��,u���tS��L�hf>�]�fJ����H
��	z�;�L��Lę�T*qjup�a'Ι3g�������r7mܸ��/��8k��r���}��3˚c�b��f���ѩ~���ng�f]r�G�T��3V(�q]�L ��Ӳ'p���@�#-Z�h�a���C0mQh��1�X����M;.�t:���-.��{�"�Lv�O�M��߹~���S��e˖-p3���B�����y��q���|I胙������������� ���L�|4ܜl:��������J�rƏeS}�s��?l��D�R }m�3ca�������hY�O��k�.�~���C� >bY����]�n����Dd�����CI)D�ݯ:@�����򱱱��ѩ�Ν{;��
�>C���,��{>�� �򔏂eY�l��l�� ��Myf�4M$����arOGR��@X��M����عsgT/�� �"��T�Ճr�ܱ�\�|���C۶�
��E"t�'�aH�.&�̟�8J���+�]�Я����&���x�w3���
"�opppG�ٶm���hg��P1��{���]&�NkӪR*��w�^�1����a�Sv��y@.�;yݺuW?��#��8��. jCF!T�=D�]L!e��7I�_���U��Dl���03{�wu"�{�+]׽�ѿLD]��L�ӡ��.%��c�St"BWW�6������d��:M��. 7�_�����rO�mۯ�M�D�<��T��)��T��m� \�:H�Y�|���6m�`a�C�-�k�"�M|�δm���[ n�pO�����8�=qfNU'�̠ONf�c���N�20�N��>��D�9f~e.�[������r���q��� ݭGB+똹�:D�h7�#������E�Ct�o��
�FCgW�\y��q����|�?����wx�����F_�8�qD��6di�ʽ�d}rR���%���[d�V�ص��/�Vd�{|��}'���Ol��l  �`Y��+�&��=|�T�ۿ\.���m��͝�"���b�Ba�뺟�
������im_�x�|��ԯՑj��%��L�iG�*Jt�vu/�k���":�\.�~��s��%6lx�]ڶ}�7����PL
���V@菈�&�ɜ�:G�ٰa�C �T0��+V�У2`�����c0�GO;��ņO4 "2M�
 K;P�DB�M�şI�.�B�Vw ؽ{7��r��>OD�3�)�bq�����\�n��{챑vXc��i ��ѱ�y��14Wu �a\�hѢ�st�RT1�~`*��+ㆂ�}�u�nY�!hm9��o۶mw�/p�D���""�R�����G&�mR�*��g�33v�څ8 �6�' �	����?�
ztl�>��� xD�z�󼆏���:����D�[ ަ:H���g�t����������0�3��f�5ul 3_�y�/����	����CWW��ה̠��ҩսR����
� 癦��\.wh.�;ob��Ћ��&�[!3]���Vu���wьS'����r��A��oY�bE,��u�hѢW8@���������1�9 � �i)��L&a������I�3a_�����f��p3�mYV&�����.|衇��ƈI��Wx��B���T�����4�����L&�U�èhs�N�RoU0��\���D������ �q]��M������Ř�3CZ�5'-�1���%�J�Z��Z��>�dv��˲�=8x���&�;���=7n�v��d�ُ1�Z�9���!�--�b���?Dt����N�����a\��w��[ ׆<�R�|�I o�d2'�� �$���>��{f2��A�|u�n����Q�{S�u.�v��wm�f ��q�9s�_���\.w���y&�9��D���    IDAT��:�a`f)�C�H$d������m��Ct���_~��Dt�QG�0�quP(�L&�+ \��5�̛7��u�m�Y��΁�I3Z���d=fT赝"��F���W�ZŎ;�͛��Gy$�D���.2�& 	�Y�wuu=�:D���߭:���3��O
��T��8>�1�r�|��y\-<��;���d�c�7�=7n,5���K�����pT�e��>�~xD{������r����3Ϝ�:G#�ȪT*7B�34�h��3��Q̌���|H�(�6M󺉽D����� ���
��J�Px��c�8�u݆��z{{��j�& �9^ӈH��vY39)�cF���N��ju�۶OWb:�m_�5�sioWC
t�*f^966&K���#�� pO��ѫ׬Y���fac������F�~�R�:�Um�4c�T
��_٧YM���S���Z�5BDteOO��;�g��w 8Gu!�DD�ޮ�a��F���?��fOQ��C��͝*��;�Y���U瘌i�H$��hW=q�+)�E���ns|߿���w?�A^,�ɼ��/S�C������Hf�E@����f��,�Es�̹�ΰ�%�w�=fTe2������ѵ�]LM
t�D*�ҭ���R�|�����r���s��V sUg"l�jU
tÐ]e>3_����(���� nU0�+V�\�*�FJ&���q+ -w_K��Z�����wL(AD���R���j��J-�R���`�9�P�Z���G�,��q�L�\�!���T����b�Y�T��2�f Tg��eYZm�<iq���B��ѧm�^�: x�w���d-�f����V�!�Hf�EЈ�s�L��9�,����Sa�KD�""�&A�m�WX�:�d��mϧIi�M���bF�'U�*IDt��8�� �|�G ��W�E��ʊ�t��a�uG������} 7):�z�j9Af�m���ix=)��]������I���W�pǲe�� �����^��>��8Y�3�}�h� W�n7!��͝����E��� |Au�z�����bj�8ft|R�c�;��r�|[oo�O���Sccc�#�;Ug"��\�0��3��uR&�9Ou��Z�n��P��O���ӿW:$�L�f� -7?��8c1R�-h���Q�j�j]��oݺu�뺧Bӣ<����I�.چ��#�ɜ�:GT��
�����{��q�c����a�`��,�tuui�-+��]E$�K�Vw0��m���5�\u]����/ �FZt�?�W�jU>WD;Dt���>3��_�h�ط������� }��ԓL&a�ZN�&I�3:��ט��k[�g�y����<�b 'Avx���A���0��������e�l�֯_�'"ʅ=.3����_�Y�v#"�T*W 8Zu�z��k���\��$z�����H$t|�G ��m�ժ���u���<���,Bh��yϪW��.Br�m۟W"�Tl�&��(W�L�� ���ٗ�.�H�3�?��}�h� !��%K�����B���4�� ֩�"D@6�g��.Btn6�}��Q��7@������f����Uu��Hk{�]h�0$�I�1^���q�ng�n޼�i˲^໪��*"ڬ:C�I��1��d��媃DI.�{��~�`��:�(-��K6�}-3Ku���z�,Z#�В�O�� �9~�fpp��y� ���#�L1�f�⌈��C�if����o�� ���ݬT*k����qj��va7���Ku�R�ǌ�-�������L���������� {U�b&�hHu�8�}_f�E�)�W�r�i��y3�QCǢͽ��w�a? ���,SI�R:Q, �՘���?"�vGJf>=��|]u��x�w����pUg�Y2���i�e�D,�5��|Ju��x��w1��
�>�#����� ̟?N�Z��e��LŲ,$	�1Z���0I�3Q����@D��l6�1�9&S(!�� �~��0c��q�����"����m��:G��hs�i��P1n����t�ff^�:�tt��jV�&�$��^*���f�/۶}������O�����Uu!U�V7��s*�f�  ���[�d�+T��]�v� �Cwd�;�֭[� �W��L'�NwLk{�&���]��4?ߑ��L&s�� ��<�4"� ���+g����E�D��1M���˗�SDwc�|�������~��Y�L�"f>Su��tJk{�蓓]D�eY�,Ku�z��a�d��᪃L���|>�i"z'd�8���� qW�T�@���T*]��F�:bf%m��Y�l6�q"�����|�jFt�UM>�b&�O����tn�ُ�~��dQ��|>�=f>Z6�{Ju��۲e����Ŷ�SBw�<��}P�`�k׮��,��f��d�U�hD:�6�uI;i[�1͟�7ㇶm۪���y�c̼�}��1	)�cf@Iu! ��8��U������=C/ٴi�k�(�q���W!�P"�й�TL�H!�e�&�ɤ�S�!��-[�l�� �
�g<��+ ��:��bf)�� m�B�{zzUDg��_�h�H��g2���@��:;,�C
t9�TJ�Vw �+��?����Ou�z�����@�=Z0�i� )Ѕ>����lW߆r �P0�i}}}��m�>�0� ��:K#���:��]LM�*G�z4ou�WU*�d2�n�A����a������"��]�]���r�|�lW3ߨ`���͛�&�$�ͮ �{h;���d2	�����	�a3��CZ��h�4o���׺}jhh�~ � ֫�"�MZܵ!��
3�l��gU��]5G�F��=��.g�8Pu�F�!��1%��*�
J������\.���i߻�Zd��T��O޲e����A=��,�:������bfiq� �q�BG��m�t�!t����N��'���Gb�A&�q��� ��҈N<Rm2�2q4�P{��ɖJ%���6ThדL&��ݍY�fMZ�w҅P��Qe:�r�BD�0�㪖�Dt�m�|� O��T*���y��BL���ʞ��Ǉ��T����u �y�43�
�;!�۔ŋ�7M�G zTgiT&���I�A�pň�"��n߾�������s (�Jرc���1666�x-��n������m�[��7���u���T r�.´{�֭{T�  �>]��}��E�-PD7�r�z ���%"���m�>в�{����4*"�8�I�A�]!"J��� �1Y�Z�3�<��{_ة؉B��2�϶��u/� ������ 6��"b��:�'3�Bs��e}?�;���c�=��}
��˕+W.Q0�z{{�#�8Lu�fġ�]LM
tE&��+�خ1�۷o�t&�Ӥ��t�׶�U�h��y{5��Vď��k��d]h����Lu�0�u
�5��no�����*�ʏ1�	ndD�(a�	P�ma��Z�މ3���J���g�ٯ�ш�[�����9/]��� "�A�c��8�s��:I$�@�)Z��/_�|^�R��ժ�4#N��5�^�̔�
L̞>��*��6R�ԋ!�H�����!3��m����(�u/'� ��":���}_f�ET|1�;Uu]<���� ܥ`�#׬Ys��q_b����J�ҏ��y-�ck{D�_C'�G u���E�Tju}�q�ϩ�Ѩ|>�K���=�:��<rĚ>d]D����e��H͔���6wT*�w�w_Q.λ��b��ީ�����O�
Di�_�� ���#�J�X\<7����O�!�n!�N�������#3蚐5�"b���6۶m�AtP,��\��ѻ�s_}}}sK����ܲ��t��pD㧁�4L��Z��:����R �C��� �l�/�R� �H(9\�e!�H�\�̒�Oضm
��s���8�q�u .C�?�BL�4M)�5!���Zb��-z�������smܸ�������<��V�\ٿaÆ\���f��pT�c�*�K"�(�ǟ���:DP�U4n�g�GI:�F�Z�̿��>�8�,"�gf�Dh�u��m{#��WuyR�k���D�Y�/��+��UD�6*�G��:�_���D�@�������{ �	sܠ�R��,��J�{G}��mO8"��; ��϶m�2"��u	��e�� ~�:��6��e�&�y��B���3����C��~��_ ����ޱv�Z3��-[�����#��y"��Eg�h^T
��� �$.3#�V��y�m��QT�[�y޳��	�y谇i"4�\�Uq4��3oW�A��"�sG�zh�&:nP0��?��O�c��K�..��?pX���"7��q�I��]n��V�T*�]1��8�w���#�t���u���T ;U���j变��"������:�JD�d7��6��Z�dIO�Z��C�=V�D��!��T.R�(NO��]]]�c4���nٲ冾��H=^���wT��W���,"R�� ��T*I�.�.	��l6�\uU֭[������N;���v��d^n��� "��M&��k����1� �@2�Tc&�V,���뛫:H3�z�!��^�BȖ�1Ϩ �l۶m�D�!�8���X�|�<�AR��>�\.�u;޸��畆a�@d�ԋ�=�QT
tY��8��$�I�fh����b��۶T��\q]�<"z+��*����@׏l':�+K��uD��V�q<(�}��A���8G���+ K�~�0%��Xއ��I�FE�@�� ��b��fG�U&�qTiV>�����É��Y��|ߗ]?��.:�_۶�M�!Tx��7x(�q���Gq�~A��mۯp/��zOU��"*���ڐ���J�.3����`�fd�t"z�a��m�`�Y�U(\�u_�s��mbr�I�~�@��}�l�c�C(�b���eYo��y�`N遼��Q)�'�qҰQ)�;�^Ղ��n�q�"�� =D��L&s�� ͚hy?���70��y�^��]K�4Etf���8m�a\7��� @E5���:��~ �M �9�2���Q�˲�G\'�C�(ֈNp���U ��7g�ge {������ g�y]�,Y��a���;�Ej˘###Q~P����S�½��̄m����/�Q�Eh���ޢ:��3�q�� n���L����,
�V$L�W������~�R�>�装���q�s\p&��i$�9U7p{��	�~|�뺑_���h���|��T�� �|�\�[����ۢ��X,��2S�ø�q�wG���<�#��m���� :�<�Md]K��.:Q�0�;l�>��?��� �]��Db-��5�""2m�����K/�{Ѹ��,k+�1V�>��Cn�o�D"�3(� ��8�'U�	f���{>3��i�y�ZR�뇙�@��@"�gѢET	K*���^C7Յ��חr�zĤ8�)��mw���I�� 3��rX�fϞ�p��J���U@ .�m�""��?�󼟕����Xu���ؘ�1C
t�ɖ%�;3�L�� a����wѝa�����W�~y#�q���⏙��v��Q\�t�A�\$o�;�� c�y��`͹\�È���"��ٶ}��8�l���y�_c|�w9�!~x˖-�!�~�@��H�4���3�b7w ��L��K��x �k�G_q,�e}rq�P�3�p
���g֬Y2{>�0:���m ~��dRd&j-� ��'�qD��3��7�)�E�c��m����a`�{��HKf~�T�8Κj�� �CB���b��R��:Fhd�prR�+�̛ ��X;��ܹ��������}�ݻ��>^m�o�y�� 3��C�bq%��Ug���v=IW���O:��A�!�-�˕���
�~�ʕ+�'��qN�3 ���ccc�*��KI��3opd*��$�����4,X��sU����,�k^���Lf�� 3�m۶ݮ��4(x�/B'��d�83g�ٷ��nG���0����g�ُ�@,�h������T��D���f��a�_�J%�J%T�U����k��a��,�R�i�8����\��k���ު:H+z{{U*���&�YD{0���u��q�ضm��:�!��x�uV�]��V�Z�	�Ґ�~jٲe�o��:q��� :�k!�T
�dRu��ٽ{wo�q���f��$fϞ�y��a���o����s��Eww���9���j�s ��f۶?�:H+�=�;��> �׋)I+��*��̠���pے%KzTiw����lڴ���ϟc����a����{��=��zAT�U������o�m۾>�;� 3��|���a�б3qED�Tg/5<<<�3�
��o�i�?�����|�YI�{�\~oWW���Y��Q&���#�����#�w ��e���Ҋ���'<�;��?@~Su�Aה�C1u��������Ui�6<`c�c�J%�ر����qT+�JR�ǈ������|�.�˹L&s�� �`��y_��M_�:�h���""�ވ�zM�\��{�f�膰�������~|�WD����=��T��dC�Fنa�2�͞�:H�����<�h �Af�#�0��3���@�ED�ض�5�9ځ����#fƞ={�k׮v;�R	Ţl���@���lW�V122"���f�[�9�"�����u/p$d6=��y��brD$G������8���~x�����̌;v`dd�]C�Z�\t�?�O
���Q[s.&e� ������7Wu�V���[��p6 yT=2K�)fު:��R6��;�!���v�i�Zų�>۱;����#>O�VR��P�_q��DtJ�X|8���:K���w]�r�4!��T���}_f�5EDR�3_��fߠ:H���� *A�����}�YT�� �V��vw�O�O
t�03*�
J�R��U*��~�;����i/7�l6��A��y�����Z��O�W�GL/�L�tM��/G�	1.��7e2��م������?��FFF�c���
Y�\�t�.&g�  "�/�J���>����'�L����g���Y��T�U�ݻWu�(��̷:���}��}ՁZU(�����E�X�<��|�i�R�����z!^`�a?t��uT�	�a�3�	�����عs���+T.������REDf�#�3�ill콭��x��Ν;1<<��וJE����sm۾}����T�	����.�u��}��U��s]7^V"-�B��| �,Z�h�� A0M�f 3�~-��x��8�@�R�\i���M
t��� �p`��[۠c���A���jJ"'�������番��P(��u�7��"��U����ޮ1���@⥖'��3�L�� �z��w�g&���o.���Q�TP,#S�Ʊ۷QR�+BD�v��s��Ig��r�6B����+|��9�󏪳�P(ܻp��# |�� "�>hLZ܅��(�0n���O���vs��|�N����J%2����O}R�+@D� .
c�N~�)�y[u��q��z{{Ӫ�%�˕]׽�R�LD���>Y���n wPBL��[�l�_"�����9s�D�G�����۷���+��rq��P���H�13wd��|���J���q^�:H��~��m�|�_��r���r��r�\�E���˶�KT�h�}��Wd�ۧ�{�#�Z�/I�C&��M
��Q7�S���m�Qo))�ˑi����`��Z�A�6<<��u���` �Bf�CEDR��O֡1�:��I�!ZaF�6�ZK��;���?�%V�H�.)��w�P7�}�;lFyS��ښ�?d��9D�=�q.[�bE(�a�<ϛ���� �@��B��R�kN֡ѐ��o��ٳ�I�U�Uii�8��t�������!�E/j��y�s�!��<��1՟���/Tx���#&	���[V��L�<d��mR�]�/_>�T*��OX�8N'�O�u�UB��8�-��K���X��-���D�7 ����cccعs�Q�4Mtw�u�@����]�= �7�E�bW7�8Eu�(�w��(Π��e��}��5��?j��<ϻFu�vx��'w�����[���CD�p��\�Ff��GD[�]��� ��?q�    IDAT�f�o���R�Y�|=� ���#���Z�b�޽���d7Qiq�E/��͖�Z�CDW;�s������.c��]�yޡ ���#u�0�@ל����.D㺘�N۶W�Y6l��R��{�9)�;T�Z���h��8�J�ޙ�)��T*Iq��w����e2�cTi'f�]׽�u���/��2�:�����d�M�GD?X�ti�� ��d2g<��sd���&Ez4D�@�� E���T*�n���c���9������1����|>�O�tz	��<�:STQ��a�Hvq�yK�����ŋϷm�v"���������C���R��z��pA�Qj�c��m�?�m�V&�\׽�� �7�@Eu�(�}��bj��K�.Ds�8�I��WOOω�e=JD��S�T�U���(�	"��J���2� �/ik����w�m��:HX������\�=ղ,�7fO��2��?iq�a% �W*����{���(����M;�s���?��T[��+mw����RQ)�e=@:_����#��m۾�q��:�b:����7f/3��� ��IS�0�A�\"��t!���M�i���O?�����9�R�� ����-!"$�I�1��rM���*E���⼳�;���L&s��,*�w]�l�����Q ��Τ�J�"�����bRDt/3����k7o�<�:�T��r�\ 8Tu��$	̚5�T
�TJu-�*�u�0T-*�̠w���1)�;-4��q�^�`�l�yT(
�x��5�u7�P �c�ͪs���,iq�3W<�:��Y�̯���'z����0�Y�d�+l��5� ĢJ5]]]H�����&�I)�먝�f�,z}Q)���}�C�o���J������H&��s�8�ATz�u����r�0^�����"ϟ??�����6w!�=����<�>�a�CD��8g����Zu��$	twwò���Y2��v�:|��H���^�����̠�Q�ƷVB�s�����x}���6����WR��-�S�q�jYֿ�v'@f���~�q>��'љ ވ�|.��������hx�+U�B�<�/x�w�DW����m�; �V�%,D�t:=ia���,���T�H���n{-3��Q�8Dԍ�[r*��I"Z��wx&",^���Yt�4���f�IIqkO2���0�l6���O'�3�y��<m����U��s� �V�C���eY�D�2�m���U �T�	K"�@*�j�������h{���S�]��M�#Q�w"z�aa��J�0���u(��CQ`|��7��⧶m��ma���9���3 ��"�y�`�u�e�C��9�� >�:�!���b���(�~r����f9�aH�R�Κ�#������k�����0��})���Ν�p�*��a(��ϟ����g�ٷ�������]�=��<����; v(�$YD4�:�!p�a�]�=?*����� x1*ΧZkިT*�D"`����t�gR���= ���vwwk�ce�XD�,�N�,a�۲�썙L� �at��U�u�y��{�w�>���T��E��� �נ��� \�H$���{����vՁe���m��ňIK{m���;����u�q��R�+ �<�S�m^��H$����O6~;��K�������JM���h��骳芙�CCC���{v:�^���) ��Ku���`f)�E�*��4�W��{ΦM����(�q�ǹ��r �U�	�eY�5kV��]]]R��Q�I�}9T+,R�+��� 8
������t��ϟ�ɢ�c�8�ϲ,��i$	̚5K���@D��F�q�\�dI��<:+
w��{�eY���o@t
ߨ�=���@���"z��gn޼yPu�fLY�(�s��!�N����m��R����>FGG-�eV�>)��(�O�OD�-���,p :蠺�:�}AHq^�i����z��k�f�,A��L�|<��~����4�����y�;-˚��̺�E�^�Dc����@��'�� ���|>�SuZ��d�f�Wa|r�`�qBc�f[f�'#Ez}2���]��W*�~>66�j��j��c6��a�4M�R)$��i_cf�
g����Y��������2�~�����¯U��E��J&�'1�i ���'~�uݳT��qg����>}�Z�~�P(�Au�fe2�3��" �:���a��{�6|/7D����wwp����]i���d2�P�����T*�ch�4�iל�f���rP�PD�a�a��8ε���P(<�:PT�`|S������K�ұ�a���=0��FD#*�M�\u!�� ~�����c�����&p� �j�Y�T�Oj�_��������`f����|�L�'-�1�!�y}���F�P��d�צ  g���q�")D���`�P(���9�����_�O�"�*Ẁl'"�����*�uO�</r������9�s��&p�)Ή�T*��Vstww��ޫ� ���V�>)�c�����5S��K֦?�  �ٶ�3�q�Bu���g7��\��3c��Xb)�#D�B� nc敮�\(Q�YDD�㼻T*����M�L�Dww�Vݤ��w��l3-�e�>����v^R��gF˻�&�Iy�;�u 68��u�q:jݑ
CCC���{����i.�"z �7��"��E�̠���1�w]�T��Uh&zzz^i���0�ɧ�eHa�a�|2A���T�"}&Kd�>�i��⼾�xF:>aV�� r�"��S� l޼y�u�K���� f�' w(<�̠G���M�Dt����N̘oPh&zzz�w������ب�Ю�=u�L:��`�&,˂i����jkқ-�e�>�$N�l�f\Y��+�J��,�Ÿ���?��m���l6{N>����@��u��� \�8N����Ll2w�%-��̠G�aO�͔�H	�`~>���3SDdٶ� >`��<ak��!���v�X�D"1e�e��J�2����L�tyC
t�fF�X�⼎ �ڧR{��QQv83��q������z�!Ձ:�뺣 ����C}�?�I Vb|#�f�z�����������y�ô¶��۶�5 �������Q+�j3�{���~��0$�Ɇ��3M�i"�L�Z��T*ͨ+���{Ծ���]�X�8���ɵk�|22��'��y��8_.��M5&644�8�����ۻ�R���d �0�� �ժ̠G���ò^P(���х�|�)�aZ�8N}��NV�E�d2�ok�v�����o��5�mh\*�P*��z��l��?�P)ڋ)ČqA�.@)�'W{����M�Y �O$��W֧�����f�u��� ����?���^CDR�GH�R�t��n 2�R�uωrq��ۻ�m���̱+�;�4�vwG�T��3��qmc�f��R#�������k�9���s��i��3ݱ1t��Z��l�>��� |��Tg�����e����� ���c
�¯��#"ö�"���%�h�6"�$�H|��'�ܩ:L+���[�l�{�t�9!�HtDa�b���u�����`Y�7G���IDH��u3X�ow]��N��]Q*Х8����R��7�b�rYu����?�#x�n���s��� ����E�B���Џ�8. [u����+Dt�ľ�ED��dN#�/X�:�
����~>�j����Q�Ez�7�k�aD���@�O
tMD�@��ڧ7k�,�~���C#>}�R�|B6��q��<`���#�g�K��w�9�7�m��a���+UgQ%�k͛��>��ı�Zِx��})��ӫ��i�CD���nk��4M̞=��<c�`��M�|�q�K-Z��C!f��:��(>��|�?�u�~��zq�����l6{#��⼓֚7�����5�a}�S�Ԍ���&�9�U"�\`���8�\m͹.m����i-75Q��������g�ϟ���Bt>)�E� \S�VW��{r�Px@u�V-]���q��}��3��:�*�D"�C�H�,+ԯw+m�/.ҥ��>)�c�ы���D6�O�5�ӱ,�f͒������/�N:�s��8]�	�))�E+�p!-s]�̧�z��Tj�m۶�8�T���pbz_]��H�ӱ�0M�������µs�}��8��LG�A��F.
��;籶�'�0���C��Q�VQ�V#�  J�yMmWM�4166&O0��@  ���8͛7�7n��b+!:��:���M .�}�ۅB�#�W\�x�|˲>FD� �"�Lm�v)��Y����n��Ώz�z�������Q��i�����1��S~��֜�Z0'��i�oL�|~F��Q*�f�	E��u�EX���E��z��;w����8��<��" 2�.�� _�<�Vf����:2��A�a�kY�?c|�Tl��T*���v������� "R�`���pN��V1�ښ�V.�D"�Y�f!�J55�LDH�R�3g��m�Q/�kjG�Ľ-��> �ڶ�G�q�"��Åh��b:cDt���Ǹ�{�����|���s�9�0�?�8b^��֚w�}P�X���{+U�mA���2�>�����T�N�aY�ŢVq-W'I$��e6�%��̶�Od��/��{-3�IĎ��O�Zx��J忟~��m��%��DD�����:�j�%r�v�.���b�ؖ�����%�k"�s�';���✈ڲ&[����J��Z���\.�����Z:�������h�Xq�9 ���!�@D��I�P���\.Z�hA"��g �� d�y+��r[�t"��ٳ��hxdZǝ�.��b������[)�j�mߵ<*��8瀬Mo@�����G���eY�����)@
����F _���S&H�L&k����� ȉ�Y� �s&}�=��A&p�O��������9o�k�F!�i"�J��Mh:�T*�yMmm�̦O)��r��)�q�eY�Ń��;T���
 V�!�X�r ׸���ݯB�t���j���0�B�weߗ̚'�H�������~��	�N^�%z�1sn��d��&�H$P.�C�`H�R���tT[�>::*�u�B ��T*�m��J����᭪s	�&r�Z�0�"�
�����4۶_ED� � �:3��dּ=��$�(�ɦR�����=�^0��K�Q��lX��6^\��"Bww���>����_�D�q��3���U�d'��Wp3�]�h��V�����8ΝD��wA���Y��Y�fIq�&�D"���J�j�c�\m�8��/���j`��a~��������C4�d6�a) g��.�q��y�uVJ��H�ޙ|"�3_�N�oإ:P�������o��1_�:�nj���i9�*�ɦR������!�n��]�q%zL�^��	�eY�}�ՓL&C�����l��Mo��$ 'e��{'v:���������! ���C�PpUj�����cccg1�9Dd�Σ�0��/d�^.����]|�o����3)�EKT�����)������X,���0�	Dt�m���\:66���[��Q�K���h� ���̷��۱����ޥ�J� �0Wqm���R)0s m㣣����~��A`f��P�W�8)�EKT<mmǇOM"��M��x�wѐ> ��J���8��Z������ͪC	ф��e�d����LDw�����L����s,3��O����e�&��t[���j����̌�����<���LƄ��EU�l�5��K�9�������x����H��+�����/��3��{���^�a�h��8��V�C�52���^�0������o�z{{��ry-}�a��茈�L&e����@f҃�K�Z�btt4
����{��A�'�B`�U_��gNf�g� p�a'9���o���]'��Bs�CT����7 d�<��1s,��N�_�� ����W�Gw2k��t:fF�Ri�}j��J�TjF���y�c�:R�k��#����JfЃdYV�gHv��Sy˲d6}f� pY*����8�ѷ���Fա��DR��R�[ 0�z˲~�y��Aա�DD�m��� �92�!rl�����0::�r���V�T`�&��$LӜvYj�ZE�RA�\�¬��ZCME
tM��'��/��䘦iJq0�0��ݍR�$��33����������:� ��g�|���`;����.`�%Lł ,RB�D�&4�6U��Ҩ�J���6Q�V�ꗪ$U�B)A�P�*bPp>ʚ$�ر��s��m`����3s��?f�@�ػ;���;�O�����#dݹ�}�=���� �
�� f�"Z���W�qyQUwx��7��=766֓����V�uW�T�,��]�I
N͓��%xs�:��Q���{H�*����&�������:C����D��z=��f���K�;u��伻��r��e�
�W �������W���Aס�籠w�������3k�O�$��u0��2-�,��r޷.�����ׇ�'Ov|%bEi]�ȂN��y��I,1�ˬ�qk�ڎ\\�(Swe2�Z�
sss<?sy6���~qa��l6�����n�Dg "դNZk xi~*�WU_�d2�\.��W���i��pj�|����NcA��ظq�G�qcI����N,�^X��∸^���O����Q1s��d��{���7T�� ~�:��(�����4���TT��b��x�W�V�㽲y�R����fff~MD�V�[�{�%��r��6D���]���P�
:�Y���g�~�4q
�BG�tx/�V��{4K�r���]�WD�����T*�|�G�Q*����~�9:m	���4�ry����7��:ORc:~6�É'8�x"��j�z���ħ��2��t,q���޶�D�-���G�����izW\���l6�������B���\6Kݠ���(�4^L# G�ީ>��Z;n����Ac��C�-�È0444h����b>�:O����,��)�0I�=�i���i��ǈ�� ���K��{w���.��ԭl�<�z��lv�q ����Z�U�';u���G��!i�L�����[U'Uu���ƍ���Q^���X,�g2���� >��ma��WN��Z���Y��w�����a�9:��x9�:�rXkq��Ɏ~Xt��r_�Fp���|FD>S*�j��?j�yx||�Y��(�D$P�8�WО|0!"GUur���Ƙp��յ={����$"�͛7�h���1�㪺�u�4�Լ�,��r��Ni|��)��w�ꃮstB'��h6����[ֹ�|�������"�_"� ߗ���}�1 ��9`JD�T�m��Z{�sDU'֯_��;>D$S,?$"w ���\gJ�k���a�o�Xk�Z�v�u�NbA���/�S�9:��\.��5�n6�h4�~B��y�Z-��u~�� �H/�C����?��E��:�%{RU��^n>`b~����y� ��1�C��pl��b�x�|)��י�haj�������oS	���!:�=FDĔJ�# 6���I"�L&��`����������Z�V��V�ձ������y�*���8M_y{<E�C�\��x+��wϿK�֢��B�V�W=ϛ�WEd�e;}D$S.�����ړ��Li%"����ԜN�$�MU���w\��4���}�Q�?�h���=:�-�� <b�yd|||��0D[�l�����оO�R6P�#N��tX�U�t�����i,�1���� ���I��y�Xk177ױ��$c��-�v�Ϫj�:�����U���""���Zיz���P(��3�^��tU��0]��4��9��.���q�#�V�Z�r�B���ƫ"���|>�̓θDD�7<<<�j�n�Q ; �&�-���bDQ����^�G:�E�Ctz̈��J� @�u�������Y)����뜦�GCU��oy����C��DDK#"^�T��	�� .u�'qjNKգ%�_� ������C�����9�����N�ck?�� �����yB�6����ͪz��|�9�3�2N�i�z��[k���j�w��X�c��������iz�D�G��mc̓�j�y��S��ÅF�����e���9Ʃ9�Wt�  	IDATuR������+�0���ނ=�|��1�+\爻��>~��0N����t��L&����Ó������0����,"����Eo�Ԝ�!�"�<��El��\����*�J_��s�#�X�	�N�	�sU�	��V������Qׁ�ҠX,^l����z����u&z'c��<�a�kR>IW�R�V��-,�1588���� �]g�#�s�E��'��`'����L��8�D{""��_� �[ko`!�?N�i��Z-�������a��:G7��ǘ��� ��s��9���bvvQģ�L��}�E�j��~ס�\�\.�Z��� l��m*:["�|>�l6�:
��f��z��:F���ӮCtz��J����s�%.
�?��8MO��D��Tu���Yc̮ R�v� ������Ƙ�D�:U�pU]"y��B���99����� �u��X�c�����]�9���Z�z��iz:�x����Zk����ܯ��u0������\� ר�"2�6u�](RT�?����m,�1����h/���5��|����i:��� �W�Qc̨��A��PD����> ��ȕ�z�+� `�KN��l,����Y�{z���h4�l6������0�N��joł� �R�oE�]�p�圖�Z���YX�k��𼈼 ��(�^���qll�OlhElٲem�Ѹ�Z{�|!��%���i�yr��Y��n݋/��v��[.������-�U]�Ƙ���ǟud%��'�ƍ�
�} ����4�s�N�i^@��w�ꋙLfo�Z��O�;�mۖ=v���(�.��D�RU��� ��|DDI�����o�αRX��\.RU��:�J��r���cP���t:�� ���>�`��v���`ett4�k�s6mڴ:��n�d2[U�"Q�_p!8'"��f�y����Q�AV
z����'Tu��+�场��hp�Ng�	���^ �E䀪V�������ӥ϶m۲�����:_ķ�`+zp%�K"�{�j�_]�XI,�	2<<<�j��p��,ݔ�fQ(\ǠE��:�M��j 8���cLEU+�Z���<8�8����LfHU�DdHD�Uu��%��p""�T��Z�����0�=a����T�1 ����\���C��p���U �Ƙ	UW�	 ���Z���!�dxx�`��`sE�Ed��=�P�����(�&������}z���W�?p���X��%N�ɑ9 � pTD�Yk�c����D�1�H��|����x�M�E��`�=�Z���`���;��&ٌv	���DD�	�A<�:�,�	422���������)�l�|�煒s��SL����¯U=n�9��3 fE�uUm��y#��"r"��4T������9��j��j��K	�iӦ�}}}�(�L&�Y7��� @E�UU�1kU5#"kUu�1f����NU׉�U]+"k �A�l�_��!""J�?��ˮC��P���p��,�%"K�n�eޘŝt�͇|oQavv����=�H��'DD��P�V�T��w�V,�	����������u�n�^yȱ�_�h4�䝈��he�,
������1;,�	W.��V��X�:���y��:�:�k��Q�T���D�v�7""""""J��l�f��6N�S��� |��3}-Q�6��[{�8���=%� xFD����BDDDDDt�-
7���z�T��=��mp�u"""""��x�P(|dll�5�A�K�S�.X�h4����k��0���G����)�J�p/���<DDDDD��Bk��Zm�� qƂ�r�ry��>�|�Y������'=��w�a��� qǂ�Ve��{ �	8M'""""��1��\���Wϳ�C���E�L�Uu��,DDDDD�Z���N���ǈ���;|ID��!""""�ty�Z{O�V��� IĂޣD���_G��_�:%��<i���0�:K�������~�����]�!""""��h��c �:ß��,�t��͛/�d2�p'��;��� �o6�NMMu&MX������ ��Rי�����ș9 ?�'U�� �\J+t:����(�nT�|�V }�cQw�`��|/���Ƙ]A̺�X�i�DD��lv��nU�� �Sյ"��* k�$""""�w�"2���8��o x�S���\DA�됽��������(�� DDDDDDDĂNDDDDDD�n|��1l�    IEND�B`�PK
     uK\��C�I  I  /   images/d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.png�PNG

   IHDR   d   S   i��A   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  �IDATx���U�u��0<��y#�W|E�b�M�5V��6�������Sc�hMl�1I�G���51jbk5IU���F06A"UE�	�0�83�c�a�������s�=�{��~]߷�{�9���^{=����7`��ɦ��ǿT+8Qp���
{w򅱬��1���z�B��O?$8=����8��}����8<�}�1A��'�s�ۥ��r����C���O��ÇM�~��._�
��54���u~www�D�
t����wK 8�Np�`�`���"�>����0�mۛ�~�3v�	�_���r�u��R��3\�g&�@]]������_9��Ѓf!=j|I�E�u��	6K��%��� 8Dp��$�Y��
��#86���F�7hР�8y'΁�	絋��'�U������uMxQ�Cͤ���ꊈ4��^&���1v���C[��@�[p��s�fm �s��y���f������Q;!�rK`\ ���͡C���&�ǂ�'k�ȭi���y���}������g"
� b����|Bp�I�?f�l-8��C�S���b��竂���/c�}�������L�7��O�3����\�`~����N�jC��+��rD��$��f�w�Q�gq��H�~k7v�R���XL�so0V� �]�q��e�o��]"ߗ
�zX	��~0�&}� �q��'�5�S�52+AJ
�`���r`~'E	hY�d��'�%����K��p!�"���D�(��?%�Y�q>#���%�	����-HDc��S�uttDc�Qv���� ���@2�<��Cs0$
���*��4n�\�P����N�/����
n�5c�!S� !�pH}���6?%���|�Up�_X��0�>1�eT�;�H��~�=dȐh��L@�3�>�`���zfWða�v�{�ƍ�˭Ok�1��36g� T;�T�4�*�E�{�7+��J���I?�I�����	��P�R��*���ݣG��b^-?뛛�omii�$�8/�3�˂�͏$.��#��0�,�	�A�@����1��O��q 1mY�bOVE<��t�҆�����,!�b�U���ۯ*c��D�@�Ϗ)S��-[��k��Mu���Qx��#��F��!��\Ey�T%��BL��|�c`�|�-�lr��?'��`S�=q�����8S���/�D�rW
�,�wq�)�,P�X��3���X/�{3�A��1.4�X}B�,Vtm۶M�Yp��%t�.�r"R-(��_�Q~�+x\X^��<P��`��:{`mt�n�{���}F� -��3�}�TF�Ǔn̛7���է�P7jԨ�{������v�?q0|�y�*�!��|�`��=\�x�9�����C)f0��0I��X ?�/,X������4�]xekk��q^����	FO�
A�4�� �#� �ϭ��"�������3g�M�6�nz�f��Y�S����2nܸ!��A�뽂��b�e�p���-�8DT���4�'YEWE�E�#0��&oV����� ��9�FP��E�������f":��y��k@Q��B,B|��	��o֊�F9��]$U�*���lM����O�� ��ޒRn{���Ks>|�� %Q���o�䎎�C2����P����a�cC�K�^�UAQE,�G�����8P-��a��w��%�MNb<.3|�����4����|�'�\&�xF��V�>*�*�����ͥ�^�+
��x������5/��r���2p�0�	�qG�2{�V*��	&���/��M4�ս�bM	w|9�
��]�W��`�/�ҠAtQ�a�k{<�%�@TUCo��"��]�n�{�tV�E,(O�M����E�"!J�z�!,(�����2T���@���I�,�K
����MG�	��̾��ZU�����<y���s�obz�9��2]@��Sf��?��}�m߾�O�/���Z"��j���Cc�"�M��IVWn�0�@l0VnF�=��E���Y�_"��&a�4'\&��W���{�d o�s�|��Y��_��kiiQ�L?N��FV �&V3�׋IAH�J����������H/"�;Y�F13��<���2�mӦMC���"�f�PF����i��7���755�?Q��h'�z�޿���5�d��l�^}����I�&�k�@8B^�7�����X�a!s��':�h���뎝;w*q�ٻf�?� z�5� [��o7v�J�J���_�=����4��x�c�E�Z*�#�r����666�'��Ῐ�7����`�}2�|3�:�g��S� �6���g)a12+a�?2v-39O蜥^�~UpP����o׆�5 �I�f���} �����}���YwY@	��TWI}ɵ32V5��D�"��s�<?!$@�Θ`�L:�b�]�
!��P��X�gJH�~)&�_�㵒L�
�hӀ4 ,�>�4�n^������[u�@�_�%��,j��9�L�:��͛7�Q6����e��@���u���* i�������U��"!� �K�ڵ�T 
��M�6��-�2��.�p	6:��mG�9GO0vB�O*�� *C��]xX�p�8l���w�c�-�e���r�D��1�|f��*��f�	
W]ƿ���������zIN�GB�y��+���lv�X��&�yR������$3�*��s?ق�Gj���M��a,�l;׸��N��!T6�X+���ٕ�^�QD
��B.�����^��!$����;�i!��g���A������L�X�%+����E�(�=�P�̒�r�X�&�B�u�$�����Դ_���ls샆�p�Dd|b�D1��������OV���9��e���ث�Ʀp��
ΪnY`�M`b�56-	O���'��� A����J�"	�Q-B��!q)DY#ˍe���fo�����I��!��W8C��VWlJT�t��y������-��
��Xfv'$B�c������u�<"qr�=���[$�r�b2�rc��z���"�M���2y�VT�9��6lX���w�G��39 JL3f�Y�zu���YZ]Ie�z��s��5���2�{SA;����BC�i����on�ԩSu	7�ayCB���Ŧ �HWID�rVqf}�A�ys�M^����S���	10]��1�F���PF��ɚ	Y���M-G�V$�j��B�e�Tͼ�{V%�� B�g8d;��4����J"�qH8(Z�цH�5G�� W������<�C��è�<;$�#H��ˍ=���IKͱ�]�:��fAG�śBd������@D���At��'v�9��~���o���Y��_0v� �.�"��W�c��Gc��Z�`�w��!��,��+�� ';˅,B8�M1�).)����f_ɇ����g�!i���K��'	 �r�o�W���dEh�D� Ib�ƾ�c	�{*�8��������z\�����i7��3?cB�`��=����I@�P̕����$e�j�%��"Z�LG�,.S���+zJ�b�F�Sɣ�Fp@1�m.F��9J�am1��r��$9`a@�����⸩���z^��֮]۫`@�\���lm^@��s���M�ِE�[ӀX�g�+T� g��������c�ql�z�?��=�q�6`�)�ω�`��z�^�\�5�ё��Ϧ�%����EB62�l�o�z�8����n�EI������VnWR/���*�������ȭwĈ��N��UQ�ó����*�JJ��Y͌�L����E9bx��:2��,"�p�}��� ±y�L��o��� �X��E��PS9�TM��ⴂE	5ֻٰ�.�R�ܪ�r�#����p.����~z����:t�۷o%��XeX1i&9��F�'nӏ;��	�ۄ�?[I��ِlV:.�`Q���XXQ��q�)�DIN<�%-71<?dȐ�tvv;R����V��B!���0駶8�a��O����y\�	v
<��p%�C{4_�L�Ę;wn�\FQ#F�@��r[Ȇ|�7�#577�ٳgG�ۺu���A�e�g�X������\�2~�x�6�Z)�9�\c�_�(��L��L�� ����u�dV���;�q�t�4���K����E��q�~�)�&�Q���!�3�Mr�����w�!)w�1��fp��?	@R::r����>��� b���e����(Z�9g�+���,�P�F��q��utJ��8�m���vD�s!�ľ�^*�C�Y�'Z�.ܒ9�FS�@�Q	!7A�%Rcu�礡rއ� f>J�"��H��y XE*ǲ����y�G�<�_�7�\c<x��H��F�]?hР�ك��I�
�V��0�Yed�K�"��t�*�@t�e��G��'��=R��]r�V���+����l�C�� v��p�"�\l��U������Q�w7:nY���K(�3^X��&8�w��{R��)XR�]"�Q>Sk���o ��Y�����d=�"~�w�H���/w655�����Fyk�u���!�*�`�$(���<sD��$Q�,i"xL��+��2T���J	�?K/-�1��	��lժU*�XGG�ÊA�����-_4V���`�RVO�. �"�a�g<)��G���{!
l}���M/R�3�B@�UI��u���� K�;` ����9;�0�~L��K� �〔����}��n����5����!r�r������Y͌#
�������ߩ����J��(�/1BQU�KJI*rgk��yԨ�!]]}䎞���<Y��5v��PI��`;3��2���pPduA���2����E8�pv�=GV�e��ұ�*͓�r#J�����ڶ��/��/j��o +F'N�Â��ޒ���t�ia�� 9�!�� )����刣=@y�Z��=��v3�>�_*3�N�eVF�hA5|�BHƜ1N�a�EoE8��g�k83Ɣ�7���[]��_�>X���o{^`v�t���]I�>�Cp`��Nu�ݙ��4���	�Ń߰{�nD��~%pF�7�a̱�鐾Lk����+����~B�|Ѓ�P�QP����]�CX3��y�$��ve���YQ�:�Y&P�~A��1>���K�3@��Uro�|_V�����!�Dx��%����d����55�B�ڤwM%3��B��*��]��v:��ń���th��)� 'e9�&��{D�%��,�*�G� 7�����zC�I_�]*�Dw�9|��Ƭ�x���Ms��Ɖ��W/����4
1Ȓ��݄(�<ĩB��;d9����b���d�x�4�����m۶�<s�̗:::NOz=�B���LT"�h2�<�?��pa���p���`89�>wn�K�"�-q�!�sF������b�8��C�Nj;v�g�3N�ed���a�{GD�bq�a�{��:��}R���#}J<�(y:����Mc�B���:b��$	;�#C�Pw����j��A�gI�G��&�,�mH�ަ�B
E7���I�
�����I(%X��g$��i��i@p�/�!�p�W�=���1���u�&�����m�__`9A��)�:�����jڪ���C�ꦯ~J{�E&O]de����=�S���eM�3{�}M����Ʀ���nu�(#�&����� ! i?��ܻ�y$���#t���ߥ��qqi'(�e���{�[�|��;�3G_&pyJ�ǩk�����U�Y����u ����+4
]�Hð��`q
{F9�]��}�ɞ�"�(L\�
����?g%�9�¯�K�T�Ǝ��w�� l}�t�H)���l��kG�v,i"��G؃��w8��>���$LF�~��#Jc7���r�.A�ϥ/݌���PPV���KAB=�_�%�+T����Z�n�,�rѓ���1�6�Db��2��GXRE$�e��Z��:�5��:Y�_�K�����}�Gd�b�"�������,�P٪��M Xn�C�9~A�<J���z^:���ۢ	��~�_ �p�,4eN��3�}��}ǔer��C�<A��GD��x!z�Nk��HE`��3o�8�4�M ���A��_��k�=d�8"%sB�[pT��?O�@g ��o�3���.8�b�W    IEND�B`�PK
     uK\��e e /   images/48caf11c-09fe-45e4-9b76-5b0bfa123a56.png�PNG

   IHDR  �  �   U�%�   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{��w}����;3�l]F#䛀n��BPhc,��C�f�R��I�n!����?���l�M���'[X.!���#ۃmᐬ�%���Hؖ53�-K��}?���`�`ْ�3����������~?�^�]     gԎ�9����P��s�ƒ��_[S�J�y5�9'����+s�Ѥt'�_�%�IR��%ud�q9���3���Lr���d�=�2���}eE�U��C�����p����'������<���VI9�-�$�]ʑ���:}�o�I��S}R��K=ܧ�=���l�}����钮�͌��#3��V����o�    ��QZ     0ƇG3��d�ڡ��Φ��ҟק����.u�OY[ҟ37 �ꒌ$u��)��:7_�ԵIJ�.�%)k������r��A�G��SI����&u���$�pM=^R��䡒2�'���K�Gjr��;<��u�K=�g�h�:=��G��]�4�    ��     Ҏ��X��+�]�tkK��}�*)�%uMR�+)����ɪ�����%Y�ߏ%9/�9O�?�E��I�N�PI���h?��hI�&u��I��:w�K���t��L���>+?����cM     ���;    ��׭�+ו̌%�X�.��%�XR�΍��ړ��������dmM�f�ת�?,�DR'�pR&3w����չ��I���#I?Y���2y,C�g�Tr���?    ��b�    �]����>���)j�o�k��z9�8��:�0�W���q�T�ɹ_e*�O>W��\I�d���Ƀg��d�i:    �d�    ,�ȥ���>�c5u,�c}��K���\WKrq��I}ZRV�����+�dR'��?)��s�����K9PR&�O̺���   ����    X��Wn���ǎ�k���zr�����ɯ��qUX�F���>'��s�����K )�����I���     ���    XV���G2ta�zqI.��E%ec�5�P�I����Umk�z"���<��`I}��<���k�׺�>��HF������l�b    `y3p    ΢+6djC�ٱA��%e�W�K��k�Ƥ^��IYѺ�L&��+��k�5eI9PS��8y~�P    `i2p    ��g��s�d��]f7�'��I�J��u���I6&�¤t�s8�jr�$�I�'9PR�הI&k��.�@���ә����    ��a�    |�h��u~zR��O��zaIyzM.(�ƚ\X���[XI�O��$��rR������k}ʽ+2�Ճ���Ij�T    `!0p   �ec|�h�7>zu=)���M����I�5�`y�Ir0������?PS�'u�7����R��m&    p��   ���cņLm����I�))�J���uS��I.�`�:>w��('��59PS�'ݾ�8���o	    �f   �"0��c�Ȧ��TR6���l���zq�g%�k�	 -��XIݟ�}sC���O�ץ?Ч�?��_8����    �;w    hn|��m��]�oJ�g��}�3J��'��x Θ�ܛ�+5��I�夿'��լ��p>|�u     ,g�    0{�=)���M5eSR7��u X0{����S�%u_��[���ݗ�n�    K��;    ��+G3�1��ƀ=)��܀�IV�. Έ�$�����7������KI��}    ���   �)�22��g>΀}cR/Nʦօ @k�D�{��{��/Nf�t�B    X��   �չ�9�5eSM�=7Z���ܘ��I�Z7 ��I����K�=IO��K��s�W���ց    К�;    ����ϱ��_��%�:w}���\غ X�f����]}�[��=w�}x�tvݓ��   ��`�   ��ed4c�Lf7%eSI�9)��]bϳ�ҵ. x��|�̍���)��Խ%�~�Pn:�:    �$w    ��l�2��O��Kݔ�M5uSM6�de�> �y0�d_R��ԓW߻}krlｹ��q    �d�   ���f�X2�)�O^c/��zI��%YӺ `��M�W���<��{������KI�ց    �x�   X v�ˡ�<�K}nMy^M�_�F�Ok] ��ԣI�BI�|��%��]��j�?;�]ӭ�    X��   �G[FF3��.3���Ks���$9�u  �L����]S����A�~(w<�:   ����   �����5�\����  x��   ��    �Cv �e��   �3��   �S0><���3d ��   ��   ���  �U�2|/ɞ��|�`vi   ��`�   �L��˞Yӽ0���~sR��d�u  �Ηk��.�tR?]2��C|>��m   ��2p   X�Ƈק<���E�lI�$6 ��e&�_H�=I�S����SG2q�u    g��;   ��.��J�wj���^RS6�=���m  p�H��$wה�]��Pn�l��u    ���   `�ڐ+7rbKM�RR.��7'���|  Xv��|!){���${�͚O��G[�   ����   `�;?�O�<�$��~KR�$yQ�U��  `$��s���)�{���=�]�Z�   ���   , r�ƙ�\27f/[��yAR��m  �DL&ٛ�=I��&wOg��&7o   ��;   @+eM�=o8�Gjʖ��(sW��Z� �rS�c%�;ɧJ�A���y�1z   ��    �`C��8ȉ-sc�lIri��5�  ��٤~>��$uOI�L�ܿ6z   8��   ΰ��׿��Zw  �m&�_�������<�:   `�0p   8��:�o)��$[j�#%��u  0_ꉤ�MRw'ݞ.�s(�}6Iߺ   `12p   8Ec�>���PM�$eK�oI�%��  ��H��$u�cF�{���a    ��;   ��ؐ��2��o��`�{
  ���'/��   |>�   ���3�z6yѷ���t��  �%m*�ݏ��kwL��{ZG   �d�   ,7�iy�)?Z�]ZS/M�%��  �qoI�����K��P��Dr���Q    ���   X����'��dk�M��u  �)�M��KrgM��K��mw��   8[�  �%e4�7��&���\��v�  Xb$ٓdOM�\����]���   8�  �E�uv  �$��   K��;   �h��  p�\y   %w   `Ar�  ��r�   X�  ��uv  �y��;   ���   ��K}I�]ާ����4ɺ�U   �[=QS�t��r� ��#����U   ��b�   �urٚ�����lMrYM��de�.   �Hݗt�kr�P��Pn��u   ���   g܆\~�L��s��rYR8)]�.   Nہ${jrgRvM�O&�[G   K��;   p�F�}S�`kIY��_Һ	  �y�P��L��&w������GZG   ���;   �du���e]���nK��u   �l�O�dWRw'#�Of�t�(   `�0p   �����9��o��+���u   ��l�O'uwM�,)���T�(   `�2p   ����h�K�֒rYMݞd�u   K� ɧ�׬��p>|�u   �p�  ��w�9c9��j�˓�,�K��j  ��pr�^nO2�gŝ�   ���  ���ch4_����+���u   ̩�J��Ovu�y2��[   ���   ���lߔ�w�������o�   �`6ɧ�O��;�����   �w   X�6��g�m�����<�u   ��z4)�ɮ.�=��e21ۺ
   8s�  `	X���J7>7h�֤\Һ	   ���$�ɮ���m�HR[G   O��;   ,B�U�r�ғ���I��t��   ���J��}����<��/�   �w   XƇGS^���en�����h]   [�W�]5�[̭_k]   |o�   � ���}sО˒�ۺ
   ����܅��LL�.   ���;   ,�پ)l��5u{���M   ���|����trg2q�u   ,w�   �Ȇ\~�l����W��+�\غ	   ��z�$w֔�K��'s�ߴ.  ����   �����d�܅�lO��xo   T����h���������   `9�!:   �E�پ)l���W%YӺ	   x*�ޒrC��ιw$7o]   K��;   �Ak2��K�v�J����}��   �3�M��j�+)��s۞�E   �T�  �iK��O^UR�Jꋓҵ�   �՗J��5݇���u(7n   ���;   <I�s�C9���5I�&�X�&   `�$�T�k�ӹ�Ij�&   X4�  �	������$�&ɋ�=5   pJ��I������LL�.  ��̇�   �8\i   ���  �	�  @W�  ��W�/�>Z���g��  ��  X�V���3|uI��rU�u��   �ek6�5�����3��A   Ђ�;   ���l�<H��$ۓ�'n�   �x�)�Ir�dλ9��x�    ��   ,i�ȥ��9����$�uI�ٺ	   �ɩG��$7v��Ľ��   �l1p  `�Y��gՔ��d{M�:���M    gN�[RnHr�d&>��o]   g��;   K�������$��䚤\Һ   `~����5���|�`vi]   ���  �Eic^s�#9|E�k��ז��M    ��&�x��]�?>�ۿ�:   �,w   �չ���_��I�LrN�&   ����-)7$�q2����E   �D�  X��g��A�5%yM���{Y   ���~�$�5ɍ�9���㭋   ��   �����&����.)�k]   ��ԣI����0��C��Z  ���  hn}�^[�ȏ%�u5�IF[7   ,�I�H��ө����A   ,o�   4�&��R~,�;�\���M    Խ%�$7Nf���5   ,?�   ̛uV�OrM��$�-{    �����?�)7L'��l�    �>w   Ϊ�ٶ����~M�-�{    xJ&妒~�dλ9��x�    �&w   ΰCcy��$���H���E    �I�hRnM�Β�Mf�t�"   �w   ΀��˱+j��L�k�lh]   ��8^So)��h��CGr˃��   X��  x��W��^Y��H�k���.   ��A��L�s8�?<�;�  `�1p  ��=#���pVl���?�����    X�j������?:��{[  �8�  �=m�k�{$��8y��uIV�n   `��{���O��ù��k   X��  ���:V2��Hre�sZ7   �T̍݇��0�k]  ��b�  @�dM�xZ����5�I�[7   ����$e� e����Z�   О�;  �2�����UIYѺ	   ��j�� ���   ˗�;  �2�.���Z�v    �G��C�w$�|�u   ���  `��њ���   ��̍���8�ۿк  ����  `�ژל�H_Q��H��L�y��    ��<:v��g⋭k   8��  ��sժ9�ښ�S5yeIV�n   �����j�e�̭_k  ��a�  �����J���Iִ.   ��S��ܕd�lV|��|�"   �:w  �ũ��Kkꎤ�>����    `$�˚�ޡ���C��p�    �w  �Ed}�m�����I.n�    UM��dWRv���?�/7?ܺ	  �'f�  ���϶�}�$?��9�{    `�GK�?O��M����i]  ��3p  X�F�(�!�O'��=    ��<PSwv)����$�u   �d�  �@�f�X2����1�K�=    �m_M�$�=S����c   0�   hl|�X�IwmM��$#��    `y�{��3�{�2��5   ˕�;  ����2�Ҥ^[S^�dM�     �Q�O�]Iv2��#����E   ˉ�;  �<Y�m�k�}�%��u    ���XIv���N�%;O�n  X��  ΢�l��>�����[�     O�TRn��Oܒ��  X��  ΰ�lK��AI}cR^ں    8��I�������[�   ,%�   gĎ��<����1�2)�.    �Ş$�$8����c   ;w  �Ӱ>�6��kk�sI.l�    4s<�Gj�{��П&{fZ  ,F�   O҆\~�l��ARߘ���    �z�$�%)��ĝ�k   w  �S2�r,�ʤ����D���E    �bP�&egҽ{*�~�u  �Bg�  �ݕ��_V��Kꎤ�m    ,Z��|�K}�dʟ$�Z  ,D�   �fC��8��kK�I�ۺ    Xr�K�$�}����u  �Bb�  �$�����*鮭��K2ܺ    X�j�$�Y���d��{   Z3p  ���ٶ��^[箵oh�    ,[�$����s����'Z  �`�  ,;k���%'�ǒ��$?ܺ    ��L�ԝ5��S����c   擁;  �L��ۺ��j�O$i]    ���ޚ��A�����@�  ����  XҞ���_L�I��u    �SQ�cI�4��3��[��   �
w  `	_9����r]�+�    ���[���S��R�  �3��  X2F�mKI��$�0)�[�     �]�Oʭ5���<��ɞ��E   ���  X�Ʋ}���Jꛒ�p�    �j�����%�w&3�{   �*w  `QͶ-]���ܵ��Z�     , {j��+3��r�íc   �w  `�8?��H~�$���9�{     �z�$�ߧ�~:��i]  p*� �����+���j�O$i    ��)ׯH��2�P�  ����  X��y��^��M�{     ��#%��}��5�[?�:  ���  �k�     ��Uw  `�1p  �[�+.���J��@�    ��.����wN��O��  �7w  ����oMʛk�Oʊ�=     �]u_��ܗ�n  ,?�  ��Z��.��ϕ���9�{     x\SI�_�wMf�o[�   ˇ�;  0/F�mK����rm�s[�     p��Ԕ�������]���  �6w  �9?�O�����r���    �t��Kʻ��������  �&w  ��[�m�N���\�d�u     gR�rkM�~:�q�sк  X:� �3dǊ����%�$W��    �����w��r��c  ����  8-r��3zcI�i�g��    ���%�����3��u  �x�  O�XƷ&��5�uI�[�     �P�O�t�Z��ܗ�n]  ,.�  �)ې���d��Kꛓln�    �BV������~0��u  �8�  Ohm^�ܡt�P�_J��u     �I�rkI}�d>zc�ں  X�� ����+J�$���     ��/��w���s�d�  `�1P  ��X�����\���n�    ��t��~0)�~2�:  X8� �$��2��A�?I�/$Yպ    �ecwM}�tʟ$��c  ��� `Y�14�����9���5     ,k_K��?����1  @�  �������j�/'yz�     ��z�$�/��q(��ݺ  �_�  �������?M�I9�u     <��5��ӹ������1  ��g�  K_7��W��-I^�     X|�{M~�$���T�  ��1l �%����>���-I��u     ��z8�{��Oe�K�c  ����  ���r�lf�K�?K���=     p��>)Q��OgbW�  ��1p �%b4۶��-I}}���=     0O>YS�9���d�X�  ��� ���ed,k~���jR^ܺ     :��?�w����1  �Sc�  ���\���#?�Է&��Z�     �r<)إ�ׇr���1  ��c�  ��h^��.�/�䗒,�kz    IDAT�k�     W�rkI}�d>zC�  ��� �"0�m[J򖤾>�p�     Xd>��ߞ��&{fZ�   ߝ�;  ,\�X^����$�[�     �p ��5�o�Ν��c  ��d�  ��_}"�]�[k���=     �I껓�7�[��:  �&w  X 6�ʍ�̼�&�%k�     ��lI�h��o��:  0p ���f�9]�?�)וde�     X�v��3��ޘ��� ����  Ͷ-%yKRߐd�u     �$�ۚ��SߛLk  ˍ�;  ̯n,/uMy[��Z�      ��&_/ɻ���T&�Z�  �ra�  �bǊu9��I���\Һ     8U�p��e��z0�~�u  ,u�  pm�ekf3���I�Ѻ     x�ꉤ���~������5  �T� �Y�*W\8��?I�$�Z�      gJ��]��8�[?ֺ  �w  8����R~-�&)+Z�      gS����7���$�u  ,�  p������֤�!�P�     `^�MR~k*������1  ��� �i��֚�-ɫ��5     ,w�$y�������H�  X�p  ��+cy�5}��Z�m     ,4�����$�=����5  ��� �)�2�.k_��oK�%�k     ���I��x _o]  ���;  <���Y�c?���")�Z�      �M}$��t��u(��u  ,d�  �]l�ekf3�j����=     ��7H��e���϶� ����  ���\~�P��ZRߜ��Z�      KM�I>T2�/&s�gZ�  �Bb�  '��U�د&�WJ���=     ��WR?6H��ù��[  `!0p `����9��t?S���=     ��S�6��<��]�[  �%w  ��uV��7��וd�u     @M�P����u  �`� ���:/�������<^     PM�/�}:w�+Im�  �Ř �ec]��'�����m�     pj�餾c*��d�u  �m�  ,yk��kK���d��[�      <5�#5����&7o]  g��;  K�����.�o+�к     �L��g����{ӑ�9غ  �4w  ���y��~[���$�kZ�      �}�g��������� �3�� �%aU^r�p��U2�ƒ��=      �f���������Wn]  ��� �EmU^�t�g�ȫJ���     ���>3_����G��}��l�"  x*�  X��Uy�+���z��e%í{      ��>����Pf��T>5պ  �w  �眳6�~����dų�     ��>�����ݑ�ߜ̞��. �Sa� ���:��.+~9�~��9��P�$     �E�O����?)�oΞ��. ���� �ku^��d��d�vY���v     ���O�����VR������$�u  |;w  �5ٲ5��J�W��S�     Ό�>5'R3�Œ���Y�d�X�.  x��;  E�&/~u����Ғ)���      g����xjf�+)�,9�����d�.  � ���+��ܟ���<)/�"%+ZG     ,5���g���݃��#�����  X�� hb}������|M���{z��v     �F3t?��?�����|ro�.  �w  �ժ�䢡�7�Է��u%+R2/M     �{�н&��>���_�j� ��aE ��X�-?ԥ�OI�ْ�d$�a;     �5� Ǔ�dOIy��<���A�0  �8k"  Ϊ�����ג򪤔.+���B     `��ϱ$}�|.)�u$S�O�x�q ���޽�u��}�>k߯g�.IH$(��	27I�$���L'����3��&�5��ز-_dE6-ۑ#;��؎�I2ө��t�������i#[ ٖ%� 	$@�������8�1H� ������̬���k=�S u��<��_:��I�$i7�O~3$?�!ȱnw
*I�$I�$I�t���A�!׃�W�72�_��\s��I�$�1]$I��YJ����~x�F�=�'8��$I�$I�$I:�"#"c�Vн�G�g����y�&I������$I�f��B���?	� �%��SNI�$I�$I���&�2"@7�oOI~���_�sq�$I:�LI�$鮭�k#��G�Sp#�^ ��'I�$I�$I��]��������񜋓$I�e�]�$I;V�c	��Ŀ,2׃��'I�$I�$I��=���G[1wH��ŗ~o��I�$��1�.I��;��#�!��a+�(�K�$I�$I�$i�HdDdt�����<�?ϫ.I�$,�%I��<�x �Q�`{���[I�$I�$I�$麔�!���;�M�m��V�wI�$��K�$�m�y��H�q�?���1����-N�$I�$I�$I��[���D��w���AwI�$݂wI�$�E���4���s�@B�;��$I�$I�$I��LI�<��?�&��ϩ4I�$�Cf�$I�����?|��?y7�]�;}�$I�$I�$I�݈׃�C�t��WZ��|a0��$I����P�$I��hB�$�o���@���Q�$I�$I�$I��2��o��J~�5���S�$I���J�$IGW���7?��7|@�@�@2��$I�$i�r��|�R9G��$
�7��R��� ŶL&C����6�g3�rw��>M#���m?�L�����~>MI'o�c<�2M���?a�F�Ӕa����$I��Hd|���\�_�e�s�yT&I���r�[�$��Ij<��"������`{�@f^�I�$I:�B�R%O.���g(�sd��\.K��%�M��>�d��,I&��m�`��%!	�!�L&B� ���yI�$c$���ܛ��S��㟼�L&�F�)I���3���`D�d�L�L'��$e:�2LH���h�h8e2I'&�Ƞ?f43����Z�$I��I��k�����6���9'I��90�.I�td���	%x��O�����%I���&���9��<�R�b)G���X�Q(f���l�|!!I��V����d+h��zM�
���q+S�10M �42L����ӭ��p0a�3N�~��'�{cF�)naH�$IGMJʐ�[�mG��H�L�߿2��$I���\�$I:��W)}g ���7~H��ϣ0I�$I3��g(Wr�]�3�@���T�
��Y�����q��z6H�\>��]�g&�)�q�d��S��t���`��|:�L�0�����c��1��NkH:��?�$I���3�tˤ������:|��
�$I�q�B�$���������7~�H(̥2I�$I����T�J��vh�T�R,m����B�\~+���b8]z��V@~4�0NSF�)��V��~wL�z ���m�H��N$I���!2!e�oz��[)�{<��\��$IҮr�V�$��y,_����:������$I������z�b9K�V�Z/luT/$d�\>C���Tʑd!I��K�ts��A̰?a<���S��	��vs@�5�ߛ�)^�$I��)c�t���)ӟ5�.I�t��["I�thl�x�͟2׃�9�&I�$�,TjJ�,�z�j�@���T�
��J9��@��%�s�-���p+���&׻鴆tZCZ�C���̻\I�$逊����n��AwI��Cƀ�$Iҁ�N���z�=;��$I���!�OXX,R[(R,e�Ts�������R�|>�/f	�eUI;7�L���FÔAJ�3�����k}ҩ�?#I�$�J$�K�$z��J�$X��k�3?<��O�@�@~�K�$I���$�EK,,����y���B�|!!WH�d�,iH�Ƞ?b4LS�	�ΈNkD�5��9dc��h��/I��#kJʐ��V� ��	�O��w��ue�$I�w�%I���۷z�灼�=I�$r�r%���2�z�J5G�Q�XJ(���Y*ռ�%J�ɔ~wD�;f8�0�t�C6��tZC6����)��$I�!��2�[}l�]�$�rgG�$�����4p����H(�4O�$I_�\�So���,.�(�
Kʵ�J�B1C�8����3���Sz�	���^{��z���>�k}�)�� I���.2"e�[}l�]�$�q�R�$i�;�������,�<���&I�$ݭH��gq���R�z�@}�@���TΒ/d�d\����c����M�w�t�#��!���k=Zb��v�$I��HʈȘ�ݧ�O�8wy���$I��")I��o���	%8s�s
�{Z�$I�t'�YXX*��\��T��(R��(���C��c%i?K�H�է���N�G�6�t;c:�kW��l/I��}(%eHdr�O#�ߊd��_���$I�t'�K�$�?I��9����)��<�N�$I�4?�r%���2������Z�B1�R���UI:�&�)��V�^wB�5��1��1���6�a�uI�$�KdBdDd�v�t���0�t�?����$I��\U�$I�?B�'�§���I�I��TN�$I{!���r��5�VJ,,���r������RI�[��v�:cz�1���ƀ���^�2G��K�$iD"S""��Nj��a�����=,N�$Io��'I��}��������;'�!P$��ei�$I:"�J��c%V�WXX.Q�f)�3,4�ds%I�5�in�h�F��[��ƀ�_k3�[X�$I��Hʈ��v'�¯e�|f�/���2I�$�����$IsT��&�g >�v�ٽ,M�$I�P6��|�ı�5�y���F�j-O��|S�4i��t;#��	͍���4����� ��J�$Iw/���ow�*��m�
�_�J�$I�M�K�$�A��� �oV !O �w�I�$���d��\bq����2���Z�|!P��%AI��4����}��!�ΘnkDkc�믵h��>�N�$Iw,2%eLow�U�3mj��/��2I�$�wI��=U��?��?{��y�8]�$I��I2)+'����t���b�j=O��7�.I:r��1��vs��z��k=�]n�n�|*�$I��VdB� ��9�W��6�_��Yq�$IG�;]�$I{��S�'ğ��m�;/�%P��$I��%8v��ʉ� {�Q�\�Po��K����1��]ڭ��!�=�^��i��K�$�HʈȘ�݁�!>���o��n��]�$I��0I��]T��A�qn�ZOH(��*I�t�e2�r_���囂�YꍢAvI�f�V��k���[c�y�'I���HIy�&��g;���^T%I�t�3&I��J<�`����n�Zr$�qj&I�t4��;Qei�D}�@���R�d�$iΆ�1��>���ƀ�k}�]n�nM|�$I��I���������uI�$%�I�$�P��+��~(���@�@���L�$鐊����α��,��Xh(�3�%I:`��k=ڛC֮��v��ڵ�n��>I�$X�)# ���@�����M����T&I�t���&I�4+��ڐ��?�ov������$I:D�;Ya�D��r�ŕ"�F�r�0��$I�.�N#��.k]6V�l����j�~wJ���$I�t�DRFDF�|"����.�~y
�$I:��K�$݃S�-w࿈[���;7�\����$I�AV,g8�@��KE�y�Kd���(I����v���ڀ���t|'fpkN�$頚�2$2}�� �C�or��^T&I�t��&I�tW��j���3��w:;�'!��/I���$R_,r�����Pk�)W3�%Bp^'I���h8ac�C�5��9�ڕ.���d:
�^$I�tpD&DD�;�:��;S�'z����I�$&��I�$�LR穿����N'2��ݯL�$Iw-���,p�5�O��7
TjY�9��K��ݑ������}�CV���|�Ű]K�$I��")#"cx�{7�n��/����'I�t(p�$I�C��h �� O�ӹ��@�@v/J�$I��$��}UN�_c�x��R��R�L�0�$I��^w��Z�͵�/����&��V#I�$�')S���NN^~�M������%I�t�p�$Izu�~:�~�swr~ OBa���$Iҝ���zp���%�Y>^%ggvI�t@��\�v���ڀի}.��b2vz�$I�"R�@������js��s�ݯN�$�`2�.I��6j����������)��޵ݍEI�������`��eW�4�JK�y&I�4Siint�X벱:���].��b:�ڔ$I�DRFD�@�����}n��$I:��K�$�I�'���
�! �N��"���'I��m����^���
��J�r��%Iґ����f����}�]�r��M�I�[��$I{%%eHdr������ڜ�v�,I����,I����Xu@�����w:k"�'!��*I���U,gyי%N>Pci�@u!G�h�]�$�v&�)�6��\���������$I�vYdB�H���@��)�u���ne�$I�I,I�$��j���I�ĝ\ȒP��$I��ER��y�K��,�YZ��s/I��{��Y�֡�>�ʥ_�d2N$�.M�$鐉DƤ��x'L ��)�=�]���$I��5w%I�Q���� � g����]�$I�f�P�p�*���|�Dc�D�dwvI�������F�kWڬ^�q��.�.w����(I�t�R������ײ��皻[�$I��䪔$I:�x�?L��|�N�	�I��J�$�^D���x�K�J4�vg�tK!2� I��$[���٭�3��[޻��L&C�׾ٍs��Ͽ��b�L�ӷ�|:���w�Ln~HӔ4M�0��֍�b�ۯo���{���K:�n�����m^yq��8�u1I����﬛;�j�O���ù�n�&I��߸
%I���*O�?!�l�o��k��]�}L�$I�Nmug�q��+'�4���vg��l6��f��a�}���lv;~��[ӵ�n���ۿ�L&�!��dr�����>7H/|iim�X��e�J��_�p��.����#I��7�����vr��#|�ù��</I�t��K I���2O�ʐ���9���[ \�gw�:I���"r�T�߽��SUKy*��AUi�!��f��\n����o����� ��M�n�����9<�q#,?��_�x�v�%�ng�����W^���&qj�wI��;���w�/B��6���ݪK�$i�p�I�$j'�P�G����;�.�#���%I���)�OU��t�㧪,/Q��]�th���L��r���*��$>�J_��m�7^��㷼���%��d<e�Z��k}�]�r��:�>>Q�$�6"R�1���Z<��.�%I�4w&�$I�a��y��#����;�,C�w��]�$�HI2p߃5N���r���2�Rn�eI֍���l�B��\��k6�%��S(�߷{�ton�?��F�F�7���)���h�x<&�M$]���ի-V_�z��+/n��F��n�$IoI��1�߉�~�×��Ve�$I��n�$I:t*<�ф�3����@B�@~��$I:hr����u�{������+��y�%�K!r��|�\.�����#�Ͽ�=����0��p�ÿ��ay��K�cds�˵�;�]����MZ#�$I�E�DDv��b��6����T�$IҞsE�$<y6%���vr] GB|\�$I:����jp���+��W�d�#�h�9�^(����A����B���$`�K�h4���C���7�/u���^o�v��k���v�K�'I���-2"e��Ӥ\��O�y��`g	yI����I�t�����L
�w���zB�"�%J�$Q�z�jp�@{c�D��\��!I�7��s����������cd<�!�>�������Cb��`�t���C�]i��z�+��\�؆��$I��I����wz�H�[��](K�$iϸc)I��%��>f��ŝ\�(8�$IGJ�����.s��:KǋT�wu8��U�P(P,�ҁ=I|:����F�����C�:���W���z�˥7Y}�O���$I::""���_�?A�G����F'ϰ    IDATQ�$I�n3�%I����S���N���@�@���F�$IT�x��<�P�c'�4�J��r��l6�Z�9�~��璎�7���vw��`�x<6���n�_�����k#�$������vz���D�?��k�Q�$I�nq�G�$(U������;�2��'��)�$I:����`��7X9Yb�D�Lƹ���vH=��S,�����y��2�Lf�eJҁt�����h4�������KIk���W7Y����t�S�$I�a5e�������m��_�$�pJ����G�����m;�6�%� vm�$I�L�DN����������R"�5У��F��T*m��o>r�ܼK��#-M����`0�>n�>M�y�(�Vk����\���寯3�E\�$I�MdD��������}nʒ$I�)�$i_[���)��(����1Œ$�Y>^��,q�t���"��s�/�l�b���{�T�P(�K��tPM&����o���!1�8`#�#�W�\���m.��d:�=*I��HJ���n���1%��.�~y
�$I�	Wp$I�>�M����)��N��I��tG�$t���^��w�Y9Y�T�õ��v]�K�٬7]H�Qcd8޲�{��g:�y�F���d���^}y��_� N��H���-2!2 {
��~��_ߍ�$I�/I���Tx��	� ����@�@�ࣇ%I�U��8�ex����"Ų���Ri�(��ہ�|>ovIҎ���7���>�^���f8s��W^����֯	d�]�$I�]�������N ���_�/f]�$I��r'J�$�5�>
��/���@B�@~�eI�$�"������48~���"I⒍�F6��R�P.����W*J��!vIҞ�L&ہ�^�����z�i:��tD�6{\y�ɕKm^za�Q?���$I:P"����w>�p�O���?�����$I�5w�$I���8��S�v�&)�%� n8I���Z�s����U�ĩ
��7�i�d2��N��b�r��}d2v)�$�_1F��!�~��`@�����>��܍vG�F�^���W6��J�˗:��ŭUI�tDF���˜���~�Ǘ��qY�$I;�*�$I��o��h}��Vv~�]�%I���$p�t��޷ĉSe�쎭�
!P(���J�b��j�$鰉1����v���^�N��t:�wy:dz�!W��x���x�A��K��}-��2 �jn�B�g)�����g\�$I�q'U�$�E�'�| �]��ws�V��"Ng$I�~�|��C�Y�����J��v�ֽ�d�T*o��^�V�iB���&�	�n�^�G�ۥ��|���Y���ڕ�]hs��q��wY�$I���拏�&�m�^ζ6I���s�K�$�Ξ��L�o��2 7�$I����gx�#�<���'�4�J�.I���+�
Ib�PI���h4���8��^�c�����׺���:�����%I�>�2eL�v���p�s�|�EI�$ݖwI��'N�J���D�ǀ�݌ȓ��)�$I�/N�_��G����:������\>��V�d�$iN�kVb��]ks��6�.������%IҾ��2�.����2%�`��2��$I���]WI���B���
�r��w5 		E 3��$I�v(I��#�<��%�{�B���wI:@��<�J�R��ݙ�V�d�$i��U��n���K�1Oy��&�������i�vw�$IsI�� ���'�S�|�5��$I�nf�]�$��<�¯B���v����Y�%I��#�j�w�g��/p�T�|����L&C�R�Z���W��$|1F��>�N�n�K�ӡ��0��]���#�W�\�����M^{�C���$i>""�]vs.C�D�g�PI�4s�%I�̕9{_��	��wג(�!P���$I����Eμ����|�B����[��+{�V�V�Q*��g$I:J&��v��n��t����xׁ!r�f�˗��z���ϯ�N��u+I���=ws8��|�_Ϫ*I�$p�D�$��c��>��f� 
�3�L�$�v�N?��C�Y���e�u� �7
!P*��T*��e��*�Z�|�y�$I������6�v{; ?�N�]����x��K�\���ů��i�6��$I{&2%e�=4b��?��8wyv�I���̀�$I��*O��@�U౻#�!��]6}�$IڑJ-���]��3u��W&��̻$��L�j�J�\~C�=I��J��{7����w:��.��`�ei��1�z�͕Km^9��k��	d�]�$I:�"�k7�n �r������@�$I�%I�=)����d���w?J !O ��I������y��˜zW�ŕI�����r�j5j��J�j�J�X�wY�$����a�N�C�ݦ��ϻ,��f���;��r����t⍹�$i�D�DĻ���| ����o��K�$=��J����X�N�{#|
���(vm�$I�)�I8��
�o�c��)��e7:�W*��P{�\�wY�$I�4�N����������]��h8��+�v�Ë_]c��{%IҬͨ�;��3�?��sfP�$I:b\�$I;V��&��<z��ص]�$�\>��]g?U&_0�~�*�^*����$I:�&�	�n�V��}���y��9�1r�J��/n����m���H�����2$2��"��/��|^ΰ8I�tȹ�'I���g�Dx&·��8�,	��.I�f%W<��ez�"'NU���%!��*�Z�j�J�^7�.I����pH������n��L&�.K{(��뗛\��䥯m�vuH��D�$i6"#RFl�v�k_����K�bFeI��C�]>I�t��Tg��H�P��qntm�Ϭ2I�ttU�9���1��H��cE2o�;
B�J�7�k�I�߿$I���h;���th6��ޏ������΋_[g�ʀ@v�%I��.^���=ts���	�����^�AY�$�3�.I�n�Ɠ���C�2N K�Hp�!I��A������8}f�c'�$�s�îP(���@�V��f�$Iڙ#�~�V�E�ݦ�j�����p� hm��|��K_��ҋ-�vv�$IwoF������-�� _̨4I�tȸ,I�n�Γ�ĭ`�_�����.I���ұ2�{�8��,P]����U�J�B�^�V����@�x�$I�ۚN�t:Z���1��]�vQ����.����-�԰�$IڹȔȀHz�C���7�<��Y�%I�w�%Iқ|c���c��c@���ʐP�k�$Iڱ��y��%N>X��l�������]���:vg�$I���`@�������v��~H��#�\����&/~m�tb�]�$�Lʐ�hC}>�����߾<��$I��`�L�$m���7C�U�{�F��N7$Iҝ!�G�y�V��t�|�9�aB�T*����ݡ�\.ϻ,I�$�ƛ��7�M&�ɼ�Ҍc.]�����6����T�$ݩ)�l����[l>/gQ�$I:��-�$I����Y2�@��{+�!��	"I�����<���>S'_t�p��r9�����%I��#�~��{�٤��ͻ,��t2��M^��翲�t��-eI�t;������~�ɹߝ�`�$��r5B��#�l���S@�^F
@�`�vI��N�_�}����jT��y��!P.������u���˒$I��ǴZ-��6�f�v�M��sO���K/��ʋ-^��:q��wI�$i�׻�s���>?!��}�xi�I������$IGT�'��@���c�:�]�%I�;Y>^��:��G(Ws�.G�(�@�Tbaa�F�A�� ���U�$I[]�;�����]�'�ɼ��=��\���+/6y�k�ĩ�I��V3����3-�{��,�$I�wI���
�p"a�K���
�*I��jq��{;��Y\)ͻ݃�J���E��:d�vo�$I�;�1���i6�lnn����x<�wY�����.�s���\�z��$I�Ͳ�{��{[<�o�2I�tPp�$��H�<���`�އ�����.I�n��\������YBp�� J��Z�F�^��h���@�8�$I�l666h6�4�M���K�]��\|i�/lr�6�̼K�$I�F$eHd&77F����9�:�%I���.�$IG@������Y�ȓ�ǩ�$I�����c<��%�yC�P&��^�o�FÿGI�$��`@�٤�j����`0�wI��V�W_i���7�x�E���$I�ȄȐ8�n��:�o��oqJ���ɝJI��i�d~>�_�Y�ZO�wmwcB����R+�Ǐ���.��R�,��r#��h4�C��%I��_�F#��&���4�Mz�޼K���=.�����ʵ��*IґI��h��G���ṯ�h@I��ϸs)I�!U��o�����Ϯ�$�X��������.���3�~�d�YX\\��hP.��]�$I�t�F����ۇ����6_j����\��$IGWdBʀ5_G��
�x�/wg1�$I�?\=�$�)����d��g3b�޵=;��$Iҁ�$�3�_�}<ƉSe�M��$IXXX����h4��.I��C���kkk�F�y��;�z�Ņ6�ꗯ��Dܮ�$�(J�ws��j��	|_�s�;�%I���b Iҡ�M�:���)�:�Y�8e�$��9�@�|�>\'_�̻���Z�F�A��`aa�@�$I���n����&4�M�ә���K�Ӕ�.n�����5҉V$I:j"#RF̨�;>�2��_�:�%I�\��)I�!P�'2�!>5�	y��'I���R�G?t�w��Am�y�~W,Y\\��h���H6k D�$I�1��t����>b�MhJ�c8s��*翶Ϋ/u z��$IGEdJ�f��}#�϶8�k@:�A%I��3�.I�v�Uz�~
�[�LV�%��I���R9��?|�w=����]���|>����F���%
�¼K�$I���4Mi6��޻ݮ��}���s��:_��U֯�	$�.I�$큔!��,��W��{:<��Y*I����֒$P5���@��#<8��(��b8I���%I���Wx��q��I���(���h4�����uj�ڼK�$I���tJ����w:�y���q��^X�k�J�qk[���m����6^�iS�|a0�A%I��p@�����2$��uVc���v�*I�av�:x����͹$�߄XXX`ii�F�A�Z�wI�$Iҡ7����>&�ɼKқL�)�/n���7���2���-I��Iͺ��	���|��堒$iw��-I����x�!�20����<	y�H�t8-�Tx���s��%
e��7�b���E�KKKd25$I��y�1��t����>b��.K7�\��������M�ɼK�$I� 2&e�n.�s)��wx����$I�ƝmI��
O$!�-�����]۳�R�$��R�?� �|`�r-��G�$aaa�F�A�ѠV��}��$I�fl<o�����f�IT����������4�&��-I���D�D���Z �p�g��,�$I��|I���o*���X$�8��ը�,	E�
H�t��~h�ǟ��SV j�/��.I�$�^���5���31F�^iq�����LF~�$�0��H1�n�������3T�$͐�6I���g�����7�@�]V^�$�Y�Q��9ΙG�(W}2�~��d��싋���y�$I�$i�&�	���������nw�}b4����U^��_l0�.I�aI�f��=B/�'�<��𹙶��$I�΀�$I��"g��� ? $�9C��l��$Is�$�3�_�9���!��~ފ�"KKK,//�h4�;�$I����`������vw�'6�:���U���V�#n�K�t�E 2$2�#<���nr�ٙ,I����%I�Gj<�-~x`���$f9�$I���j<~�>|�F6�W�y�d2�ڗ����}B�$I��-����M666X__g0̻�#m:M���*/�ɋ_� ��F���mBʐH:�A��g�4^�r`I�tw��$i�����F��َ��P�1��$`�R�Ǟ���mP_��|����v�}iiɿI�$Iw����G�3���u����l��񉧒$T���ɬ~!�_�p������$ig܉�$i�B���#?,�t`r$g9�$I�C�^�CO���%��!�@�Rayy���%j�ڼK�$I�t���c��׷��t:�#W�����_y�*��AwI���0d�+��o����:_l�vhI�t��K�4'�=	� �¬���ڞ����$i���|�ɓ�����>^Uw(I��.�������y�$I�$�JӔf����kkk��y�t$��^yi������-��.I��I������ˑ���g=�$Izg�%I�sߔ����?Tf;v�E\��$���d���
��,1l�k�B�����#�K$I�$�^�������4��y�s$�]k���7��_�ߙw5�$�NE 2$2ڍ�??a�=}�ݫ�1�$I�5wl%I�C�~0!�#�O�z�@��<�x�$�`XX*�����H2���Z�\fyy���%�]�$I�$��x<f}}}��NgޑT�1���za���p����$��wI�$�D&�؊���&ď�y��z`I�tk&�$I�gs5�a��@~�c'$]`�$� ��1{�$+'���"��F�$,,,���ıc���g<%�$I��]��)�f���5VWW�v�3����z�/���^gЍ��.I���DD&�1��2!������]\�$��oߒ$�
O|8��N�'f?z����$�k�F���S<���b2�r��\.���
���4����%I�$l1F:��vؽ��ͻ�#c2��ʋ��ѳW�r�O�$�g�)���	�G�<����F��]cN��]�M�:��ğ r�=�'!�?�%IڿN?��G��~��*�:��(
,--m!8W�$I�tx��{�ٜw9GƵ�[���5���5�C��$�_S��ٍ����%�k�<wa�K�$q�$�O|#$����'׻��h.I�~T*�������Ǘ)��ڽ��"KKK;v����y�#I�$Is1Y]]e}}���Mb�F��6N���_��ٻ�0˯����so-��k��ګ�nY�d�"˲-#���Wp��,2O3O&�bH�L�d�'a�0&�NB�I���E��^�Y���nu�ֵu�z�{�IFȲ�V׽�V���y�o}?�?����>�s���t|n/IR�D
Ԩ��'����r��ڦ�$����]��MuwW/�O� �n�O����pI����C��v�8�{��>Ǯ���nٵk��vI�$Iz�r�����W���oan�s�,���sTJ>×$��D*�(P��V?�X�/��K�Ԋ�YK��Iz9�6������ϐ#�^�-I�^�\WG�������i��޺��fxx�����q$I�$iK�T*,..�������j5u�mmc���3�<��W��J^������됚<�ӫ���{��%I�5r7-I�5��X�*��Ǩ�����.�W�J��4�����cc쿮���z	!���Ǯ]�&�˥�$I�$I[Z�V������ϳ��hٽ�b��N-��SK|�K�Ԫ���$�D R$R�ӄ�@��k�~�N$Ij	�%I��g�����z��@;:qɖ$)���,G�|�n��;z�{��Xjbxx����ԑ$I�$i[z�쾴�����r9u�mkm���//�ӗX_�CyI��A�B��W�7]�O�r�_y��$I��m9I�^�	�u�����Q��4ȑ�m��$I�*}���	��y��/��!��000���0�v�Ϳ�$I�$��b�\�r�����uT�F�/\�K�g�:�F.��$IW�F���u��o�SO�k�$IەwI��R/��
�׀��3!K�>ؖ$)�}�vqǛ'���i�uB`�Ν���044D6�MI�$I��_�����YXX�R����--̭�'x�yjU�Ē$��H�H�^#
�O�r�_z��$I��wI�^���z)}�1��>t���hI��hk�pˑ	n=6JW���f!���������ttt��$I�$Iz1F������gqq�j�N�f�X/r�+�<vb����$IJ#R�F��+�������З�4@��m�ݱ$I�A/G�̯��gB C�@[}~�$IzU}�9��y�n�I��x����0::j�]�$I���Z���˗-��I��<��_b��:5�f    IDAT��*IR
5������~z�S?��5D������$I���\/�?��Nw�f�҅�%Ij�}wq��&��E�۩,�������aFGG��r��H�$I�6ыe���9��=�fZ�[�+O,��#Ԫ�;�$��"5JDJ�r ~�
���s�$I[�wI���>��)��^3d�׏�$I� �	�|�nn;>JOƗ���R���0��ݩ�H�$I��R�������KKK�7��z�g�^��3l��N#IRk�T�Q�:�a#?�©S�!�$ma�%I���{���h�ό@�����xI��5���8��}\w� 1TR��6r��v�bll�����q$I�$I	Yv��j�ƅ��<~r����+IR�ԨR �u��Ϫd>���ź�$i��.I�K�����k��oJ�,9| -IRc�;8�o�����Z�B����N���?uI�$IR*�J��ϳ�����r�8����
�<�����H���~I��/R�D�T�!���*�?U�!�$m%�x%I�X{�E�OP�S�!�N �,IR�e�n?��[����=1n���1<<��Ȉ�vI�$I�U)
\�t���9��|�8���J��O/���Y
>��$��"ej�z��Ꮻ����L�H��%د�$����������Ȑ#�V��$��\;G����GG�d+��ly!v��������d2�@#I�$I�6���\�t���y��r�8[^�\���%}p���"V $I��H�H�H��c�⏬p���9D��f��V���B/G���ߘ�X�$�^z�s���}�q B5u�-������FFFhk�=I�$I��1���������޾v�b�L_�̣'f�>����$�N"�5�{�N�߃����Ku$IR���.IjI��¿�[�9�v2t�+IR}���r�{�sp��ׂn������066FWWW�8�$I��R�T�Zv�|�r�8[ޥ�+<��%�>ub6uI���H�%�ﻉ�@��N���"IR3�m'Ij9=�H�_v�oJ C�����$���q�;�g�H�'�]���6v�����(��H�$I�D�Xdnn���Y��|�8[��u�<��c'/Q-Y�$i�U����%�ᗻ)��K<�^�A�$5w������;vV�������2d���"I�f
n9���wO��-��N!v��������d2^Y.I�$IjN���\�t���y��r�8[��z�g�^�3��R��$i���(��{�Sj_���$IR3��.Ij	�{W~�]�9�62�p��$i�t��9r�n>:J&[���VOO������-3�$I���#�������,,,P��RGڒ��*�]�чfX�+�I�6O�"�R��T��
?	���O����c�$msww�P��u^�d��I�ZF_�7�� �n�I-�������ddd���1���RǑ$I�$�U*������˩�lI1F�/\�ч��~n�v7I�6C�J�<P�h���UN>S�A�$�bO��m�q��\_�I�,9���c$Ij#�}�y�~��A���W+��088�����H�$I�T7�|���9fgg)���lI�+<��%�<y��I��U$���{T��UN�<��6��m��$i�������g@{}ge�ҍK�$I��8z�n�ۨV���w����att�������'�$I�$IM$�ȕ+W���eaa��~j궳|e��O/��C�TJ��H���Ej���Q���*mߟ��ɺ�$��l�I���^���p�޳�r.��$]�����s��{h�(S�y���hkkcxx���qzzzRǑ$I�$)�J����<��Ӭ������l���<��,��
H�t-"ej����K���k����$IR��ɓ$m}�x$�[`G}'2t��I�����#{�󞽴uT<Y�*�عs'###��dRG�$I�$�)���2;;��ܜ��]�R�³�,p����R��$i�Ԩ�q�O��N�����6`�$Iue�]����pd8��e�C��d���%IҶ�֖Ꮋ�r��:,�_�\.���(ccctvv��#I�$IҖQ�V����ҥK,//������U�>3�#N�zٛ�$Iz}"5
D*�v��UN}��$I�-��������@��r�˧$IW�3�Λ�9����"d<1�
!044�����H�$I�����y��昝��X,���eT��g8��).ϗ�]�$IW/R�FC��� �j~N�1P����S��Eݛ�e���2��� �'�J�t�r]��������F�L�-tww�������q$I�$I�vb�\�r���Y�ћ�^�Z-r��<���ea���I��N�B�А�=��Y���F�$i3�۔$m9=�yK�����?-�!G����$I�Fz�r��M9tc?�h���hkkcxx���qzzzRǑ$I�$�e�J%��癝�e}}=u�-!����<��43�X=�$�jԨQ ҐoW!��UN��$I�,�2%I[I��؏F�Yh�q�������$i����ś�q���Q�z��k������8��Ä�6]�$I���������a~~�S�_��K�<��4翼�I�^�D
D�.%�~��Vx`�A%I�&�.%I[���P�U�҈y�62�p��$���o�����j9qdK�f����011��;RǑ$I�$I/S�T���gjj�����q�����|d�3O,��W$Iz-"%j2+����k�����$����$5��~8>6b^���LJ����?�[�q���*Ol�Fzzzgdd�l�[b$I�$Ijv1F�\����,���,-��'�ҩ9b�w-�$}c�x�\���~a���F�$��p7)IjZ�ܾc����31���@{c�I����;8ĝ��ch��j��_M&�app���	���SǑ$I�$I�S�T�ҥK���P(R�iz���y�y�|x�Z�j�$I��F�<�Z����w��З5P����.R�Ԕz��@�w�[31C�.�ƌ�$i�:|�(o���}�J��:NS���ftt���q���RǑ$I�$I��Sݯ��r�'N���#��%IzU�"{���?�p�_7j�$I���GIR�	}��?t6d Y2t�(I��w��������j;=d�	!044�����H�$I��:+����2==M�\N�����y��K|����I���DJ�(6r��g(��2�_n�PI�^�M>IR�������53�A�\%Ize����{��k����^E.�c||���1���SǑ$I�$Icd~~������S�ij�+y�~t��N\"�,�K��J"Uj䁆��y�w�r��F�$����$5���#�o��Ȑ#�֘q�$m1����-�`�P�b��B`�Ν���144Dn�%I�$Illlp��%fff�T*��4�+Kk<��%�zxѢ�$I��F�<��ݬ[	��Y��?���$���]��ؽm}���H�I�AO/3d�"4j�$I[ȋ����6j5�]����������#uI�$I�Ԥ��*���LOO����:NӺ���ӏ����9��$}�H���~4��*ߛ�ѩF�$�,�K���ɑ�U2���Q3md��(I��4�w����:��2T���q�ROO��㌎�����U�$I�$�v���LMM1??�my_��u�yl�/����I�^*R�F��# ��UN�I#�J��"�}��$z8���)`�Q3d�l�8I������o���
B111A�8�$I�$i�+�J���0==M�\N�)]^\�K�/��cK�4H���H��a�E��J�� �5T�$��.Ij���z(�� ?�ȩr�9R���6�wo�� �cT*�L}���v��Ƙ������$I�$I��1������+++��4�ˋ�<q�O?�h�]��D�/��k��D$|�'��ȡ����.P��0�?�%�p}�2t�6n�$IMld���~�u�����
zzzgtt�Lƫ�%I�$IR����255���<16�D�-���:O><�ӏ.-�K�Dj�T9t��[���6r�$�u���$5D�?��t5jf C�n\�$I���>��N��$����ccc��#I�$I�ZT�Tbff���i�e�߼܋E���<�@���"5�D�7�l�O\��r�K�Z��?IR]�⮾
�OE�w4rn��9\�$I�nh����C����q�J{{;cccLLL��ٙ:�$I�$I 1F��昜�d}}=u���pi�G����W�=�$��EJ�(6z�kd�c��4z�$�u�ۓ$�M?G����p��sd��eN���z����]o`�z(�K��4������%��/I�$I�Լ������faa�c�8Mev�
'�d�B�	I�Z[�*��+�O+��׍*Ij��$I��8��~�h��9�)IRS�̵�w���vQ�y���B111A�8�$I�$IW�P(0==���,�J%u��c���ENa��K%�@H�ZW�y"�F��,���#W=X������$m���W����ȹ�� Oa�$����w�� ��9B-ZlQ[[���LLL��ٙ:�$I�$I�5�V����155���F�8M�V�\xv�����ʢ��$I�*R�@���=�߹��/6z�$i���.I�4}�yg������NΒ���&IjA!�����R˧��4r��W���l6uI�$I��Mw��e���Y\\L�iT��s_���g.��SǑ$)�E"�F�-��N��EX�t�lJ�6C��؏F�y����i#C�4IR+��	�����P F�����{�nFFF��$I�$I��������$���>#zA�T��gy�3��
�?�$��H�����@�����R�ᒤ�÷���k�˱!�ׁ�6zv����I�Z�u7�qϻ��Y������`pp0uI�$I��$
�333LOOS�VS�i
��"g�\����Tʩ�H��h�h��.2[��:X�����$�n=y{ ��ݍ���Ih�a�$%�{� �|�!��2��B�o�>���SǑ$I�$Ij
�j���Y&'')����t�V<���>t�X�&!Ij�56ht���Ϭp��F�$m}��$I�G���O�O��&C�@[c�J����H/������\���l6���(����#uI�$I���cdnn��/����:NS������x��KH�ZG�F�H%��?�P��e��`�$is�&I�*��i����ѳ2t��%Ij�=��]�3q��r�Ӷr��w�fll�l����I�$I�$ma���LNN����:JSX�[����pf�;I�ZC�F�H�R�p!]�ԃ.IڲܩI�^�~��~8���Y�t��%Ij;zr��7q�=���q����a��݌���H�$I�$�^kkkLNN2??O�1u��.M�p�����$�5DJ�Hr�R1���p�_�.I�zlH�^�^���_ :=;�A��F��$����2��]7r�!
�־6:���]����``` uI�$I��m�T*133����J%u��b����~�"�˵�q$I��H����E��]~x�'�>\���Xp�$��an�)��ˑ�)�g�$4�S/IR��~lw߷�j��O��d2����g����RǑ$I�$I��*��W��R)u��*�*_yj����T�t{I���� &(��D·�q�K)�K�����c7��%��]�R��$�a�ﻞ��RK_��fe߾}tt�q�$I�$IR#�������} ��Z�'���s�Z&uI��F�<�$7��!��*'%�pIR��.IzE}��H�%`G�g2d��F��$�av��M﹞�=-}t{{;�޽��6?l�$I�$IJ)�����=�kkk��$uei���8ͳO^�j�$i���(I��*��*�?��v����.L��2�u���s~4��@�@7�%J��Mu��yǷ����(�
��$�b�}Ϟ=d�~�&I�$I��l�x�"+++��$5;u�?s���b�(�$�M�@�r�ٜΒ��2'�&	 IjJ�%I_��#��d��4	�Ȓ��I��� w�sG�:A���:N2�\�ݻw3>>N&�ϒ$I�$I�nyy���ISGI�V����<'>3��j-uI��"R�F��V"���8���H���BI ��V�W��)��ɐK1Z�������|�{S�yb���$����޽{!���$I�$I[���/^d~~>u�d��*�<~�����RJ�F����ɓ�mV~n��UIA��,lHR��H��s?�?	$9F5�A���%I��������7��W�Z����DOO�w��.I�$I��Mlllp�����[�0���"����K��!��K���D���C��;�5�w�sb6Q IRp�%I-��cC�}�w�I��Жf�$Iu�?��w~�fF�tP*%��1���~������`�(�$I�$I��B����$����j��q�X�_���S\8���I��R�JH��OA�#�<�@� ����aIR������>p M�@�.�4�%I����6��]7r��(7R�Ibpp��{���ח:�$I�$I��T*133���d��b83���K��Q$I�D�"�T*�?^��Ϧ
 IJǂ�$��>�<	�J� C�. �f�$I�,���7����X^O��B�ڵ�}����ۛ:�$I�$I�(��LOO355E����L�y��y���6b�8�$m�H�"�r��v��4�Z�t)IjQ�%��ܛ�e��O�JȒ�� I�vq��0���mEbl�W!FGGٷo�\.uI�$I�$5�j����SSS����p�e�|d��_�&�|&I��/�'������eN=�2�$�q�MIR���νmT�2�	�\|$I�B��������ގ�{Qg�]�$I�$I�ȋE���ɖ<�}ia��>{�ɳkX͐$m�25
)#�@��UN�A����p%I-�������J�!�A�\z$I[]6��w��-ǆ(��4T���!8@WWW�8�$I�$I���*���\�x���1F&�_恿���Rk��%I�S��B�=٭���UN�PKB�T�%i{����?2�Bd�$Бj�$I���ws�{��7�1ك����.I�$I��k��E�r��3�_��禨��iH���*U�$,��:�g����$Ց;'IڦvqW_�ʯߖ.E C�@[��$m���~���7�?(�˩�4̋�������ݝ:�$I�$I���V.�/_���&9��2�5$I[[텒{�C�#\Ȑ��N�HB�T7�$i����3��N�"���@6]I��QGg�����K�XH�a,�K�$I�$��Z��>u�2_��\�o��4$I�O$R#TS����p�7S��$m>��p����+��T9�풤-���w�X^O�a,�K�$I�$��Z��^�F�=����"�B��o%I�6ϗ�cڒ;>�J�8��c��MXp���#�q����OH����r{7�%F��E���=�v+�%�����b�$I�$I�Rkբ��Z��O��ĩyb���$ik�Q ��[��mY��K��H����#I�vqW_��oB�`��,�py�$mE;zr��C�1q��B��:NCXl�$I�$IR�iբ���e��榊��H����()��1�|x�'R�$]�����r��ܘ2G�69\Z$I[Mp�����޾���J�8B`׮]�߿�����q$I�$I���ъE�#�]��O?��jk�.)I�^j��$?H� �[����"Iz�l!J����@�-�/e�@;:qY�$m5��?td��S�i���A<��$I�$I���2/^dzz�Z��:NCe�zt���OS���M���D*D��>�J�8UN�D�t��	I��z9��d���r�$I[G_���F�bk\����ρ���OE�$I�$I�j�r���I&''[氊��u����~n=uI��J�J�<$����FJY㱹�A$IWɂ�$m1C���H�7��Β!G�=uI�^�w�s��o�Tʧ��===<x�����Q$I�$I��k���y�瘟�o��{��g����ϱ��'�K���H텓�Ӯ_.j^��I�H���wI�Bzy��P�C঴I�����1$I�
{�-����x��������NE�$I�$I�t_-�����"�>4��H|��$g�V6    IDATIW!Re�܁B ��
'#uI�kc�]���>��/�o�i�2tȦ�!I�k����}ｅC7�R,Rǩ���N������!��$I�$I���������r�J�(1;�������Q$Iz�"U�@5u |j���UI�D���l;HR�=�'��I���O��$mo<~���s?��z�(u���Ξ={ؽ{7��k�$I�$I�Z��˗9w�kkk���]�R���f9��i*ek��� R� ��G��,��-����Y$I_�;Ijb�ܾc��_��Rg�Y���CI�V�s���00��\.��SW�l���	���G6�+�$I�$Ijm���?�|>�:Jݭ,�9���{f�����Q$����D��8�T� ��W�G��Tw�i�����Y K���%I�.����w��-�)���ccc�߿�����q$I�$I���cdaa�s��Q(Rǩ������ϳ�RKE��o(R��%�U�߽��?ND���,�KR��η@�?����Ȑ�%C�����=����Sǩ����8p�\.�:�$I�$I�Դb����r���m�c�X�ӳ���D��$5�H���1 ��?Z��Ϧ"I��l+JR����'�_��h'C'.��fֽ��w�m���Tj�au�b����+uI�$I�$i˨V�LOOs����j�8u������9�/l��"Iҫ�Q"6Gɝ��? l�+�%i��(IM�#�^���㩓���vO��$5�7?��޵�bi=u�����������"I�$I�$mY�r��{����m}d�y����)j��H��uE*�h�Nyx�F��:'fS'�$Yp�����mU:~7�;Sgt�pr�$I�id���}�v:�J��ĥ��n������p�(�$I�$IҶ���9�<������Z�����G�"IjV�
�<M���T �m+�8�:�$�:w0��Xw�!��#���Y�r�$��e��{�-�p� ����b����}��111An�$I�$I��zX]]��ٳ,//��RWS.���_��b9uI�^��'��9j�@��N�V� ���lJHRB}}w$��3u��:Rǐ$��a�w더k����l6˞={سg�l6uI�$I�$�%���q��y
�B�(uS)Wy�Y���L�8�$��*U�4I�=?�ʩ� j��HR+��.I��r� �"Ж:@����1$I��m��C���nJ�b�8uB`hh�����RǑ$I�$I�ZN����YΟ?O��}O:�����?}���R�(�$}�H���9J� �����Z����A$��Xp���������	|_�$�/�ۛ�g/I��pۑ}�������3���:Ď;RG�$I�$I�Z^�R��ŋLNNnۛ$+�*O?6ˉ�NS�X�$5��'�7���V�| ω���HR+q�"I��ݻ"���M��y�]���H��7t���}����̶=-�����288�:�$I�$I���)��;w�����Q����:_����\ȧ�"I��Djl���>Z��C��HR���.I����"�O�Rgy��vIRsz����Jk���EGG���gll�ܒI�$I�$I�luu��gϲ���:J]�j�����LQ)�N#I�KEj�TSyQ1`�ӿ�:�$�[��� ;8r_ �i`O�, �@�n�풤�ҿ�����8|�J�B�8�.�Ͳg�n��f���,�K�$I�$I[@gg'ccc������F�RIiS���Ѝ���Y^*�Y�������K�·���L&uI��ܕHR��r����Sgy^�,]@&uI����݇x�;�����:ʦ!0<<̡C����HG�$I�$I��cdvv����S.�S��t1F�>�����J��:�$I/��(i��7~w����Sg���ʂ�$��G������S'�k�Nn�׿$�9����＃��"�j�\/�i8|�0��ݩ�H�$I�$I�$�J�.055E�ۯ�����g/r��e��H��E�BS�܁/�h��u��:�$mG�D$�����@���@�@��vIRS!��n��ݣl��S��t]]]:t�����Q$I�$I�$�I>�������ϧ�R�/��z���Z�(�$ь'��"��q��A$i���(I���7����G����ײd��_���f0:��|��d;�ߩ��l�={��o�>Bpݕ$I�$I�Z��+W8s���l���"��0�3�.�FIR3x��^J�V!~�*��$uI�N��H�v��;���"����(Xn�$5�l6�;?po���Tj���ޑ�n��V-�K�$I�$I-$��1>>N{{;+++���g{G��bl�.M�R,x��$)�@�@�i����LK�ܟ:�$m�%i��p������@���vIR�{`����]�֨T����k�����7���ݻ�f�bI�$I�$I�(�@__����j5���RG�T��9��eB���u|�(IJ)�m��{��NvO��S��0I�F�8$i�r�' �/4����X�j�@�����f�ｷp�wR(�S��T:t�����Q$I�$I�$5���5�}�Y���SG�t3�W�ܟ�g�r%uIR��Q"RL�e���;�5uI���=J�5�����_��wR'y�@;r�cH�Z���]|��H������!0>>���=�]�$I�$IҫZ\\��g��P(������2�>4�c������$�)Qk��;����/s�B� ��UYp���i�[z
�~xo�,/e�]��Z�{�}��9D>��:Φ�����r���$I�$I�^�Z��ŋ�x�"�Z-u�Mu��"�����X�^�.I��)S��>&�����9u:uIڊ,�K����w���'�H��2���_T�F��[�{��]�V/j���9|�0��H�$I�$Iڢ��"�Νcnn.u�M��^��=Ǚ/-�{JIR*MZr_���UN�I� ��ո��������g�ؓ:�K=_n�4YIR:w�����ȯ���i���ؿ?���I�$I�$Iҵ[^^�̙3�������.�[���<���s��$ik�T^(���Q^�����1uI�J��H�V���w��Sgy�@;�풤D�v�O���C��J��q6E���n��Vv��i�]�$I�$IҦ��r���������ʶ�����7�du%��R�\�$5Z C C��:�Ke�L�*1�g4Y�^����	Iz�z9�C~hK��d�LC�Ԣ��}�7߷�Ba��4����u�]ǎ;RG�$I�$I���U*Ο?���1n��[���_^��?�@��=�M��������c���Vi�x��IRS��.I�X���'#񓩃���vIR*;zr|�cG��r��:Φhkk���������"I�$I�$�Ŭ��q��VVVRG�4��y����L>�}H�$m%ϗܛ�S�#����\� ���,�Kҫ�7���G�h�$/g�]���mG���f��}^����p��a���SG�$I�$I���.]��ٳg���"�Z���gy�/'�V��H�+R}�$�����޷ʩ�S��f��A����9���G�L���,�K�R�����q����R)u�M����u�]G___�(�$I�$I�@�R�ܹs��̤��i./���O���d!uIR�y�侑:�+Y�d>�ƉϤ"I�Ȃ�$��^����@�(_#�I���1$I-�7���o��Bi5u�M��f9p� ��H�$I�$IR�Y^^�+_�
MYʻj�Z��Gfx�&��L�8����%�b$~|���!uIj6��$���q�.�����Y^�r�$���;�x�G�p�m#�M���r뭷200`�]�$I�$IR���r���������
1�ԑ�I���^��c��*��j�H���h#RI�����s�E��*uIj&�%�%z9���������vIR�z�(��;����T��a�U�����of�޽�����#I�$I�$I�P���>FGG)
���ԑ�YwO'��<T�4�x�$��2d����{;��Ub�π��E�$mw	��^�}�?��k�e�$Xn�$5H�{�s3�$�����g2���˾}�<�]�$I�$IҖv��Μ9����vp��"��������I��F���G��t|7<���h��kd�C� �q������A^��vIR#����#��ds�խ=��� �&�˥�"I�$I�$I��V�q��E.^�H�VK�m�y�/�s����H��J�<�Yr@��*�R'����Hjq�t���� ߝ:�+	t���.Ij�#o:�=�9���j�(׬���Ç344�:�$I�$I�$�E>��̙3\�|9u�kc�+O�q��/P�Xe�$5B3��y���2�.�"I��+�Բ����@��A|O�,�$�A���1$I-����|�c��)�J��\����<x�l6�:�$I�$I�$����"gΜ�X,��r��V�ܟ�e�R9uIR�T��ٻ��:�;���sv틵z�-[�dI���fB$@�lBH� Mߤ{��V���g�[�����w�Lwfnҷ;�I���x�����l�F^d[�%oڥ�����o�e��s��U�JU*�T����>Y���327F���C �� 
R�V68�F#-��r*\n ̔��t�=]Je'亞|��UTThѢE***��       3*��h߾}������z3�>z�O[����� �#����7r����l� �Lc����hy��<k�y�[N�q; `&c���v-]Y�xܳo؜�߯��竱�Q��+      ��5>>��;wj||�v�y��;�76�Wt<k; ��<>rO�?���l� �L�� ��T�嫍���`��T� fBYyD���j���)�J��9/������Tee%�v       /���^�@@���9}ͽ��H�Thxh\�C)q� p�92��U�vʩ�$�.��&��Wm� �La��`�h��F�iIe�[N�((G!� �<�q�\���Kiw"�?��Z�d�������k       |����2���jbbB�x�vҔC5�֨�¯{G二� Ɖ��ϫ#w#imP�UI�?/)w?��s�+ �T+��?H��n9G!.� .�@Я��Z��y%��}����A.d�       ��ȑ#���Q*���r^��k��h�Xn�}  ��UFY�����ØJ�^��o��9`� �j志���;N��� ��qn�n��2���9}�=�h��Ū����       9%�L���GG���r^����}s�vl���� �)Wie�wG�z9 ��A�=j; .� �)Պ�$���v��0n \H�]y�-[]�Xl�vΔc4g�555�~�      ����ݻ�H$l���ޞ���>ţ� r^ZO���{��7������ �� yji�L�G]���v���(l; ���ʋt�}+*N)���Ι���2�������v
       �L&�������N9/c�1���>ؓ�^  ޖ��{����v L7��  �n5ZZ�(���[l���v ����1Gw=�\��\׳o����8jjjRKK�����       ��㨺�ZS*���4%�P@�̒�˨����� �nF���\�m��N�+�P��)>b; ����b]Zg��d��[N������?� ����7��cU�b���)�����ŋ
�l�       @^s]WԾ}�r�`�$�?�מݫ�x��=  ���%���3���i��! 0]XW���)#�fI-�[N��� ���,������qe2�9S�p�B����N      ���F�s�N����N���^�G}{==@ �(W)e��q&	W��q���� �>� 0J��ÕyY��-�s�r{�v  -l�ӝ�/WF�9{a���^*++��       '���N�@@���9�^s0Psk�|���z���G �t2��ȑ������������j; �w 9�D_m� ��v���䨈�P  ���k��TW\7W�Ą�)	�jmm�ܹs�8��       (X�������V�hT񸧯Ԟ�1F���U;;�C��J'm �ɉ���+�>Qۑ�Ma�6	��j; �w 9�T+��II%�[N��'�"2�� Ө�4���\5s%���}MM�:;;UR���       Pp�~����522�����*"Z��J�c��] @2���SB<;r7�ֆ�P�T��c `���YeZ�}�<&)h��t���y� `:-X\��X��;��,���i޼y\m       �*--Umm�&&&r�{0�Wsk�|���z��g� ����%��!�nN�e��/k� &��;��T�?�����?ǌ�� �ie��7��T�k�b�q�9S��v       ��~������i����a�S��  ��,yy䮮�R˓jyR��#M �V� rN�V�{Ik��L� �[�(�;x�"e)e2�~����/^�Y�f�N       LA<�Ν;5<<l;eJ�Fcڲy�����5z �we�+���Ր��=�7�l� �����c 8S���I��b;��N���v �4iZT�{\%יȹ�8҉��*--��       ��\��
��u�dR�?8�� �ia�QV���SΤ)��7Cj|2���� 8�Z�#���j��%�#�%g��v �t���%�hM�b��{����       ���񸺻�522b;eJz�����S<��z xTV1�J��8��i����C�C �lX`�K��
?&��%gf�("��1  � R�?�D��i�Ӟ#�kjjj�h�"�)       ����_===�d2�S&mdxB�=�GG%m�  �+�UT�<�3q��{ݨ�� g����թ�xB�?�:�-gf�SDb� �M�5���N���S&���       PXb�����5:�{�i��}��A}��I�� @�s�QTR�v���J�M��Ol� ��0p�Y��"#g�d��n9#�("#�� @X}�]��Q�c�S&���       P�\���Çs����]���s��N0� �/WYE�z�>d�~gT[�d; N�W� <�X��9Jo���v˙9
3n ��@���޽Rus�J&s�q�~�_�-Rmm��       �E�x\�����2i�����=>��� �q���*���>�Ȭ�{/����� ��*�%�̫��l��͉q;Wj 秢�X?���J�9w٦��Z���*++��       �������N>�/�F�E�!-\R���	��! ��9��UF�k;�L��tgH�?I���v �k�x�G���o�<�{�yIM�{Άq; `:,no�]�/W<5j;eR�����,��_+        'cT^^������(�J�N:g��OZ���3�?0.��N �/F�2�_�]a�ޗP�G�c �,Q x��f��Ėo�q��߲�<6>����lg�������3  9�o�����i":f;eRJKK��ե��*�)        �
�����˝���1j�S��ڠ�Q6��
 �#�#wG�wC�}(��l� ��WMxī��TU;����?��ݣ�~�Q�<��F��s��((G!� ��u�.UyM6�.�c4g�555�~�        ����!uww+�L�N����	��q��x~� �0We��q.\#�ߍj�� \p`��_�~d΂�w|�?��U���^�;��-�X���Q�W��(l� �۪f���Z�pL�L�}	��Z�t�����       &%����^�DB�s�Y8Ts�,MLD5x,.�H ��ȑ�/.���Tc6���m� (l�X����~骥�������u�n��F]��[**.Ҿ�{��'f*S�d䗣Ȍ�5 ���c�n��S�T�<�U�jkk��ѡH���       ��qG�f�RQQ������fm'�����EU
�;,ɱ� �A'F�N.��e�kBj�$���� �����槿z����;W�wS��(�H���^�3��A��δ�}Չq{X��	 �
c���Ю�+���l眳@ ���UWW�N       �x<���n����N��C����ţ�K  �*��\%mg�#��Q��7�\�- 
KM V��W�����\����ch�νz�7��������x�'��.��. ����P�    IDAT����.M*����9g���Z�d�����       @r]W}}}������nndxB/oܥ�~�_� xS.��%�gc��cI��� y��;��_~��/�q�7��?���U��^w��q>���% `��+u�.R2=f;�9��h��ٶS        `llL��݊Fs�,z*��[/�֮OF�g� ���*.W)��ĕ~=��J���. 3�W� f��=��W�t�m����>m��z���������#GI��� 
B��yZ����'l��������)��N       �l6�������N9g������W���l�  rPV1�ʍ͸���/���| 9��;�����ŧ��|�-3��L&�zcJWݍEd� ��1�躛;���L�x�v�91�hΜ9jjj�1��        �chhH���J&��S���C�ze�M�M�� �ĕ�**W�)�j�J�^͍��4�+ f��?���Wݴ�����k�cϜ����dTĸ 0i�HP��r�BQe2��&D8֒%KT^^n;        �R)�ܹS�S���HL/oة��� L���%���|ٕ�W�V�1�- �w ���O������\a��g��~�r��R  WU�*��\�TvlO����^������R       �[����g�e�Y�)�$���vk��Q1� L�����Iʍ�y�y=�؍���� ��W� .�u�?=���.^{�%�[N���^m������3>>$Galg r̢��xW�&�#�SΉ����ŋU[[k;       �ӊF�ڱc�&&&l���u��;�zo�9�s  9%�LN�ܵ%������� ���;��q��%6~���5˗�n9�DRo>���?�I￾5g.� ��ź����Ɨ�KJJ��֦H$b;       ���f����Q__��s�k�a��y�2i��
 ����#���-���;�z{�v������{�u}�g?���e�[��������z���5||�v ���1��miA[����s��РE��~        ��Ǐk�ΝJ�ӶS�������nM���H ����*f;cܷ
|��;��Ʋ��ڴkWht_b[�ʥ�l���T2�7�}C���Uw ����}���
ŕ�z�q>�O---�����       ��%	�رC������ꥍ;5П�| �7�J*����x�(xݨ�8h;@�`�`ڼ�wo�XO�����m�L��=���7jӯ���1��@!��U���X��XN|����Tmmm
�öS        8o�몷�W���9�>}*�іv�g����  �U���]i���1�3`�@~��3�i����ű��ۚ��n��Rɴ�}�]m���zm���f�� 0}�[t�]m����e���F577�^�       ���А>��3�R)�)g庮>x{��㈌|�s  9"��\y������+}kL��� ��tp�ֿ�W�ID��5ϱ�2�����{QO���t��Q�9 �l���Z}�l��Q�)g��ڪ��J�)        \0�dR�����rNv�8�-��)�f� 87Y��*m;c2>r��ָ>8f;@nc��<���⒢��EK7�n�%��j�h�#�� y���-SӒHN\����Pkk�����        fġC����#�um��Ց����.E�l�  r����=c;d2vd�k�z��v�������l�{E�����m�x�������z��ґ�\u�\
t��)X�P6��/0c4o�<͛7O��2       PX��ƴc���q�)g5:�Kvj�pN]� X�*��$of�۳r��л�m� �M,_ L�/^y%\���ն|��-^������q�2��% @RլR��+�q'l��U8V[[�JKKm�        `M*��Ν;500`;�R���<�S=;��| pvYeS��ܻ3�5\r0�B0i�v�
��&w�-o�g�%|q���zZ��� 8ͭ�Ν��ż�|���j-Y�D~��v
        ���߯ݻw�u]�)g亮>��~����l�  <�UF����O�����Y�%w �����lڵ+4ޛ�n]�>�vK��f�ں��� �uk�.Ѫ���z�r��8jnnVCC��        <g||\;v�P,��rV�v֖�z��8�S  �*������+>�ʹ��;��`���}~������M�[r���=�/���_<�ý�v ����eZ�Y�x<n;�B�����UZZj;        ��d2ڹs��;f;���ŧw+c� 83WIe���1YK�vL�� 7��9a�~ap� ���st�/SU��T*e;猪�����*��o;       ��p��!����u]�)g4x|L/>�K��Y�)  �s�PVI�����9c����Ӡۯ��V�/�ݒ����r� fZ(�}u�����Y�al�Ѽy�4o�<��x        &cddD;v�P2��1`t"���LGy�  ���br���1YI�k��΀� ��2�=��A��;ZW,]h��Pd3Y���;Z�����?q� .���b��W��H�x�jK Pkk�*++m�        ��R��v�ء��a�)g�Je��s;��{\L{  ��*��$�r;#}���MF� ΄W� N��O?f����+�6�n)T_\u�����o; ���yպ�)��rF%%%jooW8��       @�s]W���ڿ��3�f]���G������ x�+W��������m� �&� N����x姝�.k��)��j����ڲ��S9�x! ��9�n]�&���SΨ��A�-�1�l       `:���[鴷?{���!���C��� pj����ܽ���Sa��LX� ���]ח~ᓏ;Vu��n��Գ�٬��\��}\u��Z��E���W,��rZ>�O---�����       @ފ�bھ}�&&&l��ўώ�g�)���N x�����)G�[}J~sD��n�-�|���Kn����K��l��̸� �w��j[Q�d2i;崊����ޮ��"�)        �l6�ݻw���öSΨ���^|f��1�> �Ss�RVq�S`�R���zs�v	 ��U/��w]_���?츸��v&g�ؐ���s�����g; <�q�n��U�K�L�v�i���j�������       �L:r�v�ڥl6k;���酧wilȻ�  ��Jȕw����VX����q�% ���; I'��ze�ۭ���݂�s]W￾U���y���kJ��� ��P8�{Z-_8&����،1jjj�ܹsm�        P���ǵ}�v��޽~;1��K�?��C)�)  ��*.W��s��}qTe7K�z�1����\�u�x��햮%�l�`���镧_�����}��v XQ^Y�{�X�w��
���֦��2�)        �L&��>�L�SN+���g?S�Ψ��  �ʕ�UT�w�n~:��y\#�H���	8��  v��ky�+����݂�
����{�V��~�������I�ދW ����t׏�+����rZ������TQQ��         �q�������Q�9���9Z��F�dL��� ��H2�K9y�]�B
/Mj�Ҿ�� �0p
ܢKn��qq�7mw�U_�57��mު��F�����a�Y p��u��Mw�)���}޼yjii���Kr        �����
���ippP٬��u��i��?�ա��2rl' <����'Wi�)S�R�=�+� mwm� ��5P��y���/[����;0s����W�o9y�}�N���/�\٢�ߙ�ht�v�)9��%K�h���2��*        xU$QMM�����Jy�
�1F���UZ�Soϰ�2r �k��L����C��T�3����;P�~��7�q�U��k��|����G4tl�v ����/��+j�z�r{(Rgg����l�        �s���UWW�X,�h4j;甪kK5�>�}{��f8� �3sr"���//
�qNR��m� �y܁��߿�w��]��x�W�o�W��뿻L�����m��Ryy�:;;UTTd;        L��8�����8��sJ�E��S��=�ʤ� ��ȯGг�S�bEP�I�?g;��b���앿]�����1�B�������S��9�Uw �g��m�^���CJ&��sN���Ammm����S        �������Tr]�v�ה�E4��T�=�Jy�# �%'F����#]RciR���n0s���}������7���qf�П����z�2��9�Uw ���9���5��s�N�m�|�1F---�?��r        �/�h֬YV*����5E�!�]X�����ٮ x��_���ő��5A�N'շ�v����(��?<��˿}��S�c���骛�<y��衣<�Uw �C~���+,�+��ޣԂ��:;;U]]m;        L�@ ���:E�Q�b�[��#A-h�V��!Eǽ�
 �##��#��c�o��0�P��l� ���৿��5�_��`(��XL�W�o���j��kd$��իt*7_��mE�!��'�K��'ZRR���.�N        ��8��������5��_M��u���GxR7 �#G����K���%տ�v	���;����c�߲�U�	�Î��Y��Zs����mj�ߠc}�4xt�v�Q^Y���F���S����ҥK��        �1F����D"��Q��-�448����$n� $ɑ�������tcP�I�j;�����c��-k;/[������qAC��]u��}��� .���r���J%R��c�`�577��        �P���JCCCJ���Y���iq���G5x4)F�  I2�Ir%em�L�cdn	k��	�����U+�����^���Ү7˫���[PX&Ƣz�/��_<�]����=�J�ߥxr�v���������v
        �$�Jiǎ���5���Wvj��� x ��������%)�*{ø>x�v���Ug ���j_tђ��j*�[PxN^u��f���6���[�xr�v�����K����S        �E>�O���r]W����s����M���:���; @F��_RZ'��9'`dn��ᅄ��m� �^\p��#�>i��T�mV}M�v���xT/>�y������ &�s�<]���J$b�S����F---����(        ����~�޽[�������H.� HRFYEss�~�qW٫���v�! �w ������ʻ��ԗ�nN��ÝZ���z�����q�^�X���S"���5s��USS���%5        ����m߾]�T�v����>��6�W6� ��*���wtn9�]9�w��0=X� yb���+})�g�����[�s�H$��soi�#��k����AkoX��U��ǽ5n7�hɒ%�����        <.�k۶m�F�w��w�1���^eR�� �d������'#]����C �?�@x�c�c�ݳ�ai����{�6�v��?�A�Cc�s x�Mw���%%	�)_��ޮ��r�)         G��im߾]��öS������r�R	F�  WY��*m;�|l3
^=�?�p~x����s�@����[̶�LUŬ
�Z�R����Z�Ѭ��q���˔@�������8�d�[��D"���RII��        �C�Qmm�R�����m�|IiYD��J��3���>� �8##��w�v�T�J����mT����0�@s]׼��'�.Y��f��~�OZ�t�����QQqD�w�W"��M�ct�}���ɯT*e;�K*++��٩P(d;        � c�������=wɽ�$��y%ڷ���)c; `��sr䞳��,���3�c Lw �-Y}�sw]a��*�O\u��u��`���X�1�Y .����5��(���/����jkk���Kg        p~���T\\�����w����8�T�=Jq 
�����#�!�;�����v���p�X� 9�э[��u�;���kq�b�tߍ���o(RQ�^%b	�i ������UԺ�d������竹�Y�p�        L���"UWWkpp�S���4gA�z�W��c��92�\y�����5T�P�F�! &��;����?��+�\���`��W�k�ڕ���;�ܱP�����=l;�yp��X��ʴ�٬휓|>�������h;        �`0���Z+�����HQPs����%�k  6�$e?�W�Z�l�P߫�C Lw ���߽�7_u�t�v
`���ӂ�&]�u���kN\u�}���@������jW�<��`0���NUVV�N        y��󩶶V�hT�X�v�I�HP�U���cJDm�  �12�KJK��g�S�6������d;��c�䐟=���V]u�?c���?_u����@��}��5
�&=5n/..ֲe�TTTd;         �qTSS#�u5::j;�P(��+up�q��@3��r��r��uA5t'���� 熁;�#~���W/�t����ہS��U�ۿ�HQ���G>������WVV���S�@�v
        ( �UVV*
ipp�v�I�P@M��u��1�'l�  l122rr}�n��-a5��P�n�1 Ύ+�@����w-\��^yU9�;`����|�M�d��}����@�
�����^.��ֻ����jnn�1�<        �iǎJ��3"�N$�ܓ�4x��[��e�������JQ#�[cz�-�- Ό�q?}Ꝺ-�v�ͩ��nrف=��W���g5||�vP�B��}�R9��픓�1jnnVcc��         IR,Ӷm���l���&���Ou�?#�F P�\e�����uܕ{ո����x�	x؆-�+��陳pn�� _��i���\ufX�(�{�T�y�X�ϧ��vUVV�N        ��d2�m۶i||�v�I�DJ�?�MG��� 
�������C��A��W���C ��6�ڴkW(v8�g�Җٶ[�|up�Am��&m���:�Uw�B).	�{_"�Dm����ѡ��R�)         ���d�c��N9)�Hk���t�7%fG P�\e�jBypRr�Q��Q��;?h�� ��w]_��#-�l]h��geUeZ�v��x�5/]���q����䕲�~���ʸ�SN
��Z�l����m�         ���8���Q2���%w��������I�\�m���)�v�=���� _���[.[��ҕ�� 
���hAk����:}��o*	�P�!Ţq�i@N+�(���r%R��SN*--ղe�
�l�         ��1F��Ւ����5'�|��/��� 
�99=�X�s�2]I]���=�����;�1�y��鼤�&�@�*�<q���ߩ�5]JƓ���+��5,0e�E���/W,1l;���jutt����N        ����
�B!�N�tb�޴h����PΏ S`䓫�����,	i�.���C �w�C~�����ei��d�ƦF]s�Z���免�Rv��؄�4��C��O.W<�q{}}�Z[[�8��        �))))QII�<q���������f� ��ȑO�ҶC��YRc"��7l� 8��;��}����}U�4�Gw^S\Z���:u�C봨s�&F'Կ�_x��HQP���JeFm��4w�\-Z�H��        ����H���P6���#�����j�?��Q�= ��f>�䞲2��aR�� ��<�_^�v�-O���r�������z��ґ�Gm� ��q�1F�-RCC��        �i����'�(��N�$%i=��6=�W| ��*���3�C�ȽyT[7�
cZ���7�X9gɜ�K�Jx����٬�n�@�٠�7nQ&ͣ�P�B�~��˕u�m�H�|>����TUUe��~�    IDAT;        ��H&�ڶm��ǽ��L"���'���A>3���*��\����i���j;(d��~��g�5��jk�l� 8_\u�����Gl� 3&��?^#���S$I�@@K�.UYY��        �*��h�����"I�Œz�m8��� �q�2�����ǌ�5�ں�vP�������q���6ϯ��`zq��$����\!��� �pX����D"�S         f��ڵk�>l;E��&�鉏5�M0 (@eS���w�J]>����
��v P�w]_f��m�͵�`�c��Ԩkn]���Q�*th�!��xc L���}�F&����%%%���R8��        0c�1����$���X����U���c�Oخ �,��ϋc�UF��+U�	Iَ
w���^z�+KWu�����+*)R�e���/oS��.%�I�s@n6/�����;������S$I������T ��        `EEE��~����m�(�k��J��;�D��� � #�N\p��N��S�-M��I�� 3��;0�y��Z�fŭ�; ̬/]u�����}���ꎜ�����S$I���joo��8g�/        䱲�2����S4Q���=�$#w (('F�i���֐���`;($܁��~���i�U��Gc��(d����U��=����7W�����.U��O�jll��ŋ��V        ����TVV������aa0PSs���=�� 
����m��3��jN��m�%@�`�̐_<��m��,�����76 ��|���ϯ������0W��M'�헩�"c;E�4w�\5773n        ��H$���JX?�4wA���>�T�'�@�02r���%��p]H�$������f�c?���uụ�e~�- �-��j����ڲ��Sy�"9��ר�"e�҇$-\�Ps�̱�        �i�hT���ɤ�Nh��?Ut��; ���r�撻bF�7F��O�C�|��������Uջkk�l� �-�G��o6k�/׫o_��0c��y`�J�R�/|c�x�b���[�         ��x\�����׳O�Pl�� WYE����`7rW�j�n�!@>�� ��[܈���h��Xi�@�G�uY�n{h��Vw)O�`�A�c�u�^��z�����1jmmU]]��        �\���USS���A�Rv/�F���=�L{wS&�� 
�����{�d�Ѭ_'t���ǀ<���@\�u��p�GZ6�n�ی1jlj�5�����߬��r������4��X��~e2��㨣�C���V;         r���Smm�����L&���T?�X=;�)�q��  f�����U�v�t�q�_�T�o�A��
 O1p.��Wߵiɲ�ն; �/�������ku�R�ϯ�g���w���Z�Yb�����Sgg�***�v         �2�qT[[���1��vΖ��5�!����r�����$���f�2?�Т���`;�G܁�7�?��Wv�c�@�����[��ש��Q}��5||�v�ĥW-��55J$V;�����TVVf�         8����O���ʋTZ�Ӿ]�b� ����=�C�|`:���^�]�^��/|��m+��Wc�� "i�E-Z���Zs�I{��+��	H��e7i�������B���Rqq��        �|b�Qmm�b���ѨՖ�Y�
������ �I~�J��NW�Ը/���l� ���;0�����-˖<X��bV}��ܰF�=x����{���%u����H����a-[�L�H�j        @>2�h֬YJ&���RSW&�$��;�� 
�����*o7I�	��ͤ��Yn�w`�l��`��9�o��� ����W�o9y�}�N�����4U�ӪD2f����H˖-S(��        �ό1���V&����Ֆ�9�Jgb:r(�� 
��OR�����ni�SI�����4��[:1�^U[Ul� ��W�8��cC���1u�Zw_��)�����Ruuu)Z�         (���rG��v�={^���1?����/  ���*-ɵ�2]"�{cH��N�?j;�u܁������>�����sl� ��|q���q�_V5�Tw��2��v�핕�������        Ph���44d�P�1F����𰆏'%F� �猌��G�y�R2�%U�k���<0p��]k�^���e�� ��/�����:5�o��CG5x���,�{\�t���}�ҥr9	        `Cii�"���5c4oa��>����@~3rd$�ʫ-���s��{�v�����W����w>d� �*:q������ɫ��w�*�ʫo��4"EA}��K���q{UU�:::�        XV\\l}��8���kt��E�\1r��f䗔���N�N�CjK����C�\����G7��ҋ�~��~�����~ۃ'���;������p�����~�b�	��f�R{{����)        �xa���;��h��?���#@���U�v�t�V��g�Σ��;�~��ת[���W�H,20l�K��q�$N&��3�=�������L:�Lw��d9��N����6�16��xc�/"�؄�P�T�PU��[u�3Hؘ����ս���p}�WI�|���EM=�:P�(������{z�IfR|�:\u�~�g���ާD��7�MMM��        ��d2��i�%�X,���=rJ�5~� �̜��WUuS��w��v׆N�r�4|�lѽ�>W��%��v��\g���]Z�=_����o_ԡ�����������5l��ݽޫ��Y�����        ����y=��N���鳺�փZY�e  ����j��>����Vu��� @%��4���~�����=�;�\g�0��sW�?��]u?��q��W��~�r5��*���2���Pn        � �tZ�\N����2$Sq�veu�Y�7)�@u�Jڔ���*r��k���ߗ4]u�}�
�������=�{��9 ����F��o�/��{Ծ�]s'�4j�u,�7�c�����t�`BKK�FFF(�        T�T*�|>���9g��3٤�Z�:����Sr�ju�I��+�Ei����\*w�5�ĝ������: l/]uׇީ+n�B��_��6�w߀.zC��Ţ�mmm��        PaR��r��Ӓ{�>�t��賧e�<@�2���Ur%h�Iuj]S�r�|�����{�u�����x
 ~���&]��7��y��z�5j^�'�]��y�C-��}Z__s����MCCC��        *T*�R]]�Ӓ{SK^�)j��Y�� �ju�A��$7�XtM\�O5}�u`��a��}��ŝ�;���ex  ������k������/i��%�qjVk{�n���Z/�8���ޮ��A��         U�̙3z���U*��������)=}`��; T1_e���*,��z*_}F�>�:��Q�~�ﾰ��'�7�']g�JS�T�����Ϳ{�wh��eM�v��������ڣ��r;��        �G2�tz����&���k�tI����ddd��צ�(A��e�W�-E�:�:�]Qp^�þ�y��c�;:Z]g�J�F�7ګ���zӻߤt6�����Z�u���G��_��ܕۻ��488�l?         ��%�Mz���Vy�4 T�so��%�]G	��ꌼ+��|ZZp�J`������]����F���� �䥫�7q��*�3��߾B�ĺ�]]]���w�         v%�I
��ͩ\�x�x��k�s�Nic�}?  F��W����.ӝP����;\'�#
��Oq����lh��� ���Wݯ{ϛ�Τt��1���+dW�w����}c���M�        �$	���kvv��%�x<�Ξz=���ʛԠ �:y��׆� 6\�T������:����
_|��?�����Q �&�7����a���wN��?�������I�        ���.���q5��u��S����� ��қ:JNSXrc\�5��� �vB�x��?13Th��'�J� !{�U�7��uJq�}�������z'������69�         w�����477�䞯K+_��C�2ԡ �*���$���-��;�j�º�\�����;8�g�./,4��� @��k���k���߬���Z~qY��N���������T*m:���֦��a'�        �^2�T.���쬓�M9���cK���*E�k�uR��!�����i.A��H�|�7x�����~�Y  ?y�U���S*�Աg�s��:�z�{��Y*:���ܬ��c��        ���J���睕�ۻ������5yN2  l22�����?˚��wu�g�'��L=�U�I�W��ёݣow� ���^��~W�_�����ڭ�Қ��MMM��         I�J�LFsssN�w�6iaaAg�7$�;, �6���Q>�o�1CI-D�5�M�I �(���}��|`���?1�� @%x�U��o~�R餎~Ak+n
�.%Sq}�w/W���d�P����v         ��t:�t:�����wc���IS'fuv�� P��"�U�T�Λ7���DQ�O�N�D	5��o��j~<��F]g \���������_��?"߯�o`~R$��������:��R���x�#         ~�S�N�g�q��������gh�4���j�kSe���a˲/�e}��� �+\pG�:8�gK����Y  �O-^u��W/U�n��:MLL(�KI         ��l6�D"��{,U[WN�>uR����jc�ɨ,_e�Ql��7����5�����3��j����8���}��  �Uא��k��߹I�c�Z<����O���7�iX���J��w��yMNNRn        �k��f�Fu����w�3	�5�u��YEC� ��ܟ�n����,�⢮�;��_�8F3	5i絿�7C�#�p� `O$Q�X�����膛߬d:��T�U���]yc���b軳٬&''���?         �v�|^�H�IɽА�����%y�� �dd�_�%w#&�����o�����;jέw?��]#��x�u @H�篺���50ѯ��5}��X[�ܚ�;�?�b1��~&�Ѯ]���B�        �ʗ��%IgΜ	}w[G���0S�} �.�$_R�u[����񢦞twԔ/|��pGO�=�T�Gr�E"��F{��_�Q7��z�y�x�V�V\G�������[{�Y^}w:�֮]���C�        ��Q__�r�����P�c��ۨ�3ZY�%J� PU�]q�Թ�{�1Fz[\mwur�u ,�Q3��ٍ���BsC�u �{�B^_u���ᛴ��T\+�س�����c�_������CߝJ��{�n��         D�PP�T
���y�z�u��	m�S���bΗ�7\�%ad�Ϩ�Sk��<8�Wk�	��;�`WO��, ���xF�zӻ���?�*4t���:�t�u�y��/Q�)���dR�w�V"�9         �V�P�������C��G��]�COM�/EC� ���;�_%�9,j*KcEM�u �Q&�}��9�.�9  �[&�Ѯ+&u�6��~�5��Ȫ\.��7�i׮]J�R��        @mhhh���VVVBݛ�$T�בgfdD� ��QD�
��z���ձY��~�A �(����z���5��g\G T��_uǯ�]���p���.�{�}p�M��ܩRi3Խ�HD����f���        @�0ƨ��IKKKZ[[uw�1+y�>�t�	 �F�'_��Xc�k��|x]S�\gl��vϡұ蓙|&�: ����e=r�����_��/߯Ҧ�WZ5��tӇv�T^��界1ڹs�
�B�{        P�J��8����P����{���\�� U����.�K:���{F�?�:`_��j���K���7r��  *�1?����_}���u��Z�p�=��뽿q�|S|��b���ؘC�        ���y�����������ʈ�u�5���ZY��
 ��("_��|�QlI��mR�'�4]�M~�.
�Z�x������Q�9  �'�Mk����ÿ�]�v��V�����_�7F�H��ͽ��6H�5���jii	}/         j[$Qcc����T*�}���y����&>tB�Ԩ �z��%���~�ev5u�� �|e�����>�'==p� P�~�U��Nh�̅�>�]�|�
-�_����Sggg�{         I�F�jhh�����rh{c�ں�t�)��hh{ vy��+��ؕP�EM=�:4
�:w}��5��"� ��GW��¯�_q͐�w�C�J!I���u'         �J�XL����������'�V�lBuqyf^�: T�sW�7%��w�7����uMO����PU{�/�K��s���, ���W���U���~�U���6]���Ő����Ң��!�sa         p/�H(��kff&Խ�Ƭ|S���/�� �l�|�}�u����[��TQ'V]��B�U��}�n�l�t�  ��W�ߣ�=�Z[]Ӊ�N����u�i��뻵^\	5_cc����(�        `[I&�J�R���uo{WAss�Z\(I�wh P~��R�i��%���Ϩ��գvPpG��}��K�H��\�  ���1��қ�:���ߡ��zM��ҋˊD<���\���-���yMLL��>        ��'��(�iaa!���u�6�gO����� �Z��⾩*�~�չQ����� A�QCT�;:����_�"|s ��rY������~yfF��7Q�tZ]t���hh;        �q��Q=z4ԝ�K���S��u/ �_%�C>>�@����E=�5�A�׋�x���mO��H����  �#_��:��J����M&�ڽ{�b�Xh;        �U__���M---��3�I(���C�2ԫ �*y:w���:�MF2��V�k:���0����kT�{}?������B�Gf e�슾���Sq}-���XL;w�T<m'         �z���5ԝCc��� _�P� ��8_t�j%E>#MPAE���TT����������u  ���[?��g�C��D499�t:�N          (���*
���w͈�v�t��/ ����-�˳J�G�!�׃w�b}���}x�ؿ6Ƹ� ������t���C�g���Ą���B�	         ����&�>}Z�b1��ݽ:��qm�GC�	 ���������.����EM?�:p!(��"��ة�����Ǔq>� �����C�û�044������         6x����F��ΪT*��3���=�COLI>%w �Q��p�:#󖔺>���Ӯ� [� l�!�O����|&�:  [1sbZ��S~9���w�ء�����         6��qMNN*�l��Q�K��RY�\� �ed�)�:F���?+&\���;*�S�|{w[��  l��ZQ�o��6�WB���Ң;v��         C:���Ą�1��ܵ�WC�9�
�r< �.���j���ެ���u
`�"� [q���w���]�  `�������������k||<��         aI&�J$���mgOo��=?��eI��p P�"�6\ǰ�H����xQSO���V�Q1�{fi��9g,�� �����������/�NkrrR�_�        �ze�YIҙ3gB��y�:z��̓/��YW���2R���H7����uM�v�x-(
�"8�gʥ���t�� ��z�I�������ڹs��Q~�        ��c�� �    IDAT�������>�7�uX�Ym' �Oq�H���,���`�u൨��JT��ǎ������:  [�����~A��f(�<���Ą��d(�         ��`xxX�B!�};ZtѾ6�
���  �"�����7��?s�x-���m���?�=��v� ����-����Pvc466��         ������&-,,hcc#��]���k�tI�	e' �O�/��:�uF�<��ǋ�z�u�g���m���˓u���"��	  *��wޡ�Ï��o``@mmm��         �����Ԥ��Y�J%���1��QгϜ��:, �tFI�:Wt�nF�1��ϭk��,���\ ^�!�O����;���q
 �(�x\G�x(�}]]]���m         ���q�ܹS�H8��T:�7�mD��B� ���(�:DX���?+M�]^�al[O>t䶖���9  ؊N��}���UIjnnV___(�         ��.��h||\ƘP�ut5�}m��> �=FQE]���7��s�x5����>�����=�o6  �����-���P����i||\��3�         �KR�������C���U�ɓ�Z~�,�� T2�H-=�tEB�5��� �+QpǶ�+ݙ\�x"��' ��|���k���Pv%�I�ڵK�h�<9         �v�lV�rY����wcԵ�A��~A�E�. Pٌ�$_%�A�`$s}Tm����%�a����'������{ӹt�u  ���<��eW,���b�X(�         �J��ק���Pv�3	]s�|��> �=Fq�ڹ���i�5�?��Hl+{���3�{��  l��=x秴Y\������	�r9�         �J��ب���E��
ml��ԉ�@E3��k�u���&tz���o����;���=z�ξ�4�q ����}}�S���|(�C�2         T:c�533�R�d}_Gw�N��ʢ$с���҃J����&�M���N��: �G�=<zگOfR�{>$ ���>�����jkkSGGG(�         �j��5>>.c��=���o�T<�f} �.Oq�P�6���L�&�� R}�a{;�ԑ��
�9  ؊�9��G	eW]]����B�         T�|>����Pves)]����; T6s��^��SV�#�s �q ���a�h�]�  `+_<��o��67֭�J&�ڵk�"�t         .T&�Q�T����]���-kvzU�� P��"�J�|�Q�2�P�EM=�:j-)8u�?������H4b�P  �+���ZY���'�h׮]J&��w         ծ��^gϞ����]�=�:v�V��$�1 P�"��:D��W��EMϹ����p���d<�z<�� PQ���/kq��=����*��X�         Ԃ�~�N���D<��퓊&׬� �c��(�:F�2F��k��g(Ù�3Gok�hmr� ��8~舎| �]���jlle         P+"��v�ܩX,f}W]}FW�0��(�@%�����q��j�߹��q ��+?8��?p� ��(����}L���w577k``��         �E�Q��y���X��Д����Ok�	 U�H2��:Hh�tyR��_��!�YP{(�#t���h4��X"�� ��|�s�h��s��d�Y�ܹS���-         ��d2�X,���뻺z���Z_�� �a�T�从#����?Yԩ��à��B���w��{ҹt�u  ����������x<���	y_�         �utt������h,�k�6.E֬� �c�t!l�F��u���B��S���>�:  [�03����U���'p=���Ą���=          ~l``@�����4��u�m�i} �#OF1�1��������-���]�����t� �����[��j�MK�����r��          �1c���ǕJ�����5wE$�=� ��SR�������!P;j�3n8�g��w�3��  ����%��=n}Oww�ZZZ��         ��E�QMLL(�X��yF׽uB�ĺ�=  ���#�-#�������z�A����:qK}S��u  ��������Y�S(���k}         �W�N�5::j}O�>���ح�(�@�2����CQ�О��C�6��g���O{o���v @�����=����W���I$����~	         �ϗN�U.����huOK[�fg�uf�$#:5 P�"��:Dخ��뾢������wX��ߔi��4�v @���s�������i||\�oo         ����^
�{��q\�,W��Ry2��·���:M���5��;�:���/��r)�9  ؊'~�f�������A�r9�{          �v����)�LZݓJ't���*k�� �=��R���×�ˊ����n�P��x����c��7]�  `+�.-i�>�҆�K	mmmڱc��          .��y���:u��=������4?�&íR �@FF���� !3��j��郮��:Qp��;�ҝ�f��c|� *�]���Vg���f��1��/         PI��b������ѨÇ���Q�]�j`��MI��(�22�G���M�Xt�Շ��8����3��Ie�1�Y  ؊�|�-�=ouG,����<�/�         ���C���Vw�b]��q�ފ�=  {"J���B}D���x:ЬB�������C�s  ��g��܁���0�httT�dM~S         T���!e�Y�;�:���M�6�� ��Q�u��醜.�m�9P}(�#P^�l����s  �U��~�6��Vw�رC�B��          ��<O����bV�\v尚�=I��=  ;<%T���͟�uɠ��.���}?��r�+�x��+ @E��׾����Vw466�����          v$�I����{�E�3���2�5k;  6y2��0�6��e>.�7�:�Ed����������u  �b��)=�m�;�ɤ������         �]�BA===vw4f���.�ڰ� `���j󊻮������A�����5�}���:  [���n��ڪ��a��         �}===*
Vw캤Wm=qI��=  ���{M����L���@��ہ�~F���|� P���״p�y�;��f��          c���ƔL&��x���2�5k;  ��ej����H��&j�����g�5==uK}��GS ���I{��Vwttt�����          �F������٫^�7dtɾN�ڰ� `�Q�u'|颼�����|��|���_l�i��  l���z��Ϫ�f��A.�������          ��d2��c��>5uD$�V�  �g�Q�u'|�_��r�9P�(��=��7���[�1��  �%���%-ο`m~4��ؘ�;         �^mmmjmm�6�󌮹qL��Z� ��(�:�+Q_���/�:*w\����|&�I�� �VL=��|����A%�5�M
         P3�N۫�44�t����am �#O�b�c�2�������E��'�~����j�9  �
���З?��⚵jii�6         ���D466&ϳWú��AշH�om ���$�:�#���7�N��D�[����$��u  �j��_������i���[�         `��d2���6?1z�['�{+�v  l12���'��J�R����Ppǖ�䭙\�?p  ev��N<�k�#����ǭ^f          �=uvv���������&���׆�  ;<�T�u�ᜊ��uT�����������m�m׹� �V��ﴹ�nm�����鴵�          ����%�Ik�/�rHuM��[� ���S�u�~?�=W���B����~]4����  l�_��ξx�����f���Y�         `��F��1���H���7��l�Z� ��(*)�:�+���J�R���rPp�k6���f���9  ؊3����߶6?�Jixx��|          �#�˩���������.j��k;  v�����6������|�S�����u  ��[���JkVfc4::�H�f��         �
]]]*
��_q�������  ;�"�/��*�_��*�)P(���:4�磉�']�  `�{�:3{�����~�r9k�         Tc�FFF�ǭ̏�"���1�ͪ��  {Lm_q�$}Tڗr�w�\�<w�|�.�:  [������������6         @����1���ΞF�,�����y2�����HN��:�?
�������/t�u��u  �j��N�g��N$�2         @u���WWW�����Q2�am> ���$;@U���J�)��Qpǫ:p��D��[l=I
 �-�~��f�?ae�K���j�iZ          �Aoo�����N$c��~��ne> ���˓��H�	�A�}Qpǫ��:�BS��W�  XR.���}w�\��*������[�         ��c4::j���h��Ғ|+� vx5�]�y��k�!�}Qp�O����k�z�or� ����w��✕�uuu���2         @uJ$�6ߵ�2�Uk� 6��%���K�*���΁퉂;����������� PYfO���G�̎F��15��,         ���Ԥ��v+��M�m��+� ��U�5�hD忕�q�OMf�[���ۺ���9  تo��g���fe�������          �_�R����{�P�ѷ2 `��j���d.���?s��w���XyCkW�\�  `���--�2���I---Vf         ��HD###V��x�w��Z	|6 ���L�Wy�2Z�=�s`{���
��C��X]Y���࿊ ��ՕUz�+��񸆇���         P[����������kV�pN�JV� �0J������e�#��8��;~����Qh�ou� ���糟��꒕�###�F�Vf         �=;v�P6��2��7�+�\�2 `�QTR�u׮�iϯ��탂;$I�-��u���:  [���O�ř������P�P�2         @m2�httT�|u+�I��+zT�z� �Dwa;��.�H3$Qp�$����Ss_�D#�� PQ�e_?���K��b/�N���?�          �N����ge��Kz���I�� ���{CD��r�w�[O�����M��s  �U���E���>����+          @�:;;U__�\�3z��c*���g �1J����/�}9��E�9���wp�o�d��:  [uznA'��잞�r9+�         �%����F���mm����&��|6 ������;�����^�*
�����m�L*�:  [����T�\|n6�UOOO�s         �����̾��Q%2E+� v�]G�:ʊ���p��{���ܻ�{:�t� ��z��Ojq�p�s=���訌1��         �����E---��M�b���>���l �\q?Ǘ~7�����w(�ר�����~�u  ���}�������g���+�N>          ~���A%�����R{OB��l ������y���Ҟ�� p��{������|C]��  l�C_��ξx*�BA��         ��'�jxx8��]yݨ�> `�'#zݒ&s�?wnPp�A�}aywkG믻� �V-/.녧��\[?,         ����Q����F/j��R� vx�K2�c8�K\���\�@�(������3+_�D#�� �8���y��,>whh����          `+����N���wߐ��b�s �x2��ᜑ�em����s���[s{s��  l������S��miiQsss�s         `�<���Ȉ�	�ve2�E�u�%w �F	q�]���r��=�S \�k���-W��#�9  ����E�67������s_          ��\.������N^ҫ|��\ �FFW��3]О:�)
�5d���[�d�u  ��;߸W�/N>w``@�85         �^����N���yFW\=��V� ��+��oH��u���{����/�v���u  �j}m]�?v�s����\          x��1�1��w���?#��\ �\q�1#����\�:�A��<<�=�|�u  .�7?���K�ΌD"
t&          )�ϫ��=�����> `W���|鯥�F\�}�k�������]�  `��N�j���;00�D"�\          R__���d�3�Y��j���@� �8w�=�:�v�'�#��u�G���=��O6w�~�u  .���?��f1Йuuujkkt&          ��D4<<��ˮV<��\ �-�_�K�6��;\�]ܫ��������#��  T����V^<�L����          l���Wkkk�3���.��Ge�: `��'Oq�1���'��\��]ܫ؃G��ECK��  \��}I�r9Й���J�R��          ��[l���W�FI�� �%.��c�d��M�s�
�U��E�1����  \��r����:3�˩��3Й          �H$���`�\z�Ѿ��U�J�s v��������'�:��^��O�~$�I%]�  `�6�7t���i���Ȉ��9V          ����QMMM���1Т���|�vm �-q�;�/�I��u�A��
=2[������9  ���~��kˁ����Q:�t&          �mhhH�X��j�p��: `ǹ+�Q�1���+�ݝ�C xܫ�������g'j ��̂�_�a�33��zzz�	          .�b1:�И���&�*: `�����I.��t���^ezv�����* ��<x��(�6����a��         �j��Ң���@g�}Ðb�b�3 �x2
�m��H����\�@�(�W�C�~�KD���  \�G�kq�P�3;;;����	          �)�6/��kץ��L �=�+�?�����Z�U��{9:5���t�u  .����66��aI*�Rooo`�          `�������t��=�Jו�	 ��p����s�����*����;[�u  .�3�pPg�t���<�/u          T���6�����E�]ti��Zl& ����$_��u��9Z_U��ܙ[#шq� ����&�����ܬB��<          �n�1�1�U��v����
 T�sW�#�clFJ������*p�3����y�u  .����VO6/�h`` �y          �]e2utt6��.�׫�V�	 ��(�:¶�K��N{op���
�����_�� ��(��z��oz����W�8�`         P����H�ۢ���=. ��W�_�,�/�k��s����^�O��y�>�w� ����_������}�           ����rm�ѥW��w �\q�G&�Z�m�!��Pp�`����M| *Rqm]Ӈ��̡�!c�	          �]ss�
�B`�z�Z�ޓ�Tl& ��sܹ��rF���.kt���{;ub���X�� ���n���r`���ڔ�&          j���</�*��oR�p� *�����M���?r�rt�����MMmM��� ��8�pF��6/����/�y          PiR��������^�R�    IDAT��|��	 ��("C%�'���hϤ��0|4W�����q� ����oWis-�y�����b��         �J��ӣT*ؼ}W�H�J`�  �ѝy��'����0�+����?���\�  �B,��iy�����y���6          *�1F����ͫo�j`�A�6�	 ��(&#�:�vs]N���ul�
sp��Ig3��:  ��;�P��Ȭ�8          ��P(���)�y�^9,]l �#)�:�6d��ڤ��
�fnv�����  \���3Z�?ؼ��Ne����         @5P$	dV.���V��@�����J}Y-�K�!�5�+ȣ����s� ���]w�����X,�;v2          �I"����{�*�\l �#���ې����u
�v�+������叹� ��:y|JK^o��           T���Ne2�@f�Rq�C���ޝI�����=yUU֑uWuu�53��43j� �6�10ư 	d�a�d����8�6,v�������x�aL`c��X#�F����H��L�wWב�}�f%��<��Of��11����w��]S�����Q�@3 '���5RDs/�_��A�����r�GWɝ z����k��W�_v,--���Z)g      L��R<��c�����sј�/�< #E%R�r�9)���?�;�Qp���b�RĿΝ z��>n^�l)g���0       ���j���f)g5�j�7�%w�Q���;�(Jſ��ǂ��8ع�s��V� Ы�J��~��ɘ��)�,      �Iw��٨V������sQ��-�, ���)�q.��}�Sp4����b}zv�gr� �^}��/��k��rV�^�3gΔr      �q�h4�ԩS���Oq/g� �c����(~9Ⱪ�98������ŋ�25��]���������_�#�ʜ,       p\�:u*���K9��<�)S�F]�j�	?й�h�T�Ε;�^�T�uiuţ [�|泱s��R�j6����Y�Y       �IJ)Ν;W�Y�3�x�S����JT��x>ί���)����.�?�j%�� �z�?�7���G���o      �kkk�j�J9�w=�ƽR�`pR�"���,��;��>�>���_\�\{g� ЫW������/�r���J,--�r      �qU�`��z��IS��C=w���">8ϼ=wL�}�jQT�^���� �����R�����G)!      ��677�����E��r �S�F�)�RKQ�b�<���:�򍿽����; �����w���u��ɘ��)�,      ����ٳQ�V�>�9;o}ǆ)� #/E%j�C���Z�o˝����>b^�P�U��; ����������ϩ�jq���      �h4�ԩS������F���0�R4rGY�(�U�{���R)���/���\s.w ��_�B�4���ٳQ���      �L���1==��9�٩x���Mqy�H��?̓�����WSp!�T�\X]�@� Џ������7��8q�D	�       �J�J%Ν;W�YO?��)� c E=w�����8�̝�/Sp!W/^���z�-2 ��7��z���|)g=�裑R*�,       ����Z�Z��ϙ���7=�E에
�AIQ��6�0'oF�T�|�+uD�t�xjy}�;s� �~�ޯ��8����s+++���TB"       ���c�}4R�w�Q���;�(���xv%w�Sp�/^���1� ��k����k�����Ri��      �����bcc��sf�Mo_�"JH���#BU�!#~>w�Sp�_����եw�� ���������������h6�%$      �(gϞ�j���9O?�HD�w�Q�""E=w�Q�S�x��!Pp��W��z��_ɝ �q��ݸ~�3}�S���̙3%$      ��F#����>ga��_��v�� ����a�h���!Pp���{?<ߚ?�; ��w��c�έ��9u�T�j�      Щ�����/<����8��%$`p*�B?��oƻ���Sp�襢h�����s� �~��ۋ+����9�F#N�t�      ��U��8}�t��o����fD��``�)T��/r�8��3���͟�kͯ�� ��o��?��;��>�̙3Q���       ����������w�?��)! ���I���;f��o͝�8suf����lT��,w �G�]��/?��9��ӱ��YB"       z�R��g��}ΙG֣���0����J�_���;�q�'�Lnܼ�Off���s @?>�߉�;W�>��ٳ���      rZ[[������H)�׽�)� #����>Lzf.����)�+���Z,N�����9 �_����FQ}�1;;kkk%%      �W)�8s�L��<��혞k����I���;�HK��E�y���3����_�jNO�� �x�����{��>�G1�      `D���D����j�o{�D�c��T BE��(��G�#�CG
�C�ɋŉ��֏�� ������h�����j���RI�       (�ٳg�>㉧�F�q��0 P%"j�C����"�q&w��F�}�޸t����u� k���W�`�B���"       ���j���r_gL����o_�"�JJ� ��~�����@�Ǎ���p�8�����r� �~}�?�z����uF��      `0Ν;)���x�]碨�-) ���I��PE�h5�i>w���9DW^��+�Z����v���ع�J_g��Lo      a���������f�}�RqPR* !��~�՝����!�e�!y�J����ʷ�� ���_��qp��#����bvv��D       �ٳg�����3�wJJ�`(�%E�������9��!�v�ʿM��� ����Ǎ7���3Lo      ���q�ĉ��X�\���fD��t)R���1�ZE����!��!�إ��ŵ�oʝ �����/q��;�8q�DLOO��      �A:}�tT�վ�x���h�ݒ0��N���xf3w��@�}�]����$x�����_�V����%�      `��F�<y��3�>��U��FY�jD�a6E��s�8��#��}ym���9 �_���'���}�����F��D       ���v�j��SJ��'OF;
�r%S�;�">Њg���1���(�t����#w (�g>�_��n���Z����v��       �Z������~2�S{%%`*�S܏�h��?�b�)��޳���X� Я7��z��z��3����^w�'      �8�w�{�Q�G޺E엘
�r�H����c�o�ǳo�b�)�ȯE�Ν��&w (�s����{o����J���      ȧZ�����;�>�t��D ��{Gj��;�$Sp�G/�wnaN�����s/n_������ڊF�QR"       r8y�dT�՞�/����ə�h�
�R�/���x�|�K���8 EQTvn����9 ����K�ܽ���J����%&       �Z�[[[}���S���?A��KQ�aT#�?�bR)���o�����& �K/������M��      &���v_S�y󉘞/JL@��Oq�h����{Ɋ�H�o����9 ��y�S��s���)%��      &H�^�'N���RI�'ND;vKL@�RT"E�73#�"��1��K�����Z^<�; ������888�y���fLOO��      �ܶ���R�z��'�DTvJL@�R4rG)⽦��O��DEQ���o���9 �ׯ\��ۯ��?��N��      `�4������MřG����0X�'��w�ZD���!&�+�D�_8�������9 ����{{��1���az;      ��:u�TSܟ:�[b" ʕ"E-w���"�.����9&��{�n^��rg �2��E\~�S=�7�      `�5�����y���+�Z�FDQ^( J���;¸�F$S�K��^���������s�s @>�_~/�n��}}=fffJL      ��9u�T��zڛR��=��Wr* ʒ�)��c���S���D��B��$��]�7�3 @Y�������v      ��ajj*N�8���ǟ؎jc��D ����U"��;ĤPp/��_����k˦�0.}�b��\�y���Z4��      0����>5U�G߲E��
�����06�Oq�m�sL�ܾu��v &�G>��coo�����      SSS������'�:�[b" ʕLq�\%E��s��
�}����X^[y4w (C�]ĝ���y���j��Ζ�      �Qw��鞧���/��ə�(�@iLq�F�x�M�S�;�>ݸr��v &�'���q������      p�LOO���Z�����V���'�0X��*��Q���C�;W[^�\|����[r� ��|�������V����%'      `�3�lE��Wb �V�z�����3�C�3�>\3��	r�ʍع�Z�����KL      �8������Ş����8���(��T ���w:Tߏ���1��{�µ�/�V�ȝ ����C�s�NO{��f,//��      �q���ǟ؎v씘�rU"��;��H?ތ�'r�W
�=�q��v &˵/}����ۑR*1       �fii)fgg{ڻ���K�l ����LW#~:w�q�'�|�j�ͭ��'s� ��|�#/Ž�W{�[��c}}��D       ���'O��/�oz�f�c��D ����0�?9�Ws�G
�=�~��/��  e��s�=���ڊJŏ       DlllD���i�[�؎"픜��$Sܻ3�"�d��H�K��Z<����l� P��7n�ޭW{�[�Tbkk��D       ���R��#�/�ĉSs�.7 �Qp�N��[���9ƍ�{��^���)y� ��#��;q����nnnF�^/9       �lkk+��jO{�d��^ɉ (����mZ��b�(�w�kŹ��ַ�� e���/��/�'O�,9       �V����FO{{�fԦ�KN@�Lq���l��f��D���߸��V��� 01���q�{���+++133Sr"       &���v��}ժZ�ƹ7�DJ� �*E=w�q�~#��b�(�w�S7��fk���s @���O������noo��      �I1==���=�}���;%'�,)���ܝ�g#������:t�k���h�� �(�.��Ӿ���XXX(9       ����i�'�����0�*��t���ŭw�1.�;��������r� �2}��/���=�5�      �����G���i��v"��-9 ��0vR?)w�q��ށ���g�9�̝ ���oQE�����ceee �       �4�P{��'���+9 eIQ���1�͓�x�_�b(�Ṣ�?�; �iw?vo�������Hɍ�       mee%���g���M������~p �R�`����sg
�GH�������R� P����ŝ�7��W��bccc �       �T'O��iߛ߶�0�`TUܻVD���x���9F���nߺ��sg ��}�3/��occ#�U�      �s���=��|����O  �D
]�n� w�Q��~��/�������9 �L�/_���=�=q�D�i       �t�j�����j�8��bD��@ILq�V�=���r�e
q��/��  e��o�v�ܽ������h6�H      ������i�co9�Wr �R�z��Q�{�C�2���ĥ♥ե'r� ��]���{�gz;       �j6�������Sg�bz�@" ʑ���Q��l<��;ǨRp�K�.�r� P��.G{�J���F���        �E/S�+�g޴E  e�(��b���1�������Kk�ߜ; ��#��������'NDJi �       8.VVVbjj��}oz�V��� P���?ɝn?��͝c)�?���W�y��`]}��ޓR�'N        �IJ)677��w��R�/����)��C�����x��������(6f�ߝ; ���Ͽ��k]�[]]�F�1�D       7�<A<��޴E( ��?ŝn�(~&����Oȟr��ퟫ�jn#`�|�;����޷��5�4       G�F#VWW�����'�;H@�ܻ�����x�B����!F���WxY��~<w �ko����f��Vk i       8�z���ي�%ӁFW��{��~��F��+T�����j�� e���_��ݫ]�;q�� �       p��Z�h6��i�}l%��@" �P	7"����[g㙧r�%
�_���[�K� 0��߉�����T�����P"       ��^�=���hǽ��I��g�h�t��D��x�r�m��s� �A�u�s]�Y__�j�c�       (���f��I�o�ba��� �+E���=��f����	���?\�|�rg �A����{׻�����       Љj�]�;��j�?�D �����U����!F��{D�t�x����M�s � |����~w�o�Z1777�D       ������G޼�7�4 �!E-w��UD���x�l��@�="��q��SJ)w ��W>����      �f��V��=뛭�_�( �K����-߉��1
�}�����������t�q����T��X]]P"       ����֧ͮ���c+Q����?S�{�~&��}�߾���tc*w �O���cww��=Q��       ���ըV���{���(�ހЯ��ޏ��)w�܎u{�(���.~6w ����������$      ��U�Vcmm��='N.�Ts@� �[�JDtw�_VD���r;��O\��<�����D�~�z�޽�՞f����J       _��Al)�8u�E���~%�~|�|<���!r:��K.��� `P^���;;;]�1�      �ak�Z�lv7���#�QĽ%�_)j�#������!r:���],޼��|>w �_�LW�SJ
�       d������ӏ�G��7�4 ����c[S.A���x�\���+�Ƶ���R� �����޽�՞���h4J       ��������j�85��B�S���x7�ߟ;D.ǲ����bqva��� ��҇?wn��j�����       ���F,..v���#�ю�%�_
��I?u�_�ϱ,�����`�^��� ���~����Z-VVV�       ����������G��FU�J����.��������ñ+��jQT�?�; J�������w��7       (���j�j�O��������&�?)����H?�;CǮ���k�W�󳫹s ��������W����]�       P�J�kkk]�9��J�7�D �+E=w�1W|�b<u6w�a;v�k���B� 0H����n�;^�l6c~~~��       �3���]�?��F��ހ� Яt���e�D�'r��cu�|�J�u��ŧr� �A�s�ծ�w��       0(���1;;�������]�0 �I����oF|�t��t�
�7����� `�.}�Rܻs���)�X__`"       �N7�c����#KQ�� ЏnD���|�xo��tl
�ϽV4����?w �O=������x���r4�&      ��lllDJ���gY�":��a��0�O�N0LǦ�^����t�X�������v�~ccc@I       �7�F#���:^�}f5jS�&�)R�)����V�g��rl
�n����3 � ��܋�������XYY`"       ����f�k��J�<���З�F9    IDAT�)�}+"�V��r,
�/^)��Zj�)w �O?���u�F����ֺz�       ���J�j��!�<�E�0 �H
�}+"޿_��;�0������Lo`�}�?E����kkkL       �K)���j��O�[�")���J��Q[���8x_��0�W�K���f�=�s ����~��SSS��p,n�      `Lu3��9;KkSL@������sg��/����{c��' &��=�޾������H)0       �gqq1�F���,FL@?��{�\��_�;ĠM|��έ[�0w �?|�����x���� �       @�RJ�������QD��0\)ja(g��H?�;àMt��W�'W�ɝ �ʗ����f3����       ��� �'��Z7�`t�H�]]���˹S�D_%W.^��� `���(��t�~mmm�i       �<133���Z�'N�8 ��?ŝ>�D����!ib�/](�f�f�7w ��~���������v       ȭ�An'O/G{L@��PD| "R��2���;w���t��; �+��d�������u|g;       ��n
�ήE;v��~��D��^�0�e.���C���wwv6w ���^�x���� �       @�fgg��lv�vyu.�Lm�O�!E�7sg��,��x�x�����9 `��޾�;W:^��      �8������#�\ ���^���Z�uK�S�Dܯ]�nz; ��|쥸}�VGk���       F���Z�k�N-E{L@?*Q�aR�D㽹C���_�P����|o� 0����(���:7�      �q��P��ӫю�'�w)&�E����a⮎�J��7���9 `vo����n�f      �Q��`����h-���~T��;¤8?�<�;D�&��~����͝ ����뱷{����f��;�      `u3�m��BDt�Dt rPp/K�����P��*��R����£�s �0|���;w�t���v       ����l���N�^�v�8 �JQ���;�DH?�-ӹs�i�
����`� 0,��G���1m       0�VVV:Z�}z5"�8 ��_r��sq�{r�(���_*�F�Z���9 `X��^�h���t���8       ^��f��X^��a� ��;�ĨD��rg(������wM�Lu�� s��ߊ�;W;Zkz;       �bnn.��zGk7N�ED1�@ ��b�{i�H�ڊ���Q��)�_�t����  ��ٗ>w���hm��g      �Q�R��}�͓Kю�'�w�H�r�������!�2�n�ˋ&w ��?��QG�e^��caaa�       `8:-��<�E�8 ���01���x�D�ş���ε�?\�V&� :�{�bG�VVV"%w9      09�����A]�9;���Ы��ۭ���Q��(������� `X�ܼ�w�v��ӻ�      `\T*�XZZ�h���\D��t r1��L?�;Cƾ������[+Kgr� �ay�����۷�\���      `�t:����r�7�4 �*E�	�3���Kq��;G�����~��O��  ���+Eq������=�       ����r���\wb{)�
� #-E5w�I2����ѯ�n�}�(jSS�ȝ �����[^^p       ȣ�h���ܑ�Z��1��8	0��˖~(w�~�u�}�j�����|� 0,����޻~五��;       mee��u�[*f �L��t�܊g��я�.�_�p��sg �a��˯č7�\777�Fc�        �N��[�(b�i �]%�xW�GM:����c{5<w�h-,��B� 0L���r���v       &���lLOO�n��b�7�D ���;�DI�������+{���j5W3 �ʍ�_�h��;       �A'm��Ro! �JQ�a�<6OC��ۂ�����n� 0l�׎\S��c~~~i        ����#�T*)�6g���^)��/E�rg��X�_�^<������9 `��^�wn^=r]'x      �I�����ѥ��͹�0�`t�H�YkYE��G<6�;G/��J�~�揧�r� ��z��;;;G����k       0	RJ�O�����B" ze�{��b�r����܋�H)ҏ�� �v��W�\�R����!�      ���ɓ�7�����!��w��&N����z1v�O\�o�]�[͝ �m���#�,,,t��5       �KKK�R:tMsv*�CJ@oƮ�<�o��g��lČݕp����  öwo/�����v       ��z����G�[�l! �JQ���oX�k������[cUp�â�������s �����/ƭ�7�\��      �q����+ksQ��� Ы��&Pz_�����ε�ˍ��t� 0l������;tM�^����!%      ���I�}��b�?�4 �*E5w�I��g��s���Xܯ]���rg ��_x��5KKK��G�       p��Z��V/E�o�"���� �K�} *�����!�16��^+�͹���A�*)b��P�Xl|�����_��j����G�Y\\B       =)�#�7�7j��2=�D ��)G�}�t��;@������ȝ��5*���Z�L-������"b���qk?����_8�w�c�Ƒ�:y�       L���Ÿ|��kV7�q���ЛjD��1i��ǻ��}&w�N���K.0wz�R��Tě"oE�����wVn���n��4qj6⭋�g����{�s_��7/�7�͘��R"       =��[]��Bi`��P�"��͝�ScQp���b������sн�"6f"�ڊ�jFL��='ED���Bģ���d{�W�����5��      p�5�͘��>t��梂;��KQ�a"�H�ϝ�ScQp�I�]��\�cf�~b��t��{ѬE<�p�@_������׎\���8�$       0ڎz�|e}!R��!s �V����)�c�8���!:1�+o\�;�3йJ�83qv.�1�+,E��Těʛ0*v��zJ)Z�֐�       ��:��^�Wcq��)� �ƣ�<v��˝�#���j�����L�tf�z�d�P�����G�#���&���~�ݽq�����       ��	�˫�!$�?�����G>��ݝw�jUW�XhD<6?���SMg�#Z��9 ����^��7/�/--)       ��F�������f�R" z��ek>��M�Ce���@�mi*��lDJ��ܗ"��l�|�I� ey��_����C�tr�9       G�����E�^< y)�N�=�3e���V,-�.?�;�[���n�/����K�3��c�ڥ�}=�CJ       �拓��F+��R z�b�k�c+E�'F��;��v��}�V���R#b��'�dUIg�#�"`L��\;������V��       ��jEJ�9�l��|m�� �E��8ۜ��&w�Ì�W�֍�?�;7_�89�;��j)���x�b�֡��Z�!%      ��P��cv������O� ""R�9(EĻsg8���?z�X[Z]|G�<�t5����@���Z��t� ݹy�Fܹu��5G=V       ����-�6#�N z���6%�/��l�|d����{S�2����J�8=w���d}&b��:`���ʫq�Ν���R����!&      ��pT�}um>�8R zS���<vN��3ߐ;�Ìl�����?�;v�15�W�å���d!`�\z��Q�[|vv6�U��      �?����|�?�4 �*�n�y�Q�'w��ɯ�'/'�ߞ;_ku*b��;E嶺�S�S t�֕�����8�$       0^��z4����Z��Ti1 �1 tPR��?���h�/�4����l��1�;E�6f"*�.`��<�����!%      ��s����j���2F]Rp���x�r�x��,�߾~�Gsg૥�857��Z�ؘΝ�p�v��7]��       wԓїV'`�'��ɪ���;w�����oK�����W[������`��"�P�&���.��[���l6��h1       ���ǵ�f"�=�0 �$E��c����O���wS��)���Dg�J��=���"VMqFإW����{��Vk�i       `�LOO���ËO�+sQ��нi�����8��͝�O�����7~8w���fDeo9X1�aW/|)��x��
�       p���__^��"�����Ts�hE�����T���������ӹs�e����z��QMK6���n_;����       ��zki6*Շ�`T(�����T���]�j�U8"RDl��N1XK��	 ���������b       O��+�K�^�� �Ѫ;O�7������F�+~�ҵΝ�/[�����R��jD��;��j��z�k��      @gfgg�Z}���֒s ����63@ߓ;�W����~���]��s�sp_5E���ݖ�r' �j��݌�7>�]�       :�R������>�jDD1�@ �hd*ϓ�s�J#�՞��o�����9�oc�~��8X���o�����q��݇�>???�4       0�$��Ԍ"���^T��O�_?_��;ğ�^��k7ߟ;��+ˍ�)���"��/0����z<��)%w       ��a�/.�+���K���+�C���(��(j���oϝ��6g"�1���'܁Qr��Ň��l6�Z��       t�	f�?�4 �"�F�y�}O� b$��k���MM7��s1]�hò�\mD~3 D��k}�?t       _��h����_��i�LӠ9�ї��?J�����b�#��y��{rg�3��5E��s� �/��<����       <�a�W�f}��������CD�H�=�ߛ;���.y��v`t�ڱw��C_Wp      ���~{kij�I 蕂�P|w� #Pp����-�����9�X�Sx���Z� �_�wn�~�k�J%�Mw�      @�������|#"���G��&^�wF|K�Fq�����]��G�t-b��O0��FԳ�� ��뗯ƽ{�����\����       ��aﹷg���!'�[&���B����!��wn�������~��h8�% �W.������|���       ��U�՘��y�k���;�(Lp�v��̝!k���������[sf b����'���	�����+}m~~~�I       `�<�}���f��;��Ka��0����;C֯r�ߙ*WZf�3��1�� �{wo<�5w       ��Þ�>�lD}J�`(�Ź�x�m9d�*_�t��9?>�JD��;�蘪FT������<�{T       p���-,N1	 �*�$�aH��3���Vp�(͹�?���s���_-�)�@^�����"%߱      �W�����0Lp��Yp߿�1՘��񉨥��z���Y˝ 8�v����;�������       �d�T*�l6���|c�i �)�Ñ��B|�r�����~�ƭ�)�����À�V��> ��o\�����6777�4       0y6`n�5���k)RD���i�#�y&����^K7��I��$[���.�,kdI>>R��93g�0�b"&f<�G�e�%j!ͥ��R�<���bWwW��"��(��d��ͪ
��@���<�~����
�լRp�(��>U�DC�^dr�ҕ8<<<�{&�      ��6`n{wU�ZN�"R���FI���Y^��/U��9��B�csǓÈ�,'���~�è���)%w       ������Ee�;@G(����?"��2Ǒ�����q\>�����+�|����+'n��QNL       ���Np�G���	&����N���9���y���q\���ߙR��y~���o���a\       g���c0<�}4�G_i�Rd*�����q��"������w���q�؅?���
�P��O����G       ��S��[N�"�H�#l��(��_���}�L���ϝb��܁,N�j�;       ��a���쪵tA�"Bɽ-_Ƿ^l����xo\���}L>���NɝGSp�VUUܾy��Lp      ��<�}�ɶɡ ]�گ@o�^�u��l��M�Z?&��w�������ݼz#������b0p�      ��<��Տ���0 ,Hѳ-U��}�^������i��1�X������wWi�=в�W������Mo      �z���H)EU/�o�ˑ�̔��JQFG�cl��ǝ+
�m��������<Ǚ�~ze��q�t����N�l�L&�       ��J)�x<~`���0Z���-�=u.���6�j������o����~��a�;ж�ׯ>pex��;       4�OTo�Rp�V+�o�m��W�o��oo���q\/ELz�StG�"��;Т�WOܮ�       �;����	� ���[V��գ�u��_�oG-�L�r'��v�m�{7O�~��       �rN��>DQ<��� ��2w�R�Ņ��n[Gk��~�w�o�:���N�-��m��=�����`�
%       ��I�SJ1�V��d�q�zG1�~[k����?�u,�K1��N�-)LqZ6?x`���       Ќ�x�)��;�i XD2��U)��u�V
�o\�vv�8��6�Ń������yʀV��4�3      ���R:q��x�$Q��hm�7QE���c�����EY�Q&;>5g!C� -:ؿ������       �q���D�
�+�Q�m��s��϶q�VJ�W?����qN��<5ʝ �{�����w       h�I��Fce+��0ɸm�����Rp�z����^2�|Q���s��)�Mp�ڍ8Tp      �V����p܏���0 ,$�S��"�m����~z�z�W�sM��m�Ĝ�<3���`��V{7o���ѱm)%w       h�I�ˏ'��b�T`��H�l�*��΀�y��i������1x8���]�	�`����fǶ�F�H�/_       Д�d����xw� ��	�-{r+��Ŧ���z������c�p��g�����;Ђ�7oDU?��       ���z��� :ߙ�@7�č�Q�o��a���{M���)b��L��
�`����)�      @�>���xb�;@���6��>@���ׯV���ٺ��1x�����ãMMpZp�w��m
�       м�dr��h<�*�� �C�=��E|�іr���Ѽ��<�V/w��3�h�t���6w       h�'ߟ/�"�2S �*5[��d;�Q}��4��^�t�?5�m��4܁6TӃ�)�      @�F��۶�J@�R4\��U�_5���^Ѫ��x{�;M�GK1r!��Lp�1=v+���0S       �'܇cw�.I�rG�8)�n�v9�l<�4�m�˵&�m(bv��p8����      �i'܇&�t�	�m���Nķ�M�	��_7�oo�˝`=(�m�N��>�g       �~�~?��x�}���)&�g1ڎ�?oj�ܯ^����7�7�;V-f��	�Mp��춂;       ����+�t�	�9���WUU����f��t�&�/mVE�4m>�����m
�       ОO�O�(Jt��vU���w#��?_�?m����7�W��c-ojz;Ђ��{1�N�mSp      �����c�{}�+�.I�rG�T߈����w;�F~���ob���������`����;       d4?q���8j    IDAT�C ݑ�~Ѳ�v���7Rp�v�����~9�I�;�z0�h�ᾂ;       ���	�a/�P��|��ld�M�t�5��&����kq�"L���1����N)E��Ϙ       6�'љ��=��J4���&vZ���ڕꕭ��'��/���^܁6���|��	g8FJ�&      ����c���^(�t��U)�/"�߫{��_�0�}��}rj)"�.B�ő�;Ђ���c�?�G3       Ь�,�,?�*�뗡��-&�g�}.�}����j^����Y�>9�aa�o=܁6����       ����~��J��c�gs�G�u����`8�n����F�����L��
�`vtx��`0Ȕ       6ױ���w��I
�9���չ��߯����l���l��c�;І��ѱ�&�      @�F�ѽ�z�Pp薪��ߜ޿�;#�k��Y�9�ſ�s��P��UD���
�`>Wp      �܎Op�E���)&�g��v|�u�ւ��/����qvC��bfz;В�����       �����LQ�� ݒ�~�G��ΝET?�w����ZL]�	�����       �}����P�kRݵh��uW�WU5�}�����g7,\{R���;Ж�㏌H)E���       6�`08~{�˔��i��"�S��j+�ߺ���J��e4�;Um܁��g�{������_�       �m�,���������^��W��kg����7o���}����{m�����)>.��e       ��^/���:]�Sp�����Hߪk_��o޸�����b�����w�-U��5�~?c       �l��+KS��&)�gV|��=ձ�������W���*��f�����<�}8fL       ��X�����5
�U�Up�ه�'���V�b1E�(�����:�0�       V�����2@�T�ԢY�7"^<�n�W��4��:����d�f
�@[��'���       �u���=�:���F�1�r;���K�~X�~X̝ܰ`�L��	��Q}|�Qp      �|�߾(�$�'��"�����K-��(LpϬ��Z�܁���{�Vp      �|�߾Tp�$g�ܪZ
�ew�w�Ɠ��Su�aq
���+�-��������3&      ��v���E���EU1{��hFi5&��n�׊���<��KNj��������-}�       ����I���<�/���N�.�߾q�����\bP���@��w       X
� ݧ��_巖��ҵ�k�o�p�}���z����@����Ԕe�_�       ������=|�n�ܳKQ����X�ྵ���e���
�6��;Т��U5��      @^�'�+dt�	�Ʋ{�=�.���ӽ���l�g�{}�ہVݽ�����      ��������t:�v��Zz�7��F�y!��`�W��Z������(�m�*�      `U�{�^����W��N|�s��`�����7����G�,G����w.RSp      ��>z�>��II�v%������*�����S���X��w�UwN:�^/s       �^�=s ��
�Q|}��/Up�����2���2w ��55&�      @~ey���	�Q)���KQ}s��/\p�����d�����G�� ȩ(�����       d��'�����U���U_��~o��/�Sx��k�>�z)�t�G����@       �WpW��0���R�d+n|a��/\��r���},��[��J�O�Eeٻ��&�      @n�޿7��Ü�WA�7삦G��.�X�e�;@w�w��6�       �������_�s_)R���ݭ�/�X��Sp���Ц�`
�       �
>z�>%��tU�]	UD���]�^�lM�=(��Y� �5#⾏8       ����^
� ݥX�"���`�.6����-�8a�{��ր6�w
�&�      @~�_(�t�&�Nb��"\�}�����_/Y� ]6��       ����Sx��*�ڕQ��+�<n��{5�g��Q��ߣj��׀G���(
�       ��e)�H�w��R]U�//��t[�[���_�*贲,c0Dru       dWE��Mg�� �0]�U��Zh���/3����ɣi�.r0��7��Ӫ*b2��       ĝAu��(����K�}u�/ǝ�:ˣ�\�>��B��i��{��ր6UU�x<�       �;�'�IL�:Lt��?_y��:s=z�ڭo��14��k�)�4�"F�Q�       �]��8�Sw���]%�(�r�ǜ��~�ڍ�<�chN����hQ5O1s�        ��&�tX���WE��>����p�ų>��g~X%�	�       �RF�QL���1 X����H��\p������z��ϟ� 4���yJ�6�")�      �
�qd�; ��+g}���_����ʳ���؍��������S        w����Ms� �u�������<�L�j>;s��f��؍8�� X�<"Rr2      �U�R2���t�VH�F��Yp���.�lyh�I���5�2��p       `���� ����J)�8Ӑ��Mp���g�C�z��%Mq� Жj�       ���`�; K��Z%U��r�3ܷ�'�=[�TZ{���m�|d       ����i�f��1 X�^�jI���޽���/W��U�{�@4�w��8܁�8�      �*1���RDT�Cp���8��r�Vݰ�W�)�+��樛�)�q       `���� ��*�W��8���i�|�V���ї�CSLpo�	�@k�2w       �>&�t������������^��bqh�	���a@[z�~�       �}��Mp�>E�USE���e��Bih��{s<�@[z�a�       �}��rG �5�@�}kg�Ӌ��)J����m��      `���6���4AWOu�{�4w����1���ф��k��h�`8���!       �{n�:���)���?�;/L��;�j�{5��l"꧄��-Ж�d�;       pw��K
�h�||�����T�ý�//��&���c!Nk@[�ۓ�       ��ܺ��; Kz�p��G��i�w����/{�84���攞[�%��0R�%       X{�sG `Ij����T_��(��\����Ƹx hSQ�rG        �}� w ������
��˅�	��6G�hS���        ܥ� M��p�{=vd����oM���Q7%�攞[�Eӹ�       ��[7�sG `i:Y�)}�4�z�����\Jɫ���*�Qp�4��N        |d�	� Аs[�gw���g�٩F�ӾǾx,�t|�MG�*w       ���rG �������c;җ?��z�P7ܛc�;Ц��%K       �*�օ2�*J��/�N�RO�²k�	�@����;       ��8<��@-�AWS�����؂�`���z�P'ƛ�|�=e9�       ����n� @MRT�#p�%'�WU����<W_ �b�x�\D ��7�        Dč�{�# P���U-7��g����p`��
Rpo��;Ж�h�;       7��FRp_U���z�Qwxd��,�O��C]�5�8w�-���       ���~�v� Ԥ�*wN�߉�ӏ��#���>_o�{�<w�-�]w       X7LpX&����#;�,�_�����C],��)�m��݉�9        ;w hCZ��>����C�hK*�H�~�       ��]��; �Q]a�{�7Yp�������<w�ME9�       6ޕ�7sG �6U� <�g��G�w��<]o�w�MG~�      �ܮ]��; 5�Lp_e�y�7Zp�����xh�슲��{�� �:8̝        �j�;��H&���OE��О�C+���G����{�܁6�R/w       �h��<n\����hۮ�r7�/=���V��O��C-��ƕ�c�E�7�       6�����2� Z�"}�a�{h���{���L�`�x�z
�@��q�       �Ѯ^��; l�Y������Ϛ��`�;Ц��v�       �Ѯ^��; �R]e)�O?�{-����WIC-,����@����        ��۹# P�*w !E:{�}<=�L莞�;В�'��        ��7rG �VJ������þwb���������\$����V���^�~/��0w       �X�.^��Z���>��o�X�\�O��P�f����EU��       6֥�&��%�w�\|񉓾qb���x��8�=܁���
       r1� ����I[O��޾t��͆aY>4�=]S�Eә�j        ����ʥ��c P��m��f�N_p�|�ڗ���Ҭ�V���i��#       �F�~�v�r� �FU�r��R��'mH}7�q�a�+Lp�T��#       �F���� ��iҫ����I�O,������ò,�v���i���;       l�K��m�,�����f�@7�����SrG       ��t���� `�8������VU���e��3��&�m:���HE�;       l���+�@�������GEY�[��4�[Q��d5 -I)E9�       ����  ���o?P�;i>��-�aI����+�-�?r�      �����~tm;!�����
�����Q���=��.h�Ѽ�;       l�������r� �vڶ]0���'�=Pݽ��?m'˰��3Pp�Ts'       ��r���8:��@�R��8�"����������8�&�m�O�rG       ����{WsG ��IwAu�	�Q�?�J�w�M�O��       6��]� 6V�x���`�|;qXF墒�(�m��̓�#       �F����;�:R���4���X��,���܁F��F�c       ��x�ݫ�# Ѐ�m�	)�On;Vݭ������n/����A�)w`���\Y       my��˹# � ���x���5���b<S�J���4�[�+"t܁6�rG       ���޿]� 6ٹ����7+���B�yX�~{�z.� ZT���       `#\�r+�n�@��q+���}�����\�	�5ת��;Т��n�       ��}��v�u�j�������j����|��8,ʢk��;Ц�O=�;       lw ȯ�xx�����n5�po�@�hѓ�>)9�       @��{�r� 4Fٶ+�GMp�MMp�ˮ=
�@�RYD9��       k�w�u�e�%������B�qXFe�F�h��Q/w       X{�)���*R������A��v������܁�U
�       Ф��i|����1 h@Ҳ�GNp��O��ḙ�֘���n�        k�ݷ/�\	`-U
Up����n7˰�ړRDO�h��yל      @������ hH���:����K�n��ﵟ�EU�2�hӓ�?�;       ����֖�m�<���G7�Uvo���<yX��׮��;Т�h�`�;       ��w~�a� 4F˶c�8����ޫ즙�{�̭�V��	�M���       My�w�5�d�5)�܋O�â,�v���m�F�#       �Z:<������ �Տ����*��.^})Oe�{��
�@�[��#       �Zz���ҿXcN�]S�Tp�u�{�̬�V܁�����       `-���K�# РJ����{��{���l�|�0,��v���"�Nl��=E��       ���~�A� 4Hݳ����e����7�hQQ���$w       X;��b� �q����S'ߗU5�`܁��>,sG       ����*���*L��*���}�������E��l���)ж�8w       X+�.ވ�7�s� �AI�����>v�daQsk�u܁�M���;       ��߿ez;��3���,���Ɠ<YX���k�	�@۞y�rG       ����|�; �S��?�G��[�h0���a
�����l4E9�       k��o)��
z2"R�݂���5����zED�r� 6��Q?w       X��b� ��z���#�܇E�ϛ�E�4ܳ�� �fZ��       u�}� .�=w W���(���[p�R<�7��Y{Y��	�M39�V       �o��~T������;��D�G�Pp�"�<Lp���K�GJ)w       輷~�^� �Bɶ�RT�#��o^��\�8,jn��n���l�5�r8�       :﷿� w �\�U�c����;������w��       :�7&�l �ڮJ��
�e�{��ED��8��w       Xƍ�{���s� �qʵv.�n���ϞΛ�E��޾S܁�M���;       t�[��l���J��S*��:jjf1,r' 6ͳ/��|~       ,�7���V(�vWq>�n��,�'�aQ&��12�h�`8�r��;       t��;�������Q}\pOe���Eͬ�,�
�@{���       ��~���rG �fGwW����������U���;�ü��5       ,���ŵ+�r� �ʵ�q�����faQ&��1,r' 6��g��       :��7�-w Z���a�܇�a�,,��<�1PrZ�̧�����       :��}7w ZR)�w���� o���Ϩ̝ �4E�bZ��       8+�6�rm����(����~��˝��(��3�j���
�       p����o?���(�v�VD��3Wb;��;��s'�\&�9��?�;       t�o~�^�f�V �C���ҳ�Iѯb'w7��|�>w �g_y1i       pjo��o�# В���M�"��B���f�a�"��1Z6�7��       N��}7w Z��'vt]��b
�]����)�@����       ����_��;�c ��ڮ��l�H=��Sp�g��dP�vsG       �Nx�������1 h�RmוQmQ�V� ,g���1����_�       :��v��R)�w�,���`�����Z�ٌ{� �h���(���1       `��sw�͢T�uE�����[�ra9G&�g3,r' 6��t�;       �<�6�	�ݗ��*n߼�D� ,g���M�"J�@�`      �G��kq���c �*�����.��G�����#k1�Q�;���~���       `�����L���V1�ύ��#k1�I/w`]x��&�c       ���ן��; -�Lp�yT[�|^m��r�f�l��	�@&��8w       XY�x��# �:��K[ET��;˙G��z�fd�;�I��!,       p�Ko��]���)�v_5,�2����饈~�;���~�S�#       �J���~�; ���@R�aE1���M�ɬ�e��&ڽp>z#?�      ��~��۹# в����PE��,�����#��&��	�M�?�A,       �I�x��# �2�u��Ei�;˛Z�Y�܁L��\�       �R�}�r\��F� �,�i�� E5,�"������5�ո̝ �TϾ�R�       �R��Lo�D&���*�aQ�B�}(��U��A�;�����Do��;       ��_������i	n    IDAT�C1(�H
�k��E'ٍ{� ���l�;       �����6�2�z��E��]t�ݖ�;��`���       `%���č�{�c ����z��EJ�Z�8�Y�����	�M����p      ����� Ȥ
Ӣ�CE�����Z�Y�ʈ�;����A���1        ��_�m� d�D�F�EQ(���#k3�"EP2٫ƹ#       @V�{�����@����aQ�J�Pp�ob5�<���#       @V�x��͔� 6S�; ��~Y�NA=���< ��_|.zCS�      �\����� ȤRp_'e�Ri���8�6�Spr:L[�#       @6�����# �I
S��HQ�e�r��G��	�V�K��       ��������Ws�  ��JQT�k���'+a�3�L���+��"w       h����� �J�}��EI�}M���z� �j<G1��       Z�ڏ�; UaJ�)�����<"�.@�n�ϝ �d{�q�       Ъ��������l�0�}�EQ路��P���V�����        ���Oފ��Y� d�ܾf�"tq�ʑ�{vE���S �깗_�rh�;       ���&w 2��ENk�(R$�5r���z� ��(m�        ��ϫ�����; U&���*�(��ȝ�)��w ���ӹ#       @+~�/�č�{�c ����:IE�R��F|��J�(�=��W���s�       �ƽ��_� @v&������߾N\���ŝ/��^it>w       h������ @fU��f�"%�ur4���e%���4-wsG       �F����x��+�c ����)̘^3UD���܁����+�SZ       Xg?���� (ͮ��྆�W��;��x{����1       �1���׹# �Yez�ZRp_C�
�+aXF�'��$w       h�������; �)ͮ#�5��R���uᅗrG       �F���M���l�J�}-)����Y�|D���³OE9��       j�ڏ�; +A�})���}kuel�s' 6�a��       jut4��_�]� � �ד��:�E����0.#ʔ;��ο��       �V�������a� ��u�྆��8�^WƤ�;�ɞ|�荷s�       �����:w V���Rp_S�����Vp2;L��#       @-��*���*w V@�ྶ�ה	�c��;��v�}!w       ����v\���; +AYv])���kve�ʈ2�Nl��^x.z���1       `i?����a���Rp_S���	��V/w`�퇂;       �VUU�������Q�@C�ה��j���N l��g^�       ���?�׮�����,�����t~�հm�;�ٳ/=�p�;       ,���_� �ʨ�2�}m)���C��1,#z)w
`�ݞo�        ��*~��o���Pn_g
�k��'/���~���;�܋�#       �B����ĵ+�r� `ET�$���Pp_k&����^���{���n�       g������ X!U(ɮ�
�km��)+e�w`T;�#       ���f�����U� ��u����Wˠ����S��l�       p&���������1 X!&��7u�56�GL��)��)�@nO<}!��n�       pj�㿾�; +�
�כ���"�����������|�       p*����߿�; +E�}�)������݋H�C ��O6R���wg1��wzߟS����\��8��p2�$�0� H� ɍc$�����w1�#{l��f���gDQ��s�H��&�)�I��N�[s�fwuUW�Y�\�,�"{���y?�n����y�<���       ����C�eu�Y:�.R��=�>��3�U��P�
��&g�281_:       N�{���t ]�������ܻ��p���3b�      @w[^Z�㏼X:�.c�������{�1p���K/�����       �{=t��i6� x�F������\������U��!�<���ёd�w       ��=�=Q:��S�JU:�-ff[��]g��d�4&v�N       ����G��S�Jg �e��ց�{��&��3=\�  9�ҋ382V:       ������r����b[�5`��}܁n004���\�       x�����]O�� �+y���k�D�t�j����� H�λ�t       ��?|)��^,�@r���k`��t���u\q����]�-�       ?w�mO�N �kuJ��k�S%k>�]�������	       �$9���Gz�t ]�J'���u`�^+����L%��� ɾ�.Kc`�t       䁻�Ls�U:�.T��^�5a�ޝ\q����x�Jg       @���	 t�F�a����&V��ؕfFJ ���S:      ��{����g�(�@�r��>�kb��T�#x�顤Q: ��K/���d�       j��v N���0p��v�4���u��p�
���hdu`�t       5�nw���?)�@��r�6�kdՋ+]i���;\�4|�       ����/�葥� t-W�����FVܻ��;�-f�2<�P:      ���'J' ��*�Z1p���]ix ,]���U:      ��9����~�|� �X#�:1p���V�N�w�[�������       �F���i�\���\p��iu���wW�)] �n`p S�Kg       P#w}���	 t�*1p���������4>��4]bz�(�      @<���y���� ��U1~��ښ9�3޵��K ��Y�����       ���7?V:�.W��^;�5��*]�����d|w�       ���#Ky�{ϖ� ���\7�5��J��|���d�Q�`ݾK/���D�       ���L��*/ ��1p��N��y��+5�#w�n00�H{x�t       }������<Q:�.W�Je�^;�5S%Y1p�Z�#� ~a���i�U      ��������Kg ���^��j��N��w����K� �`zn&�1W�      �|w|��	 ���������[�8��F25T�����N       �ϼ���<��+�3 ���d�^C+�S���dfGJ ��y�_����       ���n~,Ue���U.�ג�{��d��k�'�� ��=��t       }bm���z�t =�������V|cC�l$Så+ ~a���య�       `����Y:�R:�P�ص��kj�U��S�5p����p��Kg       ���`� z���ue�^S��mf$i�� �%3�/N�L       ��g�|-/>�f� zD'Ʈue�^S����Ŗ�5�H&]q����\Fg]q      ���v� �U\p�/�����D�t�2k�t���}�       �Qǎ.�<S:�Q�ך�{����]mv$i�� �%�/� #�3�3       �A�|�4�.rpf��;���kl�g��6���� �bro�       zL���m7?V:��b�Zg�5v��t�����H����}�-�      @y�'s���� ��������U�����f��F��_24<�����       ��[��t =����:3p���]mh �*]�^�\�Fï       ��㏼����V� zH�N�
�N���V�Ngn�t�{M�LehfO�       z�����t =Ǹ���kn��K���H�(�+&�\�F��	      ��{�ŷ��/�� ��Ti�N�0��ku�5ρ�6�H��KW ������Y:      �.v�7���r~��Q�J�t���\�䄁{כ)] �~ó�N       �K~{1��T� z���$�$Yn�.�tf��/�t��.���\�       �Э�?�v�^ Ύ�;��;I�ܻ^��>r�6��}�       �2'��r׷/�@�bԊ�;IV;I�˒]on�t������O��       ���q�c9��V:��S%1h���$U����]oj8����@#���      ����䶛-�@O2ng��,I��f����p����uɥ�5       $߻�'y��� ��*��	t	w�$�=z��h������y�3       ��\�H� zT�v����;I��N���]o|0�����20�k&       ��������t =�JCV֙ʒ$�Tɲ+�=av�t�����el�w      �:����N �G��۫�t	w~���7��]jz�%i��       ����3O<��� ��*��	tw~{OL��G�.4>=�񝮸      ���_}0U��. ����_0p���:�?t���� lr��i��      �N^{�p~��gJg У�_�r��_�@��:Ur��'̍$�� `rv&c�Kg       �����w�x; �����y�%��0�HfFJW |��]%��       ��k/���{�t =�]:�.c��{7p��@���1�����3       ���!��ؐ���_a��{4;�Z�tgbj8�	��خ��p�      ������y�^��؈����1��=:U��{Ϙs��Rs�vftnw�       ��u_�^�m�48w��|w�g���g,��. 8����       �"o:������ �8w>��;�s��T�#8##��P�
���oO�����       `����\o`ê������>�N�ꅘ��0R� ���w_�F�Q:      �M��[����� ��UI�,����>U�%/��ّd�v�R��vfl~o�       6�_(��A" �z;'c��:�,]��h$�å+ Nnt�E��      ��o/��۞(�@��.�@�2p�-��vU��35?Z� ���v���¾�       l����4�� l��;'c���T�	���3&���f��M�$q�      ��=�����z; ���x?�X>P��+��W܁n6�0��]��       `n����\3*`�\o�T�9�E�������md�����w      �u����y��� �*F����;'��N�|�C�H��KW ����\&w��      Ћ���Y[5F`3T.�sJ�T�J��N�SFK ����K���      @/y��c���v 6I�N��t]�S:�,]�٘NF|��.657����      ��o|�4�.��Y\_��La9��-����yW܁.7�����       �����y��� ��t�)N���Sju�^��)#I�t�)�OOft��3       8_���T.d�i�����0p甪$��=eh �)]pj��_��a+      �n��Ӈ����/�@�b����sZ������Q�ˍ��elׁ�       ��W��7��� l"w΄�;���N�������dԧ�r�\�����       |��~�B�|��� ��*UR9=XN�S%K^��9� Nmhx(��..�      ����*_����3 �3��vwN���3r�Y����0�4JG ���/���t�       ~�w��I^z��� ��v� z��;g�xs��;�c��̎�� 8���@Fw��      �-��N���Jg Ї��J'�#�9#�*Y�\�9�� No�26�P:      �$w�r0o:Z:�>S�J�;g���3R%9n��s&����� �7�;      @q�+�\��Kg Ї\o�l�s���8;\qz����_�S:      ��n���=�T:��d�Ι3p猭u���s�G��F�
�ӛ�wy~5      (a��Jn��� ��*ITΜg�S%K^��9�dn�t��M��gjυ�3       j醯=���+�3 �K�������sV��8;�J �����g`h�t      @����|�GKg з\W���sV�[I�S���52�Lۋ=`d|,�{/)�      P+_��=i��5:i�N���sV���ȝ޳c�t���;���O��       ��g�Z���� ��*�$.+sv�9kǛ�8����`�
�����KKg       �����Oߕ��J� Ч��r��9k�ͤ�wڞ�;�+�?�љ��       }�;~��9T:���*@2p笵�d��'͏$��� gfb��       ���J3_���� ��N�tJGЃ�9kU���=i��>r���vgb���       }醯?�w/�� ��U��s��9'�ͤ�JWp.v��. 8s{/Kc`�t      @_9��bn���� �9wΕ�;��I�ۥ+8#��p�
�3357��=��       �+_��{��jt�V�R�Дsc��9�T��f�
����� gn���346Q:      �/<�����}O�� �Ϲ��F�sΎ5��t�dj8,]pf���3����       =���|�3w���~ �Z�l��;�l������Y;\qz���2>��t      @O���'��ӇJg ���Ti�����s�:Ur���g͏&C� @�<�4<�       ���j+_����3 ���q�o��Y��!��Jp�q��-S���{�t      @O�����ۋ�3 ��*�'�1�l�j'Y�-=k�h2�(]p�λ<����      8��^̷��A� j����2pgC:U��,]��l$�#�+ ����h�Ͽ�t      @O�{O�V��z����t=���3p�m;�G܁^2����Nϕ�       �	O��<t�ӥ3 �	����l�J;Ym���\�$3��=��hd�+Jg       t�v���?ug��%] ���;����kW�qϣ��s�t�ٙٹ;S{.(�      ��n����Jg PU�I�T����)���.`#&��ɡ� gg��+20�+(       >��s헿[:���,�@�0pgS����];�J ��щ�L￼t      @W��Swfu����S�U:�>a�ΦhWɢ߇{��p2:X���̝q�fJg       t��y1��� �����*�A�0pg�[+]�F�-] pv�F�.�p~�      H��Z+W}��� Ԍ��l&k06�j'9�.]�F̏&C�
@���_�Ԟ�Jg       t�k����y�h� j����d�ʦiW�b�t�H��w��^���M��       (��W����.�@�T�#�#�l�ckQ�n�h2�(]pv���3��C�3       ���㷥�l�� �f:������Tk���TOl$��=hn��X�S:      �����q~|��� �N����Mf�ΦjW�b�t��w�GM���4Kg       l��k����-�@Ui'�Jg�g��tG�U�nh �)]p�&f�3����       ��+Wݛ�G�Jg PC�����t�N��y��v�%���h���325[:      `[�����փ�3 �����-a�Φ�T�b�t5<�̹�����@f.����5      ��UU����t:U� jh}��� 6��;[�Xs}�No�=�;Л�vff�ť3       ��m7=��>T:��r���b�Ζhv�eϭ�72�̸����?�����       [��ۋ���/�@mU�lw�D�Z��N��=V� ��g��GJg       l���X^+�@Mu���B�l��fҮJW�Qc���p�
�s3�sw&w�_:      `S=pדy���Jg Pk� �u��2���ȝ��;��f.�p�GK�%    IDATg       l��c'���]:��R�J�t}���-S%9j��&����� �ft|,3�Z�      �Mq��oϱ�˥3 �5�P���;[j���uJW�v��. 8w��.�Ď��3       6�=����t 5W�U:�>g�ΖjW��Z�
6����%w�^5{�g`h�t      �9Y^Z��>~{� j�J'Uڥ3�s�l�*ɻ���o�+] p�F''3s��3       ��>}g��s�t 5W��c���;[n��,�6��0=�L������.��ܮ�       g�G��4���d� Hb��3pg˵�d����;���Ff�F��      ��k�̟ߚ��J� PsUZ���#���;��X3�x���)W܁7>=��.�      pF�rսy��� ���v���;�b��,y����� 6ff߁���.�      pJ?y��y��� ��J�,AM��-:��w��Ԑ+�@ok4���#.�      ���V[��_|;UU�N�Ti��Hlw��b3iuJW�Y�����щ���p�      ��/ޟ7^�t $I*���F�l�Vg}�N�Z���˦�^���]�3       �㹧���)� ?�I�v�j���mS%y�����q��q�F#�^�����)       I�V�������t��) ���v���;��Dk���01�Lل=nd|"s�z�      �$�7�x^��;�3 �g�tb���2pg[���y�ʞ�� 7����.�      ��3O�����A� �%�����1pg�[K|�R��J�]q���%Wfpx�t      PS�+�|�OoIǰ�.Re�t5d�ζkVɢ+�}e�x������)�      ���?yG�x��� �K�t�*A���:Ur����������3���      @�<��gs��?*� �Q�S��;E,���v�
6�^W܁>1w�odx|�t      Pǎ�����wJg ��TY+�@M�SD��sŽ��&s#�+ 6nhx8s_�4�S      �>WUU>�g�����S �W�S�S:��2p��*ɻkIU�.a3�O�A�~0��3��]Z:      �sw|�`���3 �}��bL9���$�[�+�L#��h�
��1{���+�      ��7͗?wO� x�*I'��c�N1�*9�V��Ͷ{<p�������4K�       }�����tSVW\��5�>s�2�)�x+Y딮`35����}b|f6�~�t      �g���y��C�3 �U�e�ST��,z��]c�Cw�~0�����*�      ��}#���� p�Ti�����)�Jrt�Y�������4��_�[��      �Ƭ���?�9�v�t
 |����tw�[�$K��}g�h2�	􉑱�,\ze�      ��}�o���)� 'Q�J�t�S^�J�]+]�fk4�=��}dr��̜wI�      �G=�×r�-Kg �IUi'�-#�g�NW8�J�<���h2:X�`��]�k��-�      ��cG��?�%UU�N����Z1�����Ъ����}��d�x�
��308��4�C�S      �QUU>����#K�S पt~v��3p�+TUr��t���wf��	;P���NNe��_/�      􈛯�A~���3 ���4K'����5���q�Ǿ�;�o�����Jg       ]��g�_��t �Rw���;]�]%�z>��ɡdz�t�暿�#�(�      t������nJ��)� ��������;]e����KW���'�� �hhd$;.��4�:      �����my덣�3 �\o��Xd�UZ���Z�
���`�0Z�`s��.d���Kg       ]���˃�>U: N�J;U\&����U���۾�/�O�q����g|nW�      �K��������]: ΐ��tw�N�J�y^���F�k�t��j4����28�      u����_���i��J� ���1p���u:U��Z�
��αdē�3#���q�o'_S      uv�'n��.� g�2n�K��ҕVZɲY�R#ɞ�� �ob~g�/��t      PȽ��(����� p�\o�[�ӕ�Ur���57�L�� �|3�_��{Kg       ���kGr���,� g���S:>��;]�Jr���yv��}��}��H�/�2C�r      Pkk����n��	��������Z������dv�t����}4��f     @|�3w���,� g��*��pR�Wt�N���\�ӟ��'�� [`lv!�~�t      ������q��� pV\o����՚�d�s�o�$;�JW l����fb���      �y����_�V: �R����.g�NWkWɑ��l��cɐ3�@j4��K����x�      `������}����N���>n�Jg�)���V��R�t[e��������hv�����`�      `]��;�³o�� ��V� ��g�N�kw�wWKW��F�1�O�O�M�e�eW��       6�����y�t ��*�Ti�΀�2p��UI[ɪgj�j$�?Q�`�L�>?S{.,�      l�sO�?}g� 8'U�J'�1p�'����j_�JfGJW l���?�ѩ��      �9:�����؍i6]i�uR�U:Έ�;=�����]�.a+�O�+ ����`v\�;�6      ��N����覼���) pN:i�N�3f�N�h������]c�+ ����Dv^�Ѥ�m      �%_���<�×Jg �9���!��v����8���v�&#�L@�Xؕ��(�      �����l�u�å3 ��UY��%�Č����N�{���4�}�+ �����gbǾ�      �i���|�OoIUл:Y+� g����Ҫ�#��+�j3���p�
���h$��V�ǧJ�       '���̟���rb�(��U����5����v��*]�V�7�4JG l�������G308T:      �UU��vk^{�p� ؐ��;�wzN���bl�Lv��� �Zcӳ�q�o��       ~�M��~���� �!Uک�.�g����S%9�LV=s�ޞ�d�S
�s�;�g����       ~��_�׿p� ذ*�	ӛLG�I���:h${�JW l��������3      �������Û��T�S `�:��*�����ԩ�ŵ��)]�V[MƇJW l�F#Y���OL�N     ��j6���߿!ǎ.�N���N3p�g�U�Q��Z8o"i�� �b�C�����,�#�S      ������y��C�3 `T������Y�*9�Lھ���_r�w���u�G�O�      ��[�>�{n{�t l����ƕ�.wzZ��{]�O�<���ە���t      ���G^�W>wO� �$U�f��sQzZ�J�]�Q4�}�+ ����K2����      ��^�p��oJ�c}@��JeUI�3p��v�EW�kan$�*]�=�.�HF��Kg      @�:���?���fyi�t
 l�*�T����y�Nr��6�O$�� �`pp0s��f~]     ���nw�pC�x���) �i���tJg��YL��$'��R�t	�at0�9V�`k=���������7�4K�'J�      @߹�Sw��_.� ��r��>�8x��JG�F5�̍$�O�.a;t��cɚ̀>����ۿyG����������?������1��      6÷o�a���;Kg ����N'˥3`S��7�����P���b3y�x�
��{�ѧs�U7��_�-+�+������������6�     @�y�ї������ۮ��_:9�*���)L���Nrx-9���kaz8�N�5K� ���cK���;s�g�ͳO<w�����}8{�[�����6�     @z��#��?�Ѹ��S�c�N_1�oTI�7��v26X���"9~,��
�G�������r�wemu�������ٻ.����      ��������,/��N�MW��v(��W���F#�1��(]�vyk%9t�t��?z<w\{W���5y�G�o�55=�����%���nR      ��v��?��o�G���t
 l�N�Y*�����32�\4����^U�g��_��&O=�tn������d���]���B�����O�l�?      ��U��=���X� �UV�I�tl*w��@#�1��/]�vYn%�-�� �ŵ�o|�y����Ϲ�w.�?�ݿ���Ɩ�      �n���|��w�� �-Q�J��1�����֩�c�dat��;�obh���w6�@2�Y����o��w���������_}_��������     �^�ԏ^͗>{W� �2UV���K���f'9���qŽ6�������.�b����y����'������7~���w�B�����g     @�{��#��w]Z-C �U�*���%��K�*9��+�î���@#9o"y�x���u:�<r�s��n�}ߺ/͵����7���-L�7�@�      �&ǎ.�O��5Y:�R: �L�f�~;}�q�p������F�kl�����Rrt�t�o�y8������ߘW_x�t�{����������.�      ŭ���������S��N�-T����ӯ��kc�����P�t	ۥ�I�>��=ـ��k���|_Z���J������?�'ٱk�t
      ��T��߿>�<�\� �R����j��2����F�{,��{�YM^Y.]���x����n�k/��U��,�_~�gbr�t
      ��Oޑ�nz�t l1�����������;���br�{�-]�����ʇ�����,�      �ꆯ=��]}_� �rU��q��>g�N�l${Ɠ���Z'y�X��N�7��-_�v���y��޹�~*��]�����4��     ������ݜ�
�>W%���*��)���J�VkWɻk�܈+�u22��K�(]t�_��~�M���j�N�T��T���������)      ��~��+�ԟ�b�@M4�۩wja��YMv��.a;�K��%'�k�
��w��[���\�7����o���R�����O�����)      �e^{�p���_�f�0 �:�Re�tlwj��W�G�!W�k�������c�_��O�_k?�/|��,��G�Υ�S      `ӽ{x)�{�����) �-��RY�Q���}?�0�Hv���^G�N$o��Y��C?=���)7�[y��;�s�ʿ���\zž�)      �iVN���������,� ۤJ'K�Ԇ�;�2>�\4�{�t��c�Z�t	��:�N�o�Z��7ޓNۇ>Iff'��Gٳo�t
      lX��ɟ��k��_*� ۦJ3���J}�S+C�d�+�J�_��נ���[���n�5��6o��B�ٳo.�����ى�)      pΪ��g��;��'J� �6r���1p�v\q��ח��WKW ��������~n��]k?CW�������?���P�      8'�������+� ���v�����j�_p��{�t���cɪ,��W�57]}Sn�ҷr�wK������~��g��,����δ�,��`M�z��c�FQ&�_4���&FM�h��Ēs�&FE�"��^wiK��,������|��?VTʲ���9��uy-�u)3����>y���O��)/      �ˍ��8_9�� 0��$uR����'g�N��&��%=]�k�L]��Y���x�h#c�����3����oO�ټ�v�-�侀��7?�t
      �;n[�ӿpu� (`Ը��d�NG��-���w��=��Ӓ�#�K�G�jɪ\���]k�`W]z{f�5=���*�      �h��k��O�O�i�@g�y�}�ta�NGj���>}I�+���I�X2��}�匎��+oq�}�����}y����)      �V-ߘO}���Љ\o�s�ӱF�d�+����1+Yڿ�)7���KV��_�˾qE�nt�}2|��2sִ<���t
      ����� ;�K� ��s��Ng�N�j�;w��=��Ӓ�#�K�s��^V]�9��Wg��3�c_:      �ۖM;���m[J� @!����wn�&�su7v���Q���:Yܟ�4K�@gY�hE��教��˳mӶ�9���'���W��_9�t
      dG�p>����f���) PH�fw:��;oZwrԬ���yǓ��;���sFFF��+��Z{��1�/��?��xP�      :���xN��yY|���) PL���-�E����~}ɡ3K�P�ڡd�p�
���/\�+Ϻ*�vY�m�^:��1g���_�C߷t
      h|��g>vq����) PP�f�d+�����z����鮸w��N�'#��%05<�Z�m7|�t��~�}�u����J�      �A�����e�����S �(��a'w��+���%���ޱǓ%��+��-�sQ.=�\s���,��n:��}�'�.s��Q:     �P�uN��5�ւ�J� @Qu�T��Cw�oӺ�#f%3{J�Pʺ�����^\k�����C����&�g��N     `�;�7��W: ��3���vHb�������M��*]B)u�%ۓ�f�h}��pa�:wA�:{A��z����O�����+����/      ����ߚsϼ�t ��*���v�����+9|f2��t	��4���I�3#�������2�y��K�0	��o>1�|�����U:     �)���~�S>{Uj�% H���+�-����d�����;��δq8Y;T�Z�=?\�yg����_���pt���iy˻_�F�WF      &���kq>w�T��@v^o(-��t ��:�P3�K��ޱ����;�K�@9������r��fѝ�J�P�-��${�33�{��N     `
����O�7n���2R:Z��;���*�<��[���Yɢ�IӿO�a\k��\~�m�6�7����N     ��-�障��K3>^�N�Q��K������I��d�h�O_�J��J�����/t�������s�i�d�]�K�Т.:�;��j�^�[�S      hC��^���32<V: Z�������A�W��dNo��{�ڧ/�>��a���־�k2<8\:�6p�7����g�N     ��,�gm��.������4]o��`��N2R%[F��������g&��ɘwGc���Z�ŧ^��?ZR:�6t�7��Օ�_ul�      ����^��A�v �u�8H	���x�lI��Mz�J�PJw#9bf�lG�xl��~չWgd�[�؜{�M�6�'/:���S      ha+�ݗO|����7���y���Ux(��0ƪd�Hr���%�4�w�%�M6����v事��O�(K��tSH]��ڗ�OWW#/|�3J�      ЂV-�h� �N�l���x�lK��K�u����Cg$��p�t	<����_y���d{F]�9�Kץ�Օ���s      h!kWo�'>|A���N��Sg,����3p�G0��+��,]BI�FrĬd���.�k���\�����J��!��W���L�֓�~�SK�      �ْ֭���ٶe�t
 � ��aW��#h�Ɏ�dp<�韘�6�;9xF��洈��s��?ȼ3���o���x�$:P]'_�̕i4y��S:     ��֯ݚ���yٺٸ L��8�
��\v�X�lN��N�c(���;x�1V��N���-��Wf���zٚ�9���s�HWW#����K�      P�������-�v�N��T�J�3���:j&�cɜ��5�6wf��?�J��I����7� �:?7]~s��\k��TU�/���֛g=�	�s      �D�7����xn6��v$    IDATn�^: Z����wn������dvOr������?���s&���s�YWe���޵�s���t�o>��y�o�     t�-�v�_?pN6��V: ZV�f��΀�a��BoWr��d�i�Khk�M#�+��\k����t�]��GyƱ�/�     ��m�`>���e��M�S ��53��v��;<
�$3z���N�]q�xu��ۓ�f���M�7�ʳ�ү���宵��z�z��~e��ksK�      �l߶sܾz�q; <�:�2T:ڊ�;<J=���Ɂ�K��
F��#��gRv�k�LeӦ���>�<��F�      Sɶ���ć�Ϫ�K� @˫2�:U�h+�ft'G�N��J��
6�$�KW�n6�۔+�Y�KN�4�V�+�{Lߴ����(O�Q�S      � ۶����r; �*c�3\:ڎ�;��F�O_r���%���������^k���o�N�I��ӕ�����o=�t
      �����s�����[K� @[��#u�t��2p��4�;9bf2��t	��Y'��'��I��q��\u�չ�K�n���9PDOOW��=��7~�ɥS      �7lω</�m+� m��H긚
���vSW#�ݓ9;i���%�'���y;�$U���7������_��%y��V:     �Ga��-�ć�����S �MTif�t�-��a7Uu2�L��&�������I��l.]BI���/λ&�zq֯�P:ZJU�9�W���<���t      �`��������Fz ��*���11p��`�J6�${�&�θ��;/���.a2=�Z��oLլJ'A˪�:_9iAF����Y:     ���f��q��-�� �뚩3V:ښ�;<u��*�<��r74�̝�,ޞ�ץk����~�W.Άծ�î��:_�����:ǽ�Y�s      x˗n�'?|A���N��Re�t��Ɲ�kLx��w'G�J�u�.�U�%��(]��06:��.�9�Θ��o�Aj_F�1y͟>7�ǿY:     �X�x}��#dG�p� h+u�R��Ox�\p�	0V%G��g�.�U�ջ��}�W�2V-Y�˾~y.���r���90e���[�lVy�<�t
      I�du>�ы248Z: �L�*�~�D0p�	Ь���d�X2��t�����x�c�t	�klt<7_qs�}u~����r�Y����x����+�     ����Ѫ|�edx�t
 ��:�I��0%����M#ɬޤQ:���H2wV��?�}K[Y�dU.����Wd�F��a2̿�{��:�{��N     �Hw�~o>��.�ب+n ��U��1�(�0A�:j&[G�}����U�t���۟����FG�r˕���]~�m����4     �,wܶ,'�8ϸ vS��X���1p�	4^%�G�����<~fvOr��d�p�̊�+s�7����_�m���΁�w�w�jVy��_d�     0	n�ea������ �;�4S����&P�d�J6'�(]C+9hF20��?��Z;��o-�+�f��x�q��2r     �S������^e� �A���	0�4��l�mZwr�dzw�Z�x�,���+e�X�"W|�����eٶy{��<��O�;�wBz�<�	     0Ѯ���ڗ��� �*������H��&sg�.���'��w^�gr�����W~;�:?�����9��t̯����+2cf_�     �)c��˹g�T: �\�fb����������x���CɆ��S���s�YWeޙ�}K��1x�����U�����)      m���uڍ���� ౪3�*��3`J2p�=��dfOr�줻Q��V�lG�c�t���Z;L]�w�����C�.�     Ж�ǫ���+�ݛ�)� m�N�*�3`�2p�=��+ٿ/9��Y~�x�,���+�ݽ�,�Ug��S��������s�Q�N     h+�#�9��y����J� ��Pe0u��3`�2p�=lzw2w��_�Ǔ���O»gp�`n���\u��ڡ�̚==��W�I�V:     �-�����Y��5�S `J�3�*å3`J3p�=������9r�_�q8Y;T�����Å�wƼ\s�u�1X:(`��޼��/ϯ��ǕN     hi۶����¬Xv_� �2��NU:�4w�}]�!3���J�ЊV$[GKW�����\s�չ��˲��E�s���ӕ����7�)�S      Z�}��� ��n-� SF���1��=��t t��*�4���M��kh5��L��;��ϻ�Z���_�����1>^��~Yv�/���9      -e����G.����S `ʨS��$q�&IoW�__rЌ�%���*Y�=i������\{�u���K]kv�	������W:     �%�������(C�x 0����+�0\p�I2V%�ƒ9}����5��i]����;J��s����]�����9@���222�?�����V)     @������s�������) 0��3n�I�;L��F2�7�;�t	�j�Pr_m���ڋ��ŧ^��?ZR:hs�����/���tww�N     �t���Os�g�J�Y�N�)�N���1����;L��NǓm���}�khE��H��Ɏ��%{�k�����o�4�#y��=!�}��     :������r}����Weĸ&��0�If�$G�Nz�khE�:Y�=�b��ض#�]��\������KK� S�ѿrx������Y�J�      �Qu]缯ݒ���Z: ��:U��΀�c��t%��%�(]B�O��gJ<�w����ν:#C#�s�q���򞏼*4�t
     �1>^�+']�o맥S `ʪ2�:���qܡ�i��3��=�KhU�F�5��+v����/<�,��k�@{�;+��W��O:�t
     ����?1?w�~o� ��ꌥ�p��H�PHW#�ݓ9;i���e�H�����u�_k��3:�Z;P޴�y�{��3�	�S      &�����G/��J� �V���$&�P��;�ە8=�Z�ZUU'K���~��������r���޻�-��K��y�[_����S      �U�7�����l��_: ��*é3V::��;�H2�{�����5���*Y�=o���UU���~���Y��/���v�-��g��o~~�     ��߱"'}����ۀ@��L�����ܡ��F2�79bV�Z����K�?aoް9W�uU�9?���)\��=��O�[������)�     ��n���9��W�٬J� �W��`���%�C�֝2c��ʦ�dM���>��s��7g|l|�# &�S�>7���?��Y�J�      <���s�������N� �uFSe�tt<wh�F2�;9r�΋��PV&�'���M�6��o\�y_�,�V����$����We��*�     ��*g|��|k�]�S �CTif�twh=]�~}��3J����$����=tDݵv�������_��=��)      ?gdx,'�8/w�~o� �U�R�^
Z��;��i��3��=�Khe�U��?�&�cnZ�)W�� �~u^�._;q��M�ޛw��<��ǗN     H�l�<�O}��,_��t
 t�:c�2\:�wh!]�dvOr��Q:��6�L��'�c���k�7^vS��͉h#]]���/�_���)     @�[�|c���/����S ���if0�^wh1�]�Aӓ���.��mMV<��oӺM�����K�nź�hSǽ�Yy����F�cf     ����+r��/���h� �(U�Sg�t� =���7^%�G�Y=ɴ��5��}�v^r߸��Z;�#[0�ɟ����t��     :����$�~nA�M�c`2�i�Cr�ZPw#�ӛ1�t	���I�C|��q��\u�չ�K�n���hSO���y��}yf�5�t
     0��u����\z�wS�� ����TH�3h5�Т����g���Y'K�'#?�>�jV�����o�c*O�<j�w��C��as�/�     LQ���9�s��.� ��Hꌖ� ��;��F��=�Q��ޮ�5���f��Es��W碯\��7�Nh{�g����=>�8��S     �)f��|�cg�b�� %ԩ~v�hE���zɜ���Khe�m�7�zUN���32�B������k��wr«�t
     0E,_�!���%ټ��t
 t�f�4Kg ��t ����d`<�>�s���r��s��/�,���X����hUU��3n�}��o��tw{[     `�}��9�Wftd�t
 t�*#1n���;��F#�ٝ9+鱩�x��۞yޔs�zy��~�7<ve��U�}Z�#���#�����9{{k     �ѩ�:�]x[�;�f?����43P:x��z��}z�C��:����O��Y��{��ݼi{Vܻnr� :�A�읿��+r���K�      mbtt<�~nA�s�ݥS ��UJ�����Ĵ������%L�u�gޅ7�3���k�gͪ��a��=X�٦�����{|�q��K�      -n��|�cg����S ��UK����.0p�6��Hfv'G�N��k�SFǫ������I�g���w��,]�:۷y+�=���������W�F�     �E-_�!���%ټ��t
 t�:u�$1��v`�m��+ٷ/9xF�&����gޅ7�ܯ^����?�f�ʢ{Vfxhd� x(/x����~���J�      -�7/�)��2�#��� �cWe(u|]�va�mfZwr��dVO������������Gǳ��3>ޜ����8�W��;�B��=�t
     PX]׹���rޙ7�6���Pg<U�Jg ���;�����q���v�1�g��m���r��W��ܳ��CY�p��8��>t����(��ݿt
     P���xN�܂|熻K�  ?S�N��$�S�Nܡ�v%�OK�^��]u���/��,]�rR_{���,_�vR_�M�ї����<��ǗN     &ٖM;��$��/� <@���+�<J�Ц�w'��Lf��.�ᬿo{�]xS�>m~�ͪX��5��~�b��)�����7??/:���S     �I�䞵����4۶�N ��X��� v��;���F2�;9r��?�u��5�,)r���,_�6[6��� �����������M�$     Le�\�����k26:^: �9u�LR�()��ܡ��v%��%�(]B�:��JU�Y�hUv�N�G=���^�޻t
     0��ƚ������W�U: xU�R�hЮܡ�M�N���r ������?�ɽ�W��yD���,�{EFF�J� t��{M�_�����3�*�     L�-�v��e�=kK�  ��x�8
����\W#�՝̝�t7J�t�5��s��E�\В�����hݽ���UWW#������:6��/�     ���du>���ٶe�t
 ��43��6
ڙ�;L�]ɾ}��3J�Lm#c�|�w�˟=/+�����;��x�Ծ L��z����w�i�{K�      �����ʙ_��11 haU�Rg�t���1�;9lF2�fn­Y�5�s].���S�7*6oڞ��+��Q=b����0��_�     `�����/]���Q� �a�K����0p�)�����N���t7J״���f�w�Ը��p֬ޘ�6�� �(3f��-�~i~���T:     x�7�礏���E��@k���`�X�
�a
��J��M�Y��}�^�9�}].9�s�Vn���ٲ��t@Gi49�U���{����d     ���޵2_���l�6T: xU�Rg�t0A�a��֝6#��[��}����O��U�;�����d����,��q�q���W��9kZ�     �g������N��c�@;�3�*å3�	d�SL����N���t;���$k�mͅg]��κ&U�ٿ)�lVYt����N�8��o��/�GP:     :���XN��U�����S �]P�N���\�S��;LA=]�>�ɡ3K������|���Ϟ��k6��i)cc�Yt����z���6mzo��]/ɳ����)     бْ֭�>>/���Y2 ��f���;�Tc�SԴ��ɜ��%���������g]�������H߳����h4r����k��w���mX     `2�q۲|�S�gp��^@��3�*�v�Td�ST#�̞d��tM#��|�ֻ��O��5+ח�i���t��Ծ< ��g��z�����)     0��u�����\|��) ��:U��Wo���a
�i${�&G�*]2y��~�7��%g�־�6mܖ��= P�~�w��<�CK�     ��տ}('�����e�S �G���$���b�S\_Wr��d�i�K�,��'��5��~�� ���+������W�F�Q:     ��%��������N �*#�3Z:؃�a�k$�ޝ̝�L�.]3��$k�l��g]�KϹε�=`Ž�y���(�Y�~B���f���S     ���u����0g�vC�M?c�vS�J���\�S��;t��F2�'�;{������n�qN��Y�څ�=���,]�:��K� t���+�x�	y�ч�N    ����8'���q۲�) �n���H��Tg���+9`Zr@���dɲu9���s������k�TU��Wfp`�t
@G���ʫ���9�UǦј
��    ��Y�h]����r��m�S ��Te$uFKg ���:������̞�%�n`h47\�Ü���龭�s:��x3��Y��a� �������o�ˬ�m��     L���s�����o���k� о�if�t0Iܡ�t5�Y����Iw~���X�9g~�b��[���X߳2cc�S :�����wB���CJ�     @�ͩ�[�[oYX: xL�TH;2���az��}��Cf�.�eC��|���򙏞�Z{���{V��t� ��������n�{��J�     @�Y�x}����ٰn[� �1�2�:c�3�Id�hZwr�d���%;mܼ#�wC�:u~��p������ūSU�| ��c����o���Y�J�     @K����򵓯����?@��3�*å3�If���Hfv'G�Jz��4�u��/������%e"�m[���ޥkKg �3��o���r��,�     ����/�wo^X: �U�(`������M�5��[�u�w�=9���ȚU&�řP�ۚU+�o�*z�z��7>/ǽ�Y�S     `�ݻdC>��yٰn[� `�TL�f�� w�`}]Ɂӓ����ת����ݓ���3�v��=��L��k6e��M�3 x��~�S�~Q�M�-�     ����ӾpM�F�K�  ��H���� 
1p��H2�;9b��_����X��>qV/\��^�bV._�M]A h%���?�x��9�J�     �348�S?� �޲�t
 0��4Se�tP��;t��F2�'�;+�nL��^�xu>��s���=���R�u�/[��[�K� � �}=y������4�E     
[�p]���˳~���) �����`��tP��;�ޮd�����6�ے�O� �_}[j�b:B]�Y�xu��{r��<�YG�-�~i��wV�     x�������N�!ͦ� L5U�Sg�tP��;�$�ֽs�>�w�?F���%�ݐ������8�BU�Y�hUv�N���{F��]/�3�}|�     �m�7�狟�<��xu� `�3�*å3�`�$IIf�$sg%}]�����������k'���1>�̢{Vfdx�t
 ���h��'<3��?������9     �����9������ ��*�&1i܁�n$�{���w�w��M�s�I��˿�ڧ����g��+2::^:�q�Q���9�J�     �#�9gܔ�~P: ؃��N�t�"܁��ו�?-9`���uUU���n�i_�$;�&�n4�    IDAT'��122�����ؘ�;@+����k�����g�N    ���l��|�S�g��-�S �=��Hꌖ� Z��;�K�w'��Lf�<��z��ۿ|-wܾpr�h+CC#Y|��4�U� ±�yr��/����6     �Du]���?�٧ߐ�q?o��m<�8�
�<w��t5������IO��|�Y�ܯ_��O�4c�.s��veɢU�*_j Z�~앷��K�ԧ�-�     ٶu0�|�����e�S �=�J��Ա-~��;�z��Y��9�i4Y�pU>�/gf�O��N���o��ūS�rв�F^|�3�7�^zz�J�     С��ޜ�٫�m�@� `��v��Y:hA�������䜓������ܯ_�f�[��{�l�ϊ{����'<�����_�C۷t
     dtt<�qS���C?S�Qg4UFJg -���9#C���|!�|v��y�ӎɴ����6oڞ��+��#�>�/�翗���S     � �Wl���eYy���) ��i��z��*��܁�v�w�ȿ����j����s3g���G��Fw�2���6l��Jg ���ܧ�MoQf͞^:    �)���|k���\�ё��9 �����`��t��܁�������\��sRU�������#���1�qL9��nʺ5�Jg �8hN��w/�S�vx�     ��m[��-��-+� L�:C���6���C�[�xy>��»>�_��'=.���$U1խY�1�m.��.h4y�q��׿���S:    �6w�-s��M����) �$�2�:å3�6`���s.Ͽ���>�_��ӝ�>���N��2:��U�e��-�3 �E���/o�ۗ��O:�t
     mhp`$�|��\�]�S ��T�3�U`W�Cʿ���������<��OIW�{��iV._�M��� `uww�e�������MOOW�     �ĝ�ߛS?� [6�(� Q��`�T�C�6a�f��U����'K~�x���C=0�67Icb��Hu]gŽ�es� ���; o�ۗ���X:    �6<4��N�!�Z���) б���X����C����G���ߺ}�?F��ȓ�����k�	,���u�eK�d����) <
�}=y�<'��c����7     ~�����O_��k��N 
�2�:å3�6c����|�3s�Ǿ�����楷�'�<����N��:H��β%�ӿ}�t
 �ғ�94oy�Ks�a~     ��g}'�]��X� @g�S��@|K <Z�0ō�������rͅ&��Μ5#G}t���q�\UUg�����o��n��������g��p�    �S-Y�._�̕Y�js� ��:US�d:��;La۷l���=��o�#��C���Đ��a��ޞ�����<.��W�     &Q�Y劋���~K��� @��2�:c�3�6e�S��e��׾++/ߣ��'�}�9`������,Y�*;�J� �f������{y�K�^:    �I�zŦ���+r��S �Qe,u�Kg m�����vW���wg��m{�����r�S���i3��k�9��*K����ot�ճ�����~?{͙Q:    �=���\=��9�7fl�Y: hu�T(��9w�b��my���.�;'�5g̘���9:�]����L}�f��Wfhp�t
 �i��3򦷿8��[O*�    ��o��|�3W��.� ��:�&�J� m�������1���gddt�_���ˑG>.�4&�����ǛY�pU��������W��7??3f��N    �1��:�^~G���/� ��*C��{�3p�)�o\����T�rO���#r��{}�&#w��a�}g�o{a�}ΓK�     �6�ۖӿpu~|Ǌ�) @�2�:�=��0p�)`�7.�'���TUٷv������<93g�.���3>�̢{Vfdx�ߝ �����>%ox�3gS     �u]�[~�o������� ZP��T*�L!���.��|�o�����~ӧ�嘧����)L1���Y�peFF��@��5{z�����^���)     <�U�7���-Ȓ��J�  -�N�*ILQ��c�m욋����T����o�}��	OxRi�Na�1r�Z�q���~Q�;`��)     <@�Y劋�����팍5K�  -��`��~�X�Ц��pA����7n���G�C>,1rg����g��U-���1�/�~�s����F��     �-_�!_9iA�/�P: hquFRņ�x�Іn��ּ�u���H�~s�h4��'=.{�ٯt
S��;�����x�q9��}K�     t����\t�wr�E���LI ��We<u�Jg S��;�����'y��-C��SQOOw�y�1��7�t
S��;����דW��s��<6]]��    L�{~�*�}��]��t
 ��43P:��ܡ��Z�"o��7g�}�K��3��裏NwWO�� #w���'��x�qy�*�    0�����oȷ�(�� �K�TL��t0��C�ظ~c�������֕Ny��?`�<��%q���g�05uww�e������vz{�K�     L9wܶ,���5ټ��t
 �F���X�`�3p�6022�w�����mw�N�mGux<���LQF� S��G�7��K�ħ�>    `"l�6��O�!7_���) @��2�:#�3�`�-���|�m΂�(��4�<��'f���K�0E���gɢ��M4�T�h$�?������L��[:    �m�z���kӿ}�t
 �v�if�t�!ܡŝ��Sr�'�Θ}}�9�G��gZ��(������;����_�[:    ��l�؟����q۲�) @[�~6n77&��;��/�V���M=��1����<��OI��]:�)j|���W��0�=��O���������)     -�٬r��w���ߒ�!G�����;����{���`�$H�Ď�H%��DQ���,˲,��S�ɽ'���Mor�4�����M��N/�RK�,K����(P\Epž�;f��?H֍-Y� ���_��<�|�� ��p�((W�u�,��HQ}�z��/j~f�:e��)/����<�)�P�xB��
2r�LU�,O��܍��fy<<S       �o�j�?���qq�:  �1Ga��Yg �2܁�D���Յ��SMU�F��Zc���H8j�ا�|�: ��j�����ߡ��r�       H	���~��Cz�r&!  ���&,=�@
��o���~�)�E��z��SѲb�d0�q��֯�٠u
 `��xu�=���/�V~��:       ̴�����˚���1  pe\��(d� K1pR̳?|F��?��X��>5mj�?7�:�q\u��kv��@�+]U����ڹ;`�       KjxpJ�������n�  �%�ļ��@
�Зo���g�S�LQQ���<��d0F� �]�����WekxS      �̖H8��G����X4n�  2�+�QPR�:@c���q����<f����V�RUe�$�u
2������Ԝu
 `	��|���;t������Z�       ��;�v��῿���	�  �A��*f� �1pRķ��7�Ϳ��3+7h��r�d8F� �}6V��_�C�M�S       `ALO��G�ޯ������  , GQ��Xg  w �;~F�dߣ�ǲ��q�G�:-/*�NA�s]W=]C����N ,�ǣ�{7鳏ޢ���9       pY\�աW��o���ٰu  �8q%��  I�s�xB�sǗt��y�s��>56��gx����=��i� �*Z�����G�޵U��:       ���9�o���~~�:  d W�%1'��ƾ���o���Xg����|566*��NA����u `�5mݠ���۵~�*�       �P�H\O����ɣJ$�  ��\%�ĳ����0��֭����"��uJJ)]Y���:y�eU,���q�[g  �Xnn��}h����N���b      ���r���櫚��N  �QP�� �k�F����5�:|�:%%UT�k��
��;���Ȕ�{G�3  V�-��_ܭ�{7[�       �$i�R���Wt�X�u
  �p�"r�qV ���;`���T�G��:#���U�t�*�d��i�v[g  �l�j������PUf�       K�#z��=������  ��\��(l� ��;``~v^���I���[��4�׫ƦY� KLN̪�kH.� +��xu�=����w���o�       K���C����������9   �J�QH ���;`�?��ԏ���i���UcS���y�)�3�������� �U��|}�37�{���z�s       d�ζa}��^Q۹�  �%\9r�+� u1p�X��}���)�[����ejll���NA�����}@�� ��j���ůݦ��u�)       2��lXO�����q��   K�UB!I	� �P܁%�G��y�M댴�rU�j�k$qEKc~.���~F� ��<�v�ݤG�r�JVZ�       Hs����~qRO<vP�`�:  dW!9�0+����XB-��?�Ϭ3�VE�Z�]�^�ܱT���/�)�  ��������_/����       �tg���w���u�Y�  �,�*"G|�@z`�,�u�����3GO[���ںj��Xe��,���~�W�H�: ��U���{�����:      @������;�/��N  Y�UL��� �4��y������i������A�E�)�"�X\m�
#�) ��}g���{�juy�u
      �����Ϗ�g?:�H�cJ  �����$1�>�K�I8��V��.딌��窱�Q��<�d�D�QG[���B�) �����c�o���R^~�u      �r�H���w�htx�:  d5G	�$9�! pI�K��Ǟҿ�Ɵ[gd���|566���Y� �8�����L�[�  RHٚb}�wn�u7�[�       06�;�����j=�c�   G�r�HC܁E�$}������m��qJKKTS['�<�)�"�몷{X�3�) �S׸N���[Tߴ�:      ��������~qR�#2  `�QH��� pY���ş>�?��?���Xk׮VE�F��;�X�FG��3  )���hǍ��WoVٚb�       �,w��/O��*�Z�   H���*f� ���;�Ⱦ���p�uFF��ڠ�e���B����  ��\�O����z��s       ,0�uu��E���ktx�:  �=�br�� �+��XD�ۯ��l���<���kUR��:YhltJ}=#� ����@<�K�߳M99^�       ����������  �ߐPBA� �b܁E������<f��rr�jl��`�u
���Ԝ�;�8�J |�uV��ߨ���)       .��謞x��rV.S  �b\9r��s
����X$g����>�?6��ߟ���F���Y� ����>�D±N ��-�*��GoQe�j�       I���'�蹧�)KX�   ��+��q;� ���;�H����{�:#�櫱�Q9^�u
�P(Qg[��Ѹu
  �y<��ȗ������       �*�p����z�{53��  �@��/��܁E0=>���W�p�:%+������Ny�S���Ѹ�/�)�Z�  R\^~�Y<�Ky���9       ��G:��7_����u
  ��p�(,Wc�Y���;��������Ym��ժ��(1r��x<���~���) �4P��H�����έ�zyv      ,u����5�;�g�  ���Ǭ3 `�1p��z����?<�m��К�k�3���UWǀf��S  i��n�>��-�t�F�       �L���g?:�W�[�(  @:p���u ,
��{����n�I�G5�U*]��:Y�u]���h|l�: �F��U�Oy��U�Z�       /��珷蹧�)�[�   $�U\�B� �h|�@�y�����.�u��٣��<Y� y<m�*W�/G#C�9 �4q�p�N���4铟�Qek���      ���;��R�~��AMO�s   .AB��� ����,���9ݿi�"! R�ϗ�Ʀ&���[� ���M��gD.�v ����j��[��nRqI�u      ��\�ՑC����_#C��  �G	%�?����'�c��?�+�|��<�MM���Z� �����1�D±N �����g�>���_��      �R��}��_Uoטu
  �ep�((W�N d>���'{T������oQ��P������d����:���'�S  i���P�>q�>��k���3      ���s��ѷ��|k�u
  �er�($W�M d����CW�'������Du�u�<�)�b�HLm�����) �4U��X�?|�n�s��^�k      ���=�'xX-/X�   \Ga��Yg ��a�,�����������@֔��������:�4?�N ����Uz�7h��u
      �2�Ff����W�[,"  @�s�+�(�.܁��m_��g�3��+T��\��a�u]uwijr�: �����/߬�-�)      ���頞}�{�b��u  �s���u ,9������#�=(���RS[�����3��\��@ߨFG��S  `˶J}��[TY��:      X2�sa=�����Gq�  dW19
[g �	�u �	^{�e��i���[����NA�x<�ظF�<��{G�s  i��d���}W;n��_ޣ5kK��      �E��������G4?��  dW	.��j\p���5�8t�:�!'ǫ@ ���e�)��&g��5$��W3 ���|^�}�>��URʳ      2G"���[����ļu  ��r��QP� ً�;p�f�fto�N%�	�\��\����ϷN4?VW��b��u
  C��u�'���>~�
��Y�       ��u]���9=������  Xp��
�e� �1p���?��i��+���W��I��\�@�HLm�����) ��_���l�}����      i�u]�|�S��z:G�s   �+G!���* 0p�п�ڿ��?k��P��P�@@9��@�����A�L�ZM ��b�     �t�a��Rwǈu  �"r�(,Wq� H	܁+�8��ܩ�i�,���E�����X� r]W�����N d�����������*(�[�       ��հ�'�?��v��   �s��q; �
w�
\8yN_���,��+W���V#w��ё)����[ ��`�     �T�z�G������6l�  �$޹��� ��� ��[��X'`LLL���SE�1rG*X�f�rss��5$��{i ��57�O��^|���;      L0l  ��U�q;���b��wp������P�_<d��ER�a�֖��� �3?Vg[���u
  �-/.��^����.߉     ��j=٣�:.Y�   ,)GQ��Xg @Jb�\�D<�}�{�Z�`U�Ti��2��=�HLm�����) �W\R�}��V��r��     ��ZO����P���   ����Q�: Rw�2��rJ���Q�,2�ǣںj�(Yi��'�p��9���y� @(.)оO\��      ������t�t�u
  �	W�w��L7�a�\���?���?��u����UCC�����S�������Q��LY�  �į��wݿ]~��      �D�����ٷ{�S   %�`� ��;p���K�מ~�:K$'ǫ@ ���e�)���V_ψ\~� ��ʲ40
�    IDAT����;�玭��ͱ�     @�k=٣���]8�o�  `��� �<��ez`�������rh� ��:�5�3Auu(�p�S  Y���@��Ӭ}\��B�u      RL��=���j??h�  `Ε+GAIl;  ܁�0�;����o�y�\54��ϷN~M$SG[�"�u
  �-�ם�mם�mW�r��      ���:�V�~��7��6l�  �"����� i܁��ғ/�_?�/�3`$??O��&��|�)��������l�: ����su˝[u��v��t�u      �P"������ԏ[4�7a�  �R�����0p.��W�Y?���Yg�P�B544ȗ����u]���jlt�: ��rsst�m���#���l�u      Q,�Ё���g?:���Y�  ���Jr���u
 ���e��~]o��b�c��E��o���N�gdxR��cr�5 0�����4����׺�R�      ,�H8��^8���h��ļu  @Jr���u �%��e���.M��j=H%+JT[['��c����LP]J$x� ���#5��'>�K5���9      �s�a���q���q�͆�s   R�+Ga�� p��hlhTl��:)��l����%1rG�	���lP$�N d9�ǣ�����;U׸�:      �`f:��~qB���BA>s   �0��r�� ��� �M{�E�����	y�^Un�#w���|�M�����4� �q]W�[�u��]����j�Qk�     �162�gvT�<��bQ.�  |G�����1p.�����~�#c����n}w����j��kp`\#C�9  �~��3���[��>�S;nl���S     @���3O���[�H8�9   i�q;o������D��ڭ�����z�v�z��}<��W��� O��Cr�:	  u�����Ӫ�]�{ڡ76('�k�     ��:.�?yKG]��G	   Ise� �sj�?K�K�{w~Eg����@
��P�����ܑ��������U� �S��X�ݽM�߽M�~�     ��ຮΜ���??��-�  �T�br�� �����Dw�ݦ�������J����� ~�X,����� �z

��s����uZY��:      #����NO?qD�=��9   i�U\�B� �q��`vjF�jo��@�����ʕ��3���u]�vkb�/�  R���ծ��tσ�iCU�u     @F���R����M��Y�   �-W	9
Zg @Fb�\�3GO�����u҄��Qm]�V���N>�������H  Ha����j�Qk�     ��F����S����	Ǭs   ��;���$� �|�@:�m�N@q]W��ܑ�֔�jٲ|u�(OX�  ��.���:ӯ��5���5�us�rr��Y      )��cD�=uLo�vN��c�  ��� ����%������������@��z�jh�SQQ�u
�Ѹ�:�[�  ���붻��}W�pY�u     @Jq]WgN������v�  ����v X܁K����/�����:i('ǫ��-+�N>������Ĭu
  I)(�k��[tσ�ie�r�      S�7����o�@�u  @Fq�{���% ,6��%��O}C-/�a��4���U Pa�2��#��M��gD.�	 �4��y���&���u�PUf�     ��B����Ԫg~rD��s�9   �q�˸ �w�|�O��|�u�XN�W���1rG����cP�X�: �K�\��ڡ���)      �jtxZ�=uL��pZ�p�:   C9J($ɱ�����wUݢ��y��9�/G�@@��)�G�F���Pp>l� �%��]���ަݷn�?�g�     �`.��sO���mJ$Z  ,W��K\n�%��HRp.�;+o��@���|
4T�_`�|$�q��3����  .KqI�n�c�n��Y�V/��     �,�XB-��?}K�]c�9   Y����\.���c�$��b�>w���3�A��>546*?/�:H��Ȕ�F���  HS^�Gۮ��]�oזm��9      I�����ϞҋϜ��L�:   K�r���u d%��$irt�:&��⅋j40rGZX�f�
���1�X,n� �%sW�[�u��]�uk�w�6ݴw�r��i     ROg۰^x���x�	��  ,.��5.�Iz��W��_��d �߯@c@y�<� )�xB]���Z�  pŊK
t�[uǽ�ZY��:     d�X,��-���G�~~�:   �J($q� L1p���w~����k������@c����ܑ\�����F�x�  3�|^]s}�>��k԰i�u     �2ӓ�z��Sz�'53́   �� U�v IS�S�	�`�HD/\TC  ��:�H�G�+�TX����!9ߗ ��x�Q��j9xA5���cWk��M����     ,�ζa���q���9%�u  @c� ��O�$�LL[' Å�]�pA�@@��ܑ&V�.W~A��:E�s  X�m��l{A?y��ܾEw޷]�����     @���{�M�����Z�   @�
J�� �*<�&\N�I�w��s=��S����y�ܑv�UOא�&g�S  Xp>�W�\_�}\�����9      MMO���V���	M���t  ����v HE\p����N@��#�p��F���Z� I�z=��]��B������s ��;j9xA-/��i�n�{�v����Oj     ��Ν��K�<��o\T<�UP  ���� R܁$�o���|�u��ܑ��f���R,�N `���kO���UT���     )&�����z�������  ���r�˸ Rw I����թ�'�3�e�#]��	uwjv&h� ��l��]�o׵�ꕓ��     �:ۆ��s�t�s��c�9   �@����} ���I�ʭ���S�3���#]����	�[�  �$JJ�i�m��w��Z]^b�     �H4ב���S���>b�  ���v H܁$=���k��@����Sc##w����y�t)�C @v�x��WWjﾫ��    @����Z���okn6l�  ��ĸ �w Il�[cC���b�ܑ΢Ѹ�:��� ��R��H�oݤ;�m�ʲ��9     �
�b	oi�+ϞҙS�r��   M0n�t��H��u�ifr�:Y��;ҙ���Єu
  K���h�u������|�Fy<�$     p	�����o��[53��  �%q�PHb� i��;����o��̜u���<5��ϳN.���z���H8�)  �X��T7߹U�ܹUˋ�s     �o�8�ξݫ�~\'�tp�   -�J((�� ��@�n߰G�`�:�$��~5���o�\�p8���A�C�  ���}����n�w���[�     �w�������֫Ͽ���y�   \6W�Br�� i��;����nT4�� �����q\��kb|�:  s�6�Ԟ۷��;������     ,�x����]:��=��[H  Ҟ��: HG܁$ݼ�z%�|��%77W�*((�N.�����z��8<�  ��z�骍ڻ�j]��^99^�$     2�@��|F��ت��u   �+GA�� ���I�i���� �|>p��+���sP�`�: ���b�2ݴw�n��*��[a�    @��:����rF��[�   `�r�*$W2�t��H��p�g�N�����QCC��-[f�\6�q5�?�ё)�  RNM}�n��պ�&���Z�     ��:ۆ��s�t�s��c�9   X`���v H{܁$0pG:���!��iozjN=]CJ$�� ��TP�׵��{�fm�Vi�    @ʛ��ׁW������ V   2���Bb� ���;��H\rG��F���Pp>l� @�Z�q�n�m�n�c��K
�s     H��ǻt��3:z���*   �U��� �Q�I`��t��zU__��ˋ�S�+⺮�524a� @J������޻I��WN��:	     ��:�����i�L��s   �\9r�˸ 2
w 	ܑn�^���jU\\b�\��9�v+OX�  ��V�\���n�-w]��u+�s     Xt�`T��lӁ�Ϩ�d�u   ��+G����@@�a�$��;ґ��Umm�JJ�#�E�quwj~��;  $���i��޻I;n���o�    ��qW�Ot�Ыgu��EŢq�$   ,��
�q; d&�@�#]y<UVU�lU�u
p�\���Є�'��� @�r�>mm��t�z��x��     �,�z��y��Uc#3�9   0�*!�q; d4�@�#�y<m�ܨ�e��S�17TOא�\� ��-�׎t�m[TߴN��:	    �59>�#�.��˭�j��  �1�� ��I`��L�a����[g "�p��=���Y�  �ֺ+�kO�v�ݬ5kK�s     xO,��#:��Y�:کD±N  @
pw� �t܁$0pG�X�v�**�K�R'2�����z��8<�  p%j�˵{�f�pK��X�     ���:�v��rFG]T$�N  @
q���u `�0p����d��rUTl�� L8UWǠ¡�u
  i/77G[�Wk��M���z�|^�$    @��Ё�[���3�����  @
b� ه�;���4�W����R\rG�pW�����N  c,+������-�oZ'��gG    ���[o�i�K�����  @
s�+�@�a�$��;2�ʕ����a���2=5���a��	�  2Jٚb��Ө[�J��VX�     �P(ձ7��r�N��!��cj   |8WQ9�� +1p����jEi�jk��#�D�quwj~.d� @��x<jش^��4j��JVZ'    RX4ש�]:��9?ҡX4n�  �4�("WQ� ��@�#�/Wm]�r�9�)��q]W#Ó�ˣ  ���6Uh��v�ܤ��$    @
pWg����W����6����   pi��*f� 0��Hwd��e�j�o���NT0Qw�"a>@ `1y��7���kO�

��I    �%�8������u���Z'   -���y� d;�@�#��>�(n�u
����`��FG��S  �
��9ں�Z;w7��]��/`�    ��u]��{g�������N  @Zs�PXb� w )ܑ-�~���˷N��LP=]C���c �����iks�v�n�u74(/�/S   @��Ё�[u��3��`�  ����QH��! ���Hwd���\��׫���:Xp�xB=]C���C  �گ���n�5�����Z'    �4�;�7�סW�jx��e  `!1n �w 	ܑmrrrT__���"�`Q��M��wD��c  
�����sw@W]S����    �j~5j?��9�OZ�    #9J($ɱ ��@�#y�^��֪���:X�pTݝ�
#�)  d��B]wc�v�iT�
y<�$    �Z���zs�y�N��9   �`�r�˸ ��I`��l��xT]]��+WY� ��q\�id��C  �����j�Q���ں�Z>��   `��N�XK�N�Ѕ3��9   �
�
Jb� �`܁$0pG��ذAk�˭3�E3?VO�"��u
  xW�<mm����������Z'   @��Л�����4��   ,W	9
Zg  Rw 	�i��uZ�n�u�h�U��Ǧ�S  �o������J;w7���UP�N   ���8������u��EM��Y'   ���Q�: ��I`�����L++��x�S�E3;To���Ѹu
  � ^�G�M�sw@��PI�2�$    HI�h\��xK���^�S\�  �WQ9�Xg  �w 	܁�ߊ�������NM"�h�o�k�  �8�Gj�T����qc��׭�N    S�H\gN����=ܦP0j�   �QD�x6 $��;����[��H�uu����S�E559�����	�  ����U�]v_�q�u    ,����N����<کH8f�   ��QX�xF \�@��WPP���z��~�`Q��	�vkzj�:  \�5kKԼ�V��Ԩ��u�x<�I    �`f��z�X�Z^ԩ��J$�$   �7�����! �4��HB"��f�����~�74� ?�:XtS�����"  �Я���w֩i���x��    ���v��đkiWǅA�)/   R�+G!��m� ����H���Y' )��󩾮Nˊ��S�E����5��٠u
  �Ly���|u��w�ꚝ�*)]f�    (�p�qaH�[�u�p��'��   ���ʕ˸ p��Ip]�U܁����Qmm�JJJ�S�%1>6���9�Q  �3�G��+W�Z5�UM}�u   �,77֙S=:q�CG�)�Z'   Is��QHoF \�@����hc�F�.[m�,�H$���!�υ�S  �Y]^��͕ھ�N[�W���Z'   �#C�:q�C�[�u�t�	�@   HG	%�� p��Ip]W7��a�����
�][.�c�,:�u5<4���	�<R �Q��s���J5��5;kUR��:	   @�pW��u��]G�i��:	   �"��rb� X0܁$0p.MYY�6VV��a��
E��5�P0b�  ���QU�5�U�Z�ԗ['   H3s�a�9գG:t�p�B��u   � \��(l� �0܁$0p.݊+TSS#��k�,	�� �=V��hks���������x�   �~#C�:q�C�[�u�t�	�:	   XP�"rŗ7 ��;��q����;p��-+R}}�|>�u
�d�����R$��  d���\�7����u���:��)�N   `$���������؛���N   ���=f �P܁$0p._~^�����g�,�q5�7���)�  ��֬-іm���\����V~��:	   �"�б�v������>��\i  @�s�(,Wq� @c�$�q�)�i��-�ϧ��:-+*�N���\H=��\s  K��}
lZ�-�Uڲ�R�uk��x��    \�ٙ�ξݫ��:�V�&�笓   �%�ʕ��$��	 X\܁$0p��כ���*���Z� K�q\�OhxpB.�]  d���e�j{��w�jks�
��#    �9������щ#�x�_��   ��UB��b� X
܁$0p����ƍ�z�j�`ɅB�t)�X�  ���zTU�F[�Uj��:�7��;   �"�'�u�D���t��n���   ��;���$�� ����Hw`a�Y�F7n�� �������8�� ��Y^\�MWmԖ�*5_W��UE�I   @ֈE�pv@�'��z�G]�#��   x���\��� �w 	܁����T5���z��)���"��Vp>l�  R��#UוkKs��l�Tæ���}�Y   @�p]W=��:s�W�'�u�t�bѸu   �r\E�7 �w 	܁ű|y�jj��c���㺮FG�440&��q  �v99^U֖֬m���\��-���EQ   �R�M��d�.����ݚ���N   R���Ŭ3  Y��;�������Wm}�
��S �HL��Ú�Z�  �4������u�]x��[#��c�   ��驠η���D��>ޭ���$    M�r�+�r ���Hw`q�|>���j����)�������(�p�S  @�).)T��
l�Pæ���/�N   �\8U��!���V��u����cP   ���r�($�ϭ|G�y�Ac�$��;��<�����j�J��L,W_ψ���S  @+)]�����\�m�Vke_$  ��    IDAT@�F�xn@�'�u����r<   ���
�sB .�Yy�/�r�S���I`�,����kݺ��<�)����Y���(OX�  ��fm��l�Ԗ�*m��RE��   �K�H8��U�ɞwF�g����3   `aĕPXb��#8
+��|Z�����;����Z�j�*����0rG��������u
  � ^�G�u��|�F5mݠ�M*(�[g   �H8�jֹ�>�9իg�	Ǭ�   ���*&Ga� i�UB	�ȕ�����;����+**R]]�|>�u
`jfz^}=ÊF��)   y��۰R�M��\�MWm�ʲ��Y   �B��B�ų:w�W�`�:   �h�"r�s7�d��kF��y�w,6�@�6���U__���<��T"�h�oT�c��)   �Y[���
5l����J�./�N��ػ�����ׯ�Gc�`��v�4m�m���_���35I=�f$����\��i�&8���x����N��� �� A��|�����o<}�G  ��.�vOI��H�ߞ� pg��pw����D�<y������@�ڧgy���t���  |8�����n]F��y��F�Q�,  ��q�,�|���1�?��>EQ�=  n�*U�t��|��*����~O�Π	��
�P����<x� +wV��+�*߿���^+�O� ��Z�͓O6����O[y�������= �k��l����_=}������Y  P�*��fq;pUU�i�����;�&p�+�����q/[[�uπk����ų7��� ���d>��^��LN��= �l�u+_=}�����,��[uO  ~�J?e���"�)�����3hw��;\�������ؘ��$���z��q� ��15=�'��'����|�󭥹�g �]������������W������2  p]U�L����)s�"����	�4�;\�������<y�$SSSuO�k�⢟�_�����)  ���;��ço��?��n}���	oZ �f;�~�&_~�2_>}�o�z�����Y  ���R��*u�L�"E�S�'�wM�W p��grr2}�Q��\����y��Mz�~�S  ~���d>^�Γ���O[��_����lݳ  HRe�}������w�x������uX  �O�2g��ͩ�����?����@�����x=���۷��FYV�}s�7���i 0D\y ����  0��9KR�=BE:)s��F�Π	��
�p�mnn�޽{uπk�쬛�v�>=�{
 �o��; ���:;  ��*Eʜ%���E�9��?'pg��pw��������N��uO�k���8�^��wu ~��������<�x#�wV355Q�, �k����~�̷_��7_��?��>��c7E�#  ��2�T��=Ze�9Nu��?�4�;\������|>z�$��>y�����|�r?����  �W��c��ZΣ��f���<��n>Y� 7R��η_�ɷ_��w���WO_���'  ��2�T��=bENR��JV�Π	��
�0<����䣏2;;[��vN�;y��M�ݫ� F�-z���n&'�� ���<f���W99>�{  P�*e�S�_�`��9K��mA�Π	��
�0\��Ƴ��0���uO�k����i����T> n��G������36֨{ ���y���/^�%f  ަ�e:I|����S���>��4�;\�����ƽlmm�=��n�"/����q��)  ���������y��G�ͣ�6ro{9��� �O����g�ⳗ���|��봚�g  �P�~ʜG��>U�i�J�N���A���ax--�ΣG;�{
\KG͓�x��~��{
 @�f禲��nv������<x����w2>>V�4 `�i�ٷ{?����79�?�{  0��R�[�`9M��;�}wM�W p��6;;��O�dfz��)p-E�ׯ���{T� �kg||,[�y���l�_����<�ý�Z��{ 0$��̛WG����y�� /����_�����i  ����T9O���� #��y�t~��+pg��pw~y��I��V��,���&��wg. �Ms��|��d��J}t7�>�Ƚ��4��� 5j������|���|��7y�� /����O�  ~�*eʜ'�����)r�*�-!�3hw��;��F���ͭllܭ{
\[UUe��ׯ�Se�s  ����d6��d��Jv��ͣ������L��/ ������{�W�.c�ݼ|���׭��  #�J�*�����*���o��3hw��;���յ<xp�eE��|�r?��uO j�F���������z��e��jV�� \Q��</�������ٷ{��7�y�� �~��  ������v���H;e���!pg��pw=y��I�&'��Z�}���w�i��	 ��4;7����l=X����l_��v��7�@M�:��~�̫�y�� /�����9N��i  @�tS�W�`���H�w�s����@��izj:�?���|�S��;<8Ϋ{����  �u�w <!;  p�U)s�*��?U�9N�����;�&p�+���σ��r��)p�E�ׯ������^ �L� �N�  �*e�t����K�~�S��6�3hw��;�����<x�-�+�t�y�|7�ӳ��  �x�sS��o?\�����Y]������<߿8̋gy�l�2f?�����6  ��T��*���[�v�t��?O�Π	��
�p3,,,���'����{
�Ã�|�r?� p�LL����b��f����m����R��diy��y ����2��'y�� /�d��Qv_����AZM!;  0��tS�W�`���������A����昞�ΣǏ2?/���(�*�o���C�� �3Y�X��ݥ�o,e�������L��b4 �j5�y�� ��[�{}������~�޴�K  �h�R�,IQ�`U)R�8�{~2���A����fi4���������=���y//����S�  ~����l=X������ݼ����0"ڧ�o�7��|v�������Az]O�  n�*Eʜ%�9<x�J?ǩ��;�&p�+��ʹ�����h4�C��΋go���f4 �(��������Z���r����������LL������rt�����9�ޛV^�j���f^�j�ӫ{"  @�\�L7�v`P��/?μwM�W p��kaa!�?��O��ʲ����>LY�T �&�_����R�.������]���[�80�z�~���{�z{���яW�_�8L����   �V�n�x�/08e�S�3����A����f���ΣǏ2??_�*��E^>��q�]�  j411�;���5~��\���T��/�������G�v�O���U�D  �!T��Y���!���O��T|B���A��܁F�������=���q'/��{�  �i��������������.fem1�3�@0�~���I�O��{����/��n�yp�A  x��9OR�=iU�9N5�7��4�;\������j<��������P��*�{��~����  �nrj"�w�vw)�+��<����;�����YW�~�}z��׭���4��{}��f;̓��ie�8e�[D   B�~���2�[ENSf�����@�����|?~���麧�����y�j?��uO `��/������^����Rn�Y��;Y�X��ݥ��-f|�����>=O��I��4��[9:<����޴r�w��   �@���y�\�=�ʜ�H�������@�����xvv�����P�t�y�b/�'�  7[��,-�gu})wV����;��Y�=�6�_�ϭ�sYX��{*p����4O�j�s�l�����i���<8���I..��i   ~�*Uʜ%��*)r���!pg��pw��ظ���{IuO��t�j����t�.  P�����/μ��<�啷��ۋ��Y�������Y]�Ą�����pq�}z���i��o��7�i���}z���v�S  x�)s��ӵ��L?ǩ>���;�&p�+��dii);;;����{
��������W�� �и�4�[��r{y>K��!�|n-�eye!��f����*|��M�0���z9n��������P�u����۟[�v���9i�y�  p�T�L���R�8e���)pg��pw��LMM���Ǚ���{
�~���f��4S� �295����,�Y��;�_������K�w�|g>�3�?�s���(>�^���v7��nڧ�?�h^^Z���;:<M��41  �OU)�MO�>�"��'F|XwM�W p�b�������R�j�罼~u���I�S  �c�_��⭷?n-�f�����?�8��煙�Ϳ���D�$g�^:��e�~��㳜�:o>>�����;=>�q��ӓ�t��   �vU�������L/ENk�w�4�;\��x��k�;cccuO��vr���{9?��>  ��.�OMM\��_W����_�����LOO�ϵ򿮩���/z�\\��gNZg)
1   N��e�.�>�*E����c���A��܁w577�Ǐgzz��)0������\\��  #m||,�sS?��?�zjz2������g&377������Nev�_�������xf�2=3��	o�eUU����W���}z��ſ����Ӿ���E:�^�E��z9�t��޹��~���  ��P%��M�^�S��J?ǩRԶ@�Π	��
��o1>>��w��|��)0�ʲ����>LY��  �E�����djz"���_���Կ~����D��'399�4���f�.�'����ߛ������ߛ��J�����x���~#efv2��c���T��?�^��c�iwSUI�/r~~�$9?�,������R�e:��߄�_������>OQTo#��������s��׽��E}�@  �z�)s^k\
�\ENS����;�&p�+�����z<���wxz�~^�����q�S  �!1=3������m������cl�?�࿫n����߿���%���m���o���7�    ~�*��9��� V��9�{������܁�kn~>O?���͸��n��Ջ��O��      �e��j���\U.R��Z��F�Π��=  n�N���O�����ix��g��'�����LO{�      N�*e:�v�6U�i_��>�; | �~?_}�U^�|��Tླྀ�4�?�y'[��3>�S[      ����O�v�uOn�*ENS��{|0*  ��^��>_}�U.�����Hh4Y[��?�y'+�Ki4uO      F@�nʜ%n&5*�I�7�� jprr����999�{
���ɉ�x7���an//�=      RU��9K�^�S���y�t��� jr��端��������gff*;����?>���\�s      �!R�H��k�@�\�L��P�; Ԩ���z�*_~�uz^��4??�����'ogvn��9      �5W��2�T��5�R�H�G#n,�; \''�y��g99>�{
���[s��Ӈ�y|/�ӓu�      ��*E:�ҫ{@�~L:M���!P�; \��E���˼|�*U�����^^������frr��9      �5P��2�$E�S��`������uπZ	�a�����������W_�w�Ux��FVV���_���j��}:      7U�nʜ�R���h�=�w*s���$@��d�������I�~�i���#il���w��_e}�N�     ���J�2�T"R��r�2��g�� p�k����믿���/RU�-�011�ͭ�|��G��r��9      ��U�L;U��� ��J�"mϓ�Kw ��vw��/��y�[�YSSy���?|�0�su�      �L7e�	)p�T)r�*e�C����h�O�����U�iss����y��vf��      �e�tR�W���Px���; �~�����|�ݳ�w�� -ޚ�'�>���{����{      �U�H'��P����|�a�� ��98�K�}�G��dvv��90�n//f��B����A..�uO      ��JR��j;pmU��Y�3�Zr� ����y���ivww�#��hdeu)���Q�m�f|ܧ�      p�)���V�"E�uπkK� C�(�<�<�|�M�£�`�����q'���Q��.gl�Q�$      �g�u��{
��P��I�Tu�kK� C��l�Ϟ��Ի:�C�����Z���<����;      \Uʜ�L7��V�~NSy�"�; ��^��/��"/_�JUy����x6�V��??����4Bw      �C�~�tR�_��_T��c\�� FDUUy���|�ŗ9�v�7���D���ӿ<����      >�2ݔ9s���>e�W�
w 1��i>�4��Q�S�F������w��?����-�;      T�"�TbQ`T��Y�3`h�`E�o��G���)K�R�izz2v6�ɟ
�     ` ��S����{
���R�H;U�C`��`����gOszک{
�833S?��      #�J���+�RQ`T)r���,x'w q���|�������SU>Y�mff*;��	�     �w��䋺� \�۸��&�]	����*�^��_|��n��9p#��N�     �7(�M�N\m�I�vJoʁ�D� 7H�}�ϟ~���������C������|�s      �ڪR�H'Ur�K�����=��� n��(��~�o��6EQ�=n����<�h+r?�su�     �k�J��j{Q��wR��"guπ�6Q�  ���a��vvvv���P����f����>=˫��i�z�     �MV��y�����޾9�]�z.����u��_�������9p��/���O����ۙ���{      |pU���ہ�T�L��T�����; ���7?^s���B�o��[�::ׇ͛���      U%��M�^�S ~�*ENR��{�����k�_S�e���׺g ���x�ݻ����uO.�O�������t�      �]��2n/��9I���g|0YL#�u�`���=  �>ʲ�˗/��W_����x��f�����'�ski��9      ��T�̙�jE�7*n�A� ����V�~�Y���\�_��㏶�O���b�s      �w(S��2�$U�c ~�2�ˀ�I� �WEQ���.�|�M��~�s�Kss��y|/���a��J�Ѩ{      \Y�^�t\m��ۧPt�#I� ��f���>{�V��)�O��N��Ά�     ��P�J�3Wہ�P��"m�`@� ������믿�?��<eY�=�����<���������Bw      ��*��i����ïJ�"����00w ����w�����>m�=�����l�_ϧy�����     P������v`4T)r�*D� 	��wr�=�_~�W��OU�\7SSBw      j��j{��v`����^�=F^���4�5eY�o��{��3;;��������=���"�{G�{�LQx9      �V�L/Uzux���S�[��ka"�id���0����쬓�?�W/]s��jbb<�V���q�m�fbb��I      ��*E�t����)s&n�h�� �p��*߿~�V�(;�evv��I�1>>��w������Vv_����      ���$U��v`$���Y�3�Fq� x/:g�|��Ӽy��;\ccc����Χy���LMy�+      �]�"e��v`$U�H�v�3��i��P���,��m��u� ��������t�S�_QUU��'�}����ǩ     p5����J?ENREf�sYL#�u�`�	��
� �nll<������ݺ� W�>=˛ׇ9ny�9      ��H��T)�0UZ�F    IDAT�9�q��3hu  FSYy��E�Z���ܧ�������<�h+�N7���4ORy?,      ?Q��2�����r���2V�  `��OO���ϲ��W������`g#��NVV�26֨{      5�R�H[�������!p�5�~�$#���,�տ�=`�-,,�����LO�=x�~���������"     �f�.����0p��s5YL#�u�`�	��
� ����x�ݻ��w��h�
ä,�췲��0�^��9      X�"eΓ�uO�"�ˏy��;�6Q�  �f)�"/_��Q����33�;���F��ogm�v�[�|�j?g�\     5U�*�T��7D�sq;\#.����0����k��������uO     �=�R��y*Wہ�L/EN�1T\pg�\p j��5�������Ch~a6�?�J����n3�ÓT�C     0t\mn�*)��p��W��;���5�{�^�mn��C�۽��n3�����      àJ�2牫���TIF���O��T��w�;�&p�+�|8s�sy�����ٺ� �C�_d�(��G�����      �_U)�s��q��q�7��wM�W p���F�ݻ����aؕe���V�w��v/�     ���)ҍ����S��cq�� pg�&�  �sUU�իWi6�y�p'��suO~���F��ogm�v�[���6srܩ{     �V�L7U'n�*}����� ����Y>��iVW׳};�c���0��4�[K��t�9�;J��8e�R      J�~�t���U��I�u~E��~EY����_�p�MMM��Ç�uk��)�{��9�oe�(���      ��*U������ 7W�Ӕ��=c$Ld1�L�=�&p�+�\��w����LLx�����::��f:���      ��*��9O"n�"���=cd�4e 0T��ôOO������;u�ރF���ˋ������Y�v��::M彸      �C�2]Wہ�̙���� :���|�ݷi6����~�����'���_�M�{���V��Reݳ      �J�^���j;pӕ9O���g ���Cg�הe������ ����������z�S�(�2G͓�i�{ޫ{     ��V���R\�=�vez)s�>0��42Y�F�� �P+�"ϟ?O�y��fff��I�{4>>��ե��.�ut��ݣ��t�     p�TI�tS�� �$�r!n�!�;\�� á���ݍ���H�Ѩ{0 gg����yx���r     ���^m?OR�=�Z�r�"�����;�&p�+�����<xp?���P�_�`���ݣ\\��     ��U)�s��'��S�D�>`wM�W pN++k������D�S���*����i��>�{     ��U�_^m�~��Jq�{�Š	�4� 0��r�jf���ܹ�\�`@�Fn//���bNO:��k�ut��{y    ��S�L7U<�৪��v!w `�]�����o��+<���tݓ�ZX����\..�9<8���Qz=_�     �_�^���j;��U�v1��:k��,��m��u� �w���F66��h�=�@N�;��m�ծ{
     �;��O��p࿪�ω'[|`YL#�u�`��� �eY�ի�9j��Ç����{�,ޚ�⭹t�9�o�p��~��{     ���R��*��� \S?\n�èq���w�Ѵ����������=��ʲJ��8�{G9�t�     ���S�<���)r�2uϸ�\pg�\p n���ݴ�������ʝ�� ��X#+�KYY]J�����Q���)K_      �U�L��T�4Z�_R�T�#�w��F���b>|���麧 5(�2G͓�i�{�1�     ��U%��M�����ˊ�S�Ӻ��;�&p�+��c�FV�ֳ�������� 599��`����i*/�     ���O���~]����L�$pg�&�  p]�U���7i�Zyp�~n-ݪ{P��[sY�5���~�[��=J��1�     ��U�L����v ~M)n��w��n���۹��A����n����::��~+'ǝ��      #�J/ezq��jʜ��Y�3��;��; ���j���N�������i4uOj�h4r{y1��s~����Q�[)K_p     �M�"U�S��{
��(s.n��w������Ç3??_��(�2��9�o���[�     �ګR��*��� ��q�'m_7.�3hw��; ?XYY���V&&<x���y����q�µ     ��U��y���(�M����א��A��������lnngmm%�F��9�5Q�U�[�9�o���     �H��$� ��*�9�_Sw��Q �wTE�?�g�������/��=	��������ˋ9?����8�����E��     ��J�^���0����.��M�;\�� �����lmmer�{�WUUZG�9<8��q'��_     0ªT)R�<�e�&U../��8z���Π��  ~����5�������4��'�D���^?��������=     x���&�dW�ߪJ_�$q���w �jvn>�����|�S�k�专��VZG���    �P�R��*��� ��q���}H��Π�� ��u���ϳ������LN�d�O���xk.��p��n���Y     �;��K�^"��]���Ϲ�W��; ����x677����F�Q���;=y{����;     \gU���K���) CO�>�\pg��pw ~�ٙ�l��[����(s�<���Q�:ݺ�      ��T��MOe�JrSN�U)R�X�>�����@���������ۙ���{
0$:�n��r�<IQ�u�    ��J���q��}�7�;�&p�+�𾌍�����llldll��9�������qڧgu�    ��Jqy���{
��x����#_�J�Π	��
� �o��S�����ʝ�� C���yx���V�]�@    ��(S��*��� �q�h�3hw��; ���x+������L�S�!��t�<h�yx�~��     ������EY��$nwM�W p`�VVֲ�������� C����wrxp���i*/�     ��U��y�� }��4 �5pp��V��{��emm-�F��I�i4��4�[K������N��w��N��i     0ʔ9OOKq;�\p�+p��iff&��?ȭ[�uO���y/��i��_�     �V����K���� �,q�hr��A��������ܿ����麧 C�������yx���I���@     n�*U.RƓPI�>�����@�@]�����es�^�������(�::M��8'ǝ��     �U��2�I$S �$nmwm��  �oUUfw�M���ٸ�����4��gCl||,wVn��ʭ�z�4�s��J���     ��"ez�ү{������p.�p]���f{{;KK������Y�s�<IQ�B     ��J�*�ҫ{
�� n�\pg��pw ��۷�������麧 #�,���Nsx����Y*/    JU�\�L��! 7�����3hu  ��5�j�������{�{0"��Y����;������i��S�4     ��*�˰]`	�ہ�I� 0������dss3���i4u�F���x��ʝ�[���9j��yx���k7     \GE�tS��{��"n޷��=o~MY����_� �hvf&�6���|��)�����i���8��^�s     ��T��M���� �8���i"�id���0�;\���a��x+��ۙ���{
p����^v?8N��     |HU��.�v	��&n������@��0Z^^���V���� >���Y��'9j���_�     FX�^�\$�J�ZT�_��ԛH�ΠM�=  ��h6�je}}=�{0��f3�0���t��9<8�Q�$E�     �U�)Ӎ��>�v`�\p�+p��a791��{Y[[K�Ѩ{p��e�ӓ��e������     �E��R�D�$n'q�������3��������uOn��(�::�Q�$'ǝT^�    ��˰���! 7^��9�#pg��pw Fͭ[���}?��3uOn�~��Q�$�Ó�O��    ��S�$l�7�M��O	�4�;\���Q�������LMM�=��z�~��'9j���>�{     ��R�"ez�\ez)���#�;�&p�+�0������fk�^&&&��p�^?����Nszr��KV    ��J?e�Iʺ� p�m�~*m���4�;\����`||<���������� ��/r�j�y����    `DU).����) �D����v�wwM�W p�&���ν{YYYI�Ѩ{@�;    �(�R�J7U�uO�g����;�&p�+�p������V��o�=��E��ѩ�    `h�)s�*��� �_�9O�N�3������@��M�����������=�?�e�ӓN��'9j��,��    ������E�&0��$n�*����@� ɝ;w������麧 �WeY�u���i�[�bw    �k�J����E�p}�9K���g0��D�  ���i6�YYY˽�{����$p���5r{y1����{��4EQ�=    �F�һ�!l�ΊtR�� I�  ���������Ã���gc�n�������wg�mj��?� 'p%׊�諨�������{��Z�dY"%�������dK65���y" !H����I o�	�'�f#{����SUUƣY.��y�n����{<    �G��:eI, ��L6߳�ƿ���	�,�����= �;�v'/^��gώ�l6��o]��W����     ?�eؾL��W����x�}n���4ҩ{1�;܀� �Z���O��/9::J�Ѩ{��N�8���8���     ߪJ�*�T�v�������s��pw ��^��?�K����-�\�Orq>�x4K��2    �ߪRn��uݣ pcU����7�s��pw �:[�A^��/98د{�o�^���8����8EQ�=    �=S��*U�u�U�$O����&nw������&p��������?��loo�=
�7+�*��4�ƹ8�d���    x��T���<@U��v~ �;�M�7 p�ﳷ������ڪ{��6�/���(�ƙMu�    pG��Y&YFl��T)6q�+����6�;܀� ~��p?���?2����X.�]Lr�a���4���    ��S��j�{�!��	ܹm�  ��8?����988�?��/��zu��]��v���9:�(ʌ.&�8�ދ��    �C&lx��7q�����!p �ν�.>����q^��<}�;��Z���f�`7UUe:����Q�?��\��    ��.����< �*��ہ����\?�NY�����{ x���V�����鴝	<N��"�ƹ8g6]�=    �gUYn>�D ]�e�L|O�V���F:u��#&p����k6[999ɋ��j���֬�Eƣi.�'�8�d�.�	    xҪT)Rf����(����T�έ�s��pw �;�V+ϟ?��ɉ�x����t2����vw    ��	��2���=�����&p����k�[99�O�����?�S�T    ~�*�TY��+L<&E&���v	ܹmw��; ԧ�n���D�<9UUe6[ft1���$��M    �����>��� �O�q�,��'B��m����~�vg���X�<I��    ߪ�z=����T��}U� <!wn��n@� �G�����/rr�,�f��q ja�;    p6�<ve��ʺ�Axb��6�;܀� ��;��lw    >&lx���)2J���@��m������ݟ���D���   �)�<U�M���=��s��pw ��:�N^��"ώ���h�=���Z�3�2��d<�f�t�J    xl.��Eb�/��We�"cq;��s��pw x8lt�k��*��4��iF��?   ��<-U�)2I�'��s��pw xx��vNNNrrr�V�U�8 �RUU�͖���ǣY*/    ��We�2����2���H۹��6�;܀� �����&t��௔e��x���r��l��{$    �Z�*E�,S	���2���=\�s��pw x�lt�z��:���z��r��{$   �N��v��N�����N��V��f��V��f��V��V��F���?���E��(S�eʲJQY���V�W�V�˯��Ey��� ��2l/�H���SSd�9��!p�	��� �x�Z�<�<�NN��|��|��h���4��T   ��4�t{��������6�w{��ۭ��o�j��b��b��b��|��l��j�$o�~���<YU��SfU� �'wn��n@� �O�����I�����n�=��SUU���f��,��,��   ��^���V?��^�^z�n��v���X.יM�N��g�Nf)K�{��bc; e���/����6�;܀� �V��gϞ���$��'_ ߪ,�LƳ�.&���f>s�L  �Ǯ��fk���V����j�=֭��*��<��ԉ��-�Re�*�T�=੪R��8U��G�/�s��pw x��F���O/������+�������$���  �!k4����d{g��ݭ�ۭ�ǪMYV��9�0���$��͚���OS��a]���UYo�vW��~�s��pw x:.C��<�S}�;���q�~yi��Mw   ��Uо��}�?���?�d<˻��|x?JQ������L�e"lx�,Sd�d'�;�M�7 p����h��� /^��`0�{�G�(�LƳ�Gӌǳ̦�;  �j�[�ބ��;�?mc�t�i6���ZeY���8��]dt1�\��*e������$)�H�������&p����6��O?e{{��Q ���2�lx  �%�N;;��탁�޶�j���9;=�|��{�^(Sf%l�ef)2�{�*wn��n@� $���N~z�S�ý�Gx�ʲ�l:�x��}2��,��  pS�^���~���t��7�����	��U)S]ol������!yx��6�;܀� ����V^��)�u��dTU��l���D�  ��F#�~7���l�����n�]�X|�j�λ�������r]�8�-��eU��S:F�@	ܹmw��; �9�� /^<���a��F�� <)UUe:�g����  �S�h4�u�o6��Zͺ��+TU���Fy����g6v�cS�؄�Nd�Ϫ�)2J���Q��	ܹmw��; �W��^N�����q�Mo$��*x�g�N晌gY��0  <�f#ۛ�}ww+��~�M���4�=�d<�{�T�R��2,�U�)2N���Q�ܹmw��; p�v;'''y��Y�m����|����'���x  �����=����n� ��]�O����� UYm6����*����d��O��m������l����qNNN��v����(�c��x��d����  P�F���V/���렽ӱ<�);;=ϯ/O]��*UV)�J�� ��2�J�y4��6�;܀� ��F#���y��E�~�� �UUe6[^���,���  �G��ig�*f��g��O�i;;�Z�����4g��u��I�2�TY%2E n��4e�u�?����&p�� �k8�ŋ��٩{ ��j��l��x<ۄ��T^:  �Q��H����V�z;{����x4�?����^(7�ڗ�v n�J�I�,�~8�;�M�7 p ~����<�"��^ݣ peYe6���D<  �%�v+[��lm���3����vv�[Q��埿���Qݣ�U|�� n�?H�    IDAT�:�Tq�"�����&p�� ?Z�����I���l�= _a�Zg�	���Yf�E�#  5��:כ�mg綽;��/��-e�-~�U֩�L� �:U��JY�(pk��6�;܀� �-�N''''9~v�v�]�8 |��(/��O�N涼 �#�鴯��oo�3��ղ���5�.�_��2˥M�p;�T)Re!J��TY��8Ud�<nwn��n@� ܶf���ã<�<�~��q �N��:��B�  T��L���V/��~�w���q���^���x��xV�(��T���|��6e)3��$ܹmw��; p���a~��loo�=
 ?�b��d<�l:�t��l:wYy  ��Fz�n��/C���~��n�c�_*�*���������Q���Rf�*�D��w(3K' �tܹmw��; P��ݝ<�S�ý�G�TUu�O'���b�L�  �5�샭^���i4u�_�����߿���Eݣ�T��ll��S��$e�uwJ��mk�=   �y��8����֠�gϟ���ț� �H�Ѹ���O�]�W�U��Y��E��yf�yo� ���v��ھ��~���lz}�ǡ�h����^$��n�J�"U��R�= �@�2EƩ��{�G�w��������ٳgy��Y�m�<�u���>�DV^, �?�t�l�2غ�ٷ��i�[u�w���Z�_T��*eVIʺ��������-<M6�s��pw �>i6�9<<������u�@����6��� x:z�N[��z��܊�yʪ���ǫ\�O��*�f[�*�4���2e&�_x���6�;܀� ��vvv���Ow���6�S�Z�3�.2�-��/3�.2�-�  ���f���~��lf�/)�*�����d^�(P�*e�,R������<E�u���s��pw �999���Q�; ����l:��ݧ�����r  �P��Hн��>�2����Z��j������r��{�c�&l_����p;�LR�bH��>�;܀� x(��V��O���Y�O&�����X�2�̯���t���  w��h���fk�2b������L������Nn�ɸ��W�R�=
��Uŵ��Z�"��N��kwn��n@� <4�f3��999�`�U�8 < ���z��l:�|��j��z  �_��J��`��`�����
ܢ7��ϫ_��=ܢ2eV���e�	 ��J�"#'R�ܹm�   ~��,szz��ӳ������Y���6/ �E�~7�~7�����V�̦��f����<�Ū�) �Ϯ�����lm��t��xK����G�\�O�~�*�fc����}UV)2N�d*�;g�;܀� �c������$GGGi�Zu��U������2~_̗)
�k  ��N�}��}��`�Kе���j������k<�Ga{Q�0 <e�)3������m����Ǥ�j��� 'ϟg���= ��j��|��|��|��|��l:OYz�	 �!��ʾ���lg�e�ճ��ӷ��?��=|�*UV�'j pW���̢�A�^�sۼ�  OLQ9==���i��aNN�eooX�X <p�N;�N;�{[��UU��bu��g��f�,�Tv.  �;�^'���V�n[��zެ�����~޿e2��=
|�"eV��N���N�Yg�9P'�;  <a���9??Ϡ����I����j���G��h�����~rUU������bUӤ  OK��No�s��A{/�f��р[����$�����ǀ�Q�J�*�T)��'��:EƮpO4���uY�wʲ̿�k�c  ܺV������<�A�_�8 <1���>���  |�N���������d��K���vxj��?^��ø�1�O�TIV��P�2˔�l�K�M���F\���c�;  p�(�������4����<;���0��p���(ʏ��Ef�����F7 �F��n������V�~�Fv��O�8���$��w�E�M� u*3K�Y�c �w  ��?|������9~�,�G�i�<� ��Z�l���3����(3�/��/�o�U�h xt�F��N��~7�A7����k�~7���|x?�{��*U�TY�����[�"��Y�= ��N  ��|>�/?��W/_���0Ϟ�d0��o�[�j5�����v������r��ߗ��u �Z�k� �f��F���M쿇�����>�N��ԢJ��z[���_�2EFN����  ���e��oO���i���rr�<���\��i4��:��:�n�kUUe�Xe>[\o{��Y̗)Ko� w��h��m�����|������=�Hm�2��e6]�=
OB��H�U�8�����*EƩ�tp�5����5��)�2�v��u� p�t:�<{�,G���v��������|����v��F< �m:��u�~����9�	�@N�~�/�|S�<j�f[��V\ �2���H��hg7�h�=6�  �l�Z�իW���_����g'��٩{, �&�n;�n;�{[��_�U��e������|��r��ڛ� �ԵZ��D엷ͦ��_�v��緩���+Rf�*�D6��S��4e\�����UI��p�����w�����lmr��Y��l�� �[����V/[[�?�ZQ�Y,VY.���U�˫۵h �V��N�s����Q��n{�<�v+�;��GӺG��|ƻN��m� �[U���+u<$w =q;�ݚNg���3/�%999�`���� �V�������,�����*�_,�Y.V)�����/i����:�����N����� ���p[��w*Sfe[; �^��&n�Z,�C#p  nEQ�9==���Y�wvr��8�i4�z���h4.7�~!�[��,��>��/���V��� ��]ma�:>_��n;�^��U������/o���J�r���\ �2����r2��$p  n�d<�����?���a�??I�߯{, �U��J��J��|L�� ��-� ����ne�.���2
���n�- C�"ӔY�= �A�  ܙ�(rz�6��o����gϞe8ܷ% ��&�ߗ�uV�է���(~��M�ǧ�h��i����m_���������8��=��m� <LU�;~<w  ��\\���stt��g����� ����[�?vVU����jUd�Xf�*����b���k �O��F:�v����n�����n�-`�A[w��j[{�Ub[; L��&nwx�  @�V�u^��-���&��0��G�ID �.7�^F�[_�����r��j���]�_U�O�c����W!{��I�լ{L�'�K�x�lk��+�H���d- �;  p/TU�>�Ç�v;9>~����tmu�[�j53�2|�X�Z�?	ޯoW묖�ׅ��x�ݹڸ�N�j��&f�tZ���#�n������ڗ���J�i�,��L�  �;��*�^�ʫW�����g�G��?C ������S�u�Z���^�6!�f3|Q�40�C�j5��N�}��u���|���tZu�@-lk��R���1���  ����"���t:����(G�G���� w��j��������ʲ�s�������} ܾf��`��i������N��{�+2=�Q�:�m� <UV���q��  �j�ʯ�_��ׯ����gώ3�- ��h6��:��:�����\�R��,����׫����U��jo���/��v����ͦ�R O]��r��#W����G��<e��v�GN�  <8���H�����a���ӷ� �f�q�~�o[eV�u�u��(?�᯾.�2��:���vJ�Aj���t;�+f4/��w�i�~�֯��V�Y�� < �F<Veʬ6Q{Y�0 �U)2I�e݃ p�  ���Z����oy�����n���Y���l�� ���g�Ə�����"��v��}#��(� ���h4�n��l5/���ԯ���u���� ���m�v��S�H����"p  ��h��h��[����8[[�� xJ���z�=���O������(�O6ŗE��(R�6��c��P������Z�����  ��2j_��*��! <Ne�)3I�X�� �G�(ʼ}{��oO��5���q���jy� |�F��N��N��~���*EQ^��W��_�w�_��y��F�::o���1���v�2Lo}�7[��?o6� x��TYm�v[lx���RdV� �@�  <Z��,���y��e���9>~��ݝ$b ��\mvn�[7������(?��q_eʲ��_��[�>/����~_
ӛ�FZ��澫����f���fS�����ʇ���֞���	(��xs��)�  �^Y�y��}޽{�^���������= ��|���c������?�>�ʫh���_����S��$5��F�q�7�47�Wq���W��l6>��f����Ga��� ��"�*U�Uʬ�������:EƩ� �4�;  �,��z�k^��5�{�9>>���A�fݣ �p���������8�����eQ������~l�{p��}WQ���+�#����|\u�ث�����R�u�s�U,���z[�Ǜ˯B�?���ǟ���]��q|�h\�z룈 �ߜ�xm~
N���� <9e�)3u� �  ��5�et1���sxx������c$ �߻ڦ}��q��f��{\����k}�'�F��l6�h��������q��Ux pSE�m?�p�����=�> ��*E&)��{ �	�;  ���E޼9͛7���{9<<���az�^ݣ �>����z ���s'�q��T�fS{' �4U)Rd�X�'�   ��y��U^�z������� Ϳٲ	    ���N�&h�� ����"e���� �ww  �/����b�_~�99::���vu    ߡ*�w�J�Q������J�i�,��{J�  �7��"oߞ����������(�n���    ૭VE�#<	U��z[�s H.��"c�F ���  �+�狼z�k~��uv�vsxx����4���G   �Y��u��hUI.���f[; p��2E&�6GL ��;  �7��*��8��ϭf���spp���a�F��   ���?X�*�fS�*�����̼�1 x �   ߩ(ʜ����ٻt��������8��Vݣ   �����c\F�W��˺��{�J�"cW6��  ~��r�7o��͛��rpx�ã�t;ݺG   �$�jU�=U�J�J�u�� �W��6q��� �u�   �d:�e��e^�z������� �f���    x��ka�׸L��mk �N�i����J�  p˪����E...���?��� GG����MҨ{<    ���rU�B�⣨��Y ��*eʌ7W;�o#p  �CEQ���,��g�v������0;;��   p�V�u���{�{�H���.j��Se�"�T�� |'�; �3U� O�r�̛7o����������0�^���    x��e�#�Ce��Sf�D� ߢ�,ef�v ~�; �3�v��i>_�ի_��կ�����8��v�u�   �#2�-��^��,���w�Rn�����GD�  p�L��L�?��/�d{{;�G�9<8H��)    �g���*U�TY�� ���L����1 �q�   �TUU�������_����ã����h�=    �S��~�ۭ7Q{q} �}�LSf^� <Rw  ��,˜�_���"?����~����F�Q�x    < UUe1_�=���Ծ�lj���R��lmw5 n��  ��Y��������,�v+��0������K"v   ��y����U����}Q; �xU����q��%p  x���"gg�rv�.�n'��988��Ύ�   �O�FӺG��I�)�NR�= <RU��Rf^�  <w  �Gb�\�͛7y��M��nspp��`��   ]<���J���.j��V�H���2 �w  �Gh�X��__��__g0���`?�����   <=��:���1��� �^�E�LS��{ ��;  �#7��3��ΫW�3��p��{���   ����u���D� P�*E&)��{ �(�;  �2���r:�˗�n6�d���fw   �G�����nD� ���N�q*�a j$p  x�.7���W�~M���p8���Avv�#v   x<ƣi�E�c|�� �2�����{ �<�; <rU$� ���b�7o��͛7��z988���~����H   ���}�#|�e�^���vUʔo�� P?�; <r�D ��b���ׯ����t����spph�;   �4��sq>�{�$6��}Te�"�T��p��  ���r�7o��͛��u;���   �W����o�R����T�v �G���̼�A �O�   ��b������V����goo�FC�   pߜ��g2����{��=Y� �P�"EƩR�=
 |��  ���^9;;���Y��V���spp���=�;   �=�\��t{�U�^e�����*3O���� ���   |������YNO��j5��p���)v   �seY���W)��V��˘}�2ED� pߕ)2I�U݃ ���  ��Ey�ٽ�jf8����A�{{i6=   ����L'�[���ͦ�U*Q; <U�)2M��=� ~u   ��(ʼ{�!��}H����p7���i�ZIlw   ��^��6��.~��X��z�Q��? �}U��R�6N|��#p  �֕e������y�Fvv������p�^��;   ��{��ۼ���w�9�!{!j���:E&�� <Hw   �TUU]�3�������������[[[�   |�����?����U��6�'� �ce�)3K���Q ���  ��l6�l�k^��5�^7������gk{7͆�   �,������l����w��]mh_	� ��R��8e�u� �E�  ���X,��oo��oo�n�2�eo8��p�f�SX   ��}x?����[��׫T)Re�	�E� �X�Y���Ik <
�    ����������O�����n��a�ýt;�$��   O�|��˟�dt1����TYo>�[� �kU�LS��� ���  �{�,˜8����$���V��{��?�`0��   x
��"�_����<U���[�/���������*E&��xd�   <8��4��4�^�N�����0�������h�=   ��X�rq>���8���a{�2E��fK���w �1�Rf�2sG} %�;   �r����iNOO�l6���������t;���   <$eYe2���|���,��/=�zK���Vy <U����/��  ��  �G�,�\�_���"I������^�ý��i��  �{h>_ft1��-�A�e�v� OI�y��R9��GN�  ��5O2O����t��ݻ�݇{ôZ�   ����>Ms�a��|��GV��}�*Eli���J�2㔶��Dx7  �'a�Z��ٻ�;{�F����������lmm�=   ��-��.&]L3���(>���2d���~�9 �Y����v ��;   ONUU�Mg�Mgy���t;����7��po�vw   �UU��d���IF�̦�/=�:f���-� ��2E�)�+� ���{   ���j�������m��6��������Q��   ��^���8����ؖv ���Yn���g	 x�� ���"�a���>�l:ͫW�6���2�������   �FUU�͖]Lrq>�d<��#7ڋ$k� ��fk���� O�w��;!nࡺ���.gg��h4������0{{���ڮ{<   ��]mi]\nj_�֟}�-� �ר�J���  w   ����2�3���e6�݇��������   ��|��}<�f<�����=r��}�	��i �M�� �w   �F����rvv�F���������ekk+�a   �b����>���(����ݖv ��UYo���9 >&p  �����Ǔ�Ǔ�|�*�n'{�a��v�������   po�V�G��.&]L�Z�����:f��>�� ��T)3O���& �3��   .��    IDAT�`�\���iNߞ��h�?�g���www�h4�   ����2�2]nh�M_xd��:j_E� |/[���	�  ��UU��t��t�ׯߤ�lf{g;{�{������V�F�c  ���X�2Ms�a��h���R�^l6��S��� �1lm���  �+�2��QF��|��z����fwo'��{�;u�   �j����~1���$�������د��"�v �G�� ���   j�X,�X,rzz�F�������nvw�����F��  ௕eu���]L2�.>��*U>�Ҟ�w:' ��� �B�   �HUU�Mg�Mgy��M��f�w������0[[[I�u�	   ��t���b��h��h���\:Vmb�b�5��T ��U)Rdlk; |�;   �ceYft1��b��/_��negw'������M�7���   <��*��4��iƣi���cU����� ��}k��� �-�   ����E>�?χ��I�N����������^��;   ��j��d<��b���$������оN�2� 5�� ~�;   <`�������fgw'{{{���K�Վ�  ����}<�f�X}�WA�e� P7[����  �#�X,�X����4���������Nvvv�j���   ���:��e�>��"h/7�ً�FT� p?TY����v ���   �HUU��d��d����2x�����흝��7�  �n|��}2�g>[|�q��O�b��M� �=T}�� ����   ODUU�N�N�ɛ�4��������v����  �r�OƳ�ǳ̦��/7����=)�rL ��bk; �.�;   <QUUe6�e6�%���}7;;��w   ��z]d:�g<�et1�b����u*A; � �� wA�   $�c��&�F#[�[������Nvvv�   |b�.2M3�2M��/��ȫ�E��cC; ��TYm���9 n��   ����2O2Or�����lgg�r�{�ݑ�  <!�u��x��h��h�����/���u�.h �*E�)�{ �M�   ����߼9M��{����{{��v���  ��X�֙�g�Q�x�����b�Ww9& ���� �!p   ��|��|�.gg�$�N;;;���fgg'�~?�w  �����,�߃��4���s��D^�� x����� 5�   ?�j�����y��<������Nvwv��l�j�  �$)�2��<�M�>��R���/��*�\F�e� �cUf�2S[��Fw   ���1xo6�l�������l���jŖw  �۷Z�3�.>
�穪?��U�|�����Y �Z�2e&)��{ x��   ��)�2��$��$�oi4���������n�w����"x  �~��*�M�>��3�-���˼�2b���K�J�'��<ef�� ��	� >��� �BUU����9==K�t��l�lggg'�;���i6Z�?{w��ؙnkt�#�}����.W�R����`����l$-@cD(��x��Q�ˏ�&�  ��Z�:~����_/��\g~ ��j�yJM?�) �w �o��tڶK����;I2���{���!����������r�� �mJ�O�<=.+�|kq��ה1ܲJ
 ��q��h� ���   �j��<}z�ӧ����o�d���������[��I� �;Uk���f�t��c����ץ&�SS�1j� |��W��& �Vw   ���M��&����$����n��~;E�e�\��e  nQ��9����K����
��� |��!��|��� �u�   7���O�>�ӧO���u�{|�o���><d>[Lx%  ��J�9�O�짘����z�i�}�F��  ?��W��ԧ  �A�   ܥ��������H��f�l�����{���c��Xy  �S��y�t�ӧC��&��cj�����u�!c ��2���S � �;   �!�Zs�r���o�d�����1���[v���wY.W�w  �UC��阧�ø�~L���^�%��b���5  ?��I�~�M8 �-�   �0��������<�ݮO��������n��l!z  �V���Ⱦ����~]j��칬���  ^K͐!O��> �Iw   ���6�c���G�d6�e�]g���a����Cv������  >���s�7��鐧O��ǔ�y�.f xO5%ǔ���'p   ���M������l6���)z�lD�  p���?-����쟎����|��$e�s >��n\m�� ��   ��R�:d�tH�{�S���{�����?>f��d�YD�  p;���xx��ޤ��/^U�x��c� ��*�OI;�! �+�   ��RJ�>=���S��M�,�<�y�=�a���n7F��i�  �����&�����t�����#  S*9����	�   ��0�|��>���O���</��v�S������Cf3�;  ��/c������V�>$)���]� pMj�٧���r ���   ���K��o��g�Y��Mv�]v�y�m��e>_f6�  p�^����c�c���>{�i���[f �~5C�9�l�;'p   �X�5��1��1��_I���:��.ۇ�����CV�U"{ �$����c���a�~\f��C��*�y���ˢ  nEI���H�B�   p�N�{�áI�����z�����vc����f�Y��  �{�㡹��MJy�����O��� nU͐�}J�~1 p7�    7�m��m������s���Mv��<��{��n��|k�  ܢa(9��"�)loS��P����\�v!; �}�)9���= |@w   �wZ{?�p8&�?��o6�S��pZ{x�Y{ જ�˶9�������z��^s^g�� p�j�ُ?� |Dw   �;�4m�������b1�f����!ۇ]v�lvY.W�� xS]��xh��s<49�4��W���y��9f ��Ք��S�N}
 01�;   �2%��}�O�$�_�_,��>���޷��͗�w  ~�0�4MwZe?����&]�_^s
ٿ\e��	 �Q�Sr� ��   �C�ӧOy�����l6�z�����o����&�-��  \�u���)h?4i[!;  ߧ�ː��� �g�    |S�5MӦi��;��<?�Ͳ٬.K��w ��VkM���%�Cs	�ۦK���M!;  ?�d�!%�ԇ  WH�   ��,u����U6�mv���v��|)| �r琽9>��c����R��U�Bv  ~A�1%���$ ���    ����������/߷�����f��|!| xo�Xl�Z<����E�o��%! �j�y�� �?�   �^.����{����l��l6�l���}�^'�w �_R��!��e�琽�������� ��S2䐒f�C �!p   `2mۦm�$�����b��v����o���כu2[H� ^������ض����S�^ǵ�rYe ��TrL�a|�	 �}�    \�a(�?�����j���C6�u6�mN��f��l6��w ��ZӶ�g+��c���0������5v;  ﯦː���  ?F�   �M�>]��/6ߓ�|��f��f���v|�d�}�r��L� ܀s��4���]��k=������˴� @����CJ��O n��   ��PJ��p��p��Ͼ�X�O+�c���l��l�٬�\.c� xOmۧm���f\co�.�����x���  ר�䘒�� ��	�   �{�P��g���_|o��g����6��:��&��&��*�w �gt]���>��O�mJ9G�5����&�   nHM�!O~  x5w    >�a(9��9����ߛ�f�l����:��6��&��&��:��|�����Z�%�.M�^b���ƈ�e�~~|� �m�R�OI7�) ���   �_���xlr<6���?��o��l�����/�x �m���{�v9��{�v���p��5  ܯ��cJ���_ ��%p   ��tZ?�?|���l��z��f��z��f��j��j����5 0��+�m{Z_���7M+�  �I�!��a �	�   ��Z�4M�������|��j��f��z��z��j��z����8����n �'���7Mw��ۦ˱i3KI��%Ic�  ����OM?�) � p   �	�Rrl����?/��֧����o�Z��Y�3����j �.�PҶ]��?E�m�n|<=ߎk�/��"���  �_+rHɷ�?, �� p   �+�r��_�f�Zf��d�Ze�^e��d=>�Z��^��xK� ܦ���6��q�כ�K����&�p�՟���G�:  ����&%��=6 ���   ���>]���z�Ze�^g�Ze=F��*��:��*��:� ��w���s�ޝ�׻��6��|��RSS�>  �VM�!O�w ��   ��.]�e�7�Y,�٬�Y�V� ~�X�N�i)�� �֚��uC�񇱚�{�y��mS�ie����}��# �m�)yJ��*  �5�;    |p�P�?��_�f6�}��ן}�Z��\-�Z.���Q�5]7���K��uC��K��i�6C?��<��?G��_  ץf�!5G���� p    �Q�5mۦmۿ}�l6�j��b�>-�/�Y��Y,�Y��Y��Y.�Y��Y�g�L�����)\o�>}?����mO�];F�I�Z]  nQ�1%��� �'p    ^M�5m�']�w��I��|��j��j��r��j��r��r\�_.�#��r�.�܋R�%X������;-�w}���Ҷ]�2$/�֟��.  p�j�q�}�� ���   �I�2��I���k�Y��U��E�eVc�\.N�j}�|q	���㼲��C�����u]��K���>]w�֓���9V��� �C�R�OI7�)  I�    \�RkڮM���u�\d�\e�\f�X�A���^,Y,NQ�l&��^�5�P��ջ~�����n|�O?��������R��  �(�b{�w5 WO�    ܥn�E�)t_����c�\f�X^B��b��r��b\��>�ZO���P2���0}Ώ���}�0���0��s��c��   �>5%MJ�
 �vw    ��0��>i~쯛%Y.W����s������s��"˅�x��yI����0}(�!exԇa�;bڇ�kρz.�����  ୕�)���O ���    ����뻤�~�Ϙ����c�ɟ��e�8�������cH�8}>��.����p��Az)��PR�)8/����1D?���PN�굼��iI�yE=��  ���ːCj��O �)w    �+PʐR���ɟ͒,� ~1�%�E��yf��%�?>��Ɛ~��|9>����>��/�$�b|��2��XkM)%����kR��7&�R2��2�kN1z�5������ׇ�d��Y��G�rv  �^�)9���� �_"p    �35I?���Km��#Y,I��b����g6����g�l>F���|�8�	�Sp�������Yf�ӟ?��$�/�_?��.���x~���şs�J���9�>���ה�^RS��<y~])C�D?�����W�$���<�=�����K�>��?��S�^j����}_>�a:  �YM�1%��� �ew     ~��Z�s����?����VϾzn>�/�[�q��8��ߣ�7��;}��O>.��S�~��{�  �ޜ���� �+w     n����~�������I�|   �9%�����  �O�        pj���S�O}
 ���        \��!%���S� ���         W�d�!5M�ԧ  ��;        �U�)iRrH�� ��        �J<��e�S  &!p        �XM�!��S� 0)�;        �Dj��R�M}
 �U�        ���a�۩O �*w        �wRSRrHM�:�1  WH�        ��jJ�)9�J� ���        ��Ԕ4�j�� ���        ��s�^�> �f�       `5�l�#x%��S� ps�        0q����2䐚~�S  n��        ���)9���� ��'p        �	5���S� p7�         ?���䐚&u�c  ��        �;� ޞ�        �oՔSrL�� �)�;        �7	� ޛ�        �35%MJ�v �w&p        =��e�S  >$�;        ��	� ���        ����  �E�        |8%��S� �w        ��� \7�;        p���  �A�        ܭ�.C��v �!p        ��)l?����  ~��        ��v ��&p        n�� �>�       ��U�f�Q� p'�        �ͱ� p��        ��� �7�;        p�JڔR3L}
  oH�        \-a; ��"p        �NI���� ���        WC� �	�       �ɝ��Cj�ԧ  0!�;        0��b�]� ��        xw�v  �M�        ���"l�S ��        o���Q{#l �o	�       �7q
��i��  |�;        �j���  ���        ����SrLI;�)  �(�;        �Kj��R�O}
  7N�       �ߪIfS�U��2�*l ���       �[�v�TҤ䘚a�S  �3w        �;�a{��  ��        ��E�^�> �;'p        �R3��IM#l ���       ����E�  �K�        ��KI��v�S  ���        �����cj��O  �;        |<�E�^�>  .�        �AԔ1joRS�>  �"p       �;W3�� �z	�       �N�t)9����  �.w        �3%͸�>L}
  ��;        ܅�"l/S  ?E�        7�f��65u�s  ���       ���)9����  x5w        �!%͸�>L}
  �:�;        \���v����  ���       ���ƨ�MM��  xsw        �25]J���S�  �J�        W���ۇ�� �I�       `B5%5ǔ4��S�  ��       �j�q���� �H�        簾���a�c  ���       ��Ք�4c�n�  ���        �HM?F�  ���        ^UMI;�����  �M�       �+�)�iư�^;  ��;        ���n��;Y;  �"�;        ����vۇ�� ��!p       ��Tӧ�IM�j�  ^��        �AI��cJ��O ��&p       �o�)�i���2�9  �!�       ���n���ԩ� �F�        �)���a�c  ���       �a��/��� ���        |05%mJ��� ���       ��� ���       p��k�Mj���  ���       ��S3��M��Z;  ��;        w���KM��n�c  �� p       �Yk ��!p       �Yk �{$p       �f��)iS�Xk �;$p       ��Ք�)iR�O}  ���        \��Z{���Z;  |w        ��y����a�c  �w&p       `r5ݸ��Yk �L�       �$jJj�1l/S�  \�;        都�KM;~   <�       ��j��K�n�  �6�;        o���MI��a�c  � p       �U�tc�ޥ�N}  pC�        ���!���^�>  �Qw        ~R5�ɞ    IDATMI��&%���   w@�       ���ư�MM��  ���       �G5Cjڔ4�)S�  �)�;        ��������  > �;        /Ԕt�i�  ��#p        5���ޤ�� ���       >����6%Mj���  �       |,5���S  ��;       �ݫ��Ǩ�KM��   �o�       ܩ稽�  7A�       pGj�Դc�^�>  ���       n\My�S�  ���        7�����n�c   ^��       �fԔt�iRӧ�N}  ���  �S�̦>   �R�]��E�  �=�  �#n   �5����L}  ���       \	Q;  ��	�       &T3����a�s   &%p       xg�v  �o�       ��S�ޥ��  ��;       ��)�iǵ�~�s   ���       ���  ~��       ���  ^��       �'��  ^��       �;��  ޖ�       �o���RҦ��  ޔ�       ���R;  ���       ����R�0�9   ��       ��j��t�v  �+!p       >��~��Ԕ��  ��;       p��W�;Q;  ��       w�~��^�>  �� p       �D}��މ�  n��       �Y5e\hoS�K�  n��       �)5Cjڔt��>  �W$p       �^M�rYj/S�  ��       W���mj��ԩ  ��      ��PSƘ��  |Pw       `25}j�q����   &&p       �QMM��v\i/S  ��       o���1���N}   WJ�       ���>5ݸ�>L}   7B�       ����~ڻԔ�  �	�      ��RSR/A{��:�I   �8�;       ��+���[i  �u	�      ��tZi�^|Xi  ���      ������ƥ�~�s   �@�       ��Yi  �Z�      �é�J{o�  ��"p      ��J;   �@�       w�������  �$p      �;Q3�Xhﭴ  ps�       p�j�A��v   n��       nFC�>e��  ���      �������:�I   �f�       pEj���?�   |w       �TM�,h/S   ��      �����Sӧ�K��h  ���       ��9h?-����v   �&�;       ������  �{�      �Ք1d��   ��       ��>��Ԕ�O  �� p      �TRҿ���   ��       ����^�   �H�      ��'h  �� p    �s5�l�#  ���   ���    �Ή� ���E���  �J	�      �;���几   n��      �W_,��W���G   ?A�      ���_�샠   ��      ��VS�
�  ��$p      જ���v   �(�       L�~�����G   �      ��Jʋu����   w       �HW��e�   �+&p      ���A{7~n�   �~w       ~�uv   ��	�      �G5�ʞ���  �7!p      ���  �i�      �̐O)�>   ���S            ��          �+!p          �*�          �
w           ���          �� p          �*�          �
w           ���          �� p          �*�          �
w           ���          �� p          �*�          �
w           ���          �� p          �*�        ���k�    ������8 w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w           w    �];    �o=��      � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � &<{    IDAT�          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          � �          �v,    0��z;���          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          �����(    IDAT          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��     �صc   �A����Q    ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,�           ,� Į    �Ǝ�         `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `A�s�    IDATp          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap       �];� ���7��}�SP   ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;,���          ����          p��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @��          ��;           	w           �           $�          H0�          �`p           ��          @�� 8�ڱ    � �i�(�         `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          0�y�    IDAT`Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap          `Ap       �ع�帎3��9(R� v8����݀o������[�inJ)��)�X@�Pu2{C�01�:t>Ϫ�'�m�{# ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R�          ���          ��           � p           �;           )�          HA�          @
w           R��2j{          ���W�.���O          �����;           �+}�45           �+}�w           F7��T�;           c+}�Z�^          @�J_K�;           c+})U�          �؆�T/�          0���Z��+           h^��P��          �؆>j��;           c+})��           ���(}�1�=          ��Ոy����           м���*p          `l�>"��W           мYQc�           �y���;           ����a1��          @�jt�����C           h�A?�"p          `T]T/�          0�ݬ�%�c          �uݬ_����3           h[�:��P��          ����Y���d�!           �����k����C           h[�������c          �m]t����/�          @�j�I�ݛw           FU���߻wg{�!           ���n�������           жä�=          ���E���}x�          �Q��v����           �k�~#bg�!           �m3�v��yl�=          ��m�����noXe�1           4k�yq0���^          @��#"�����l�-           4�M�~0;�w           {�*p��n          �U]to��0�;          �V�(�^p�/�ǝ          @���^�{6�           �&p���q�           Ъ��*p_�蟎;          �V��_p�y�'��          �]ݛ������q�           Ъz���͵g��          �U5�7�{�=�           ZU�;�{'p          `%6�E�
ܧ]�w           �����"^�_܎絔:�$           �2��#^��a�;�w           �����������q�           а����O���l          �aG_p_�ߏ�          ��}����8[           h������f�-           4�hྐྵ��p�-           4�h�~ok��q�           Ю���_?�7nm>g           ;��{��Q�           в����f<=�.           \���߾��C���w�yJg           �>�?l������:ݛN��          @���?����tg�[           h�Ɂ�|>��-           4������j�           ЪzZ��E��j�           Ъ��������          �]����K�~����1           ������־^�   >z	    IDAT        Z5D=9p�>�           �D�Ɂ����G�u��           h�bw��_�_t��t2��v           z��A�����ɋ��          �U_�}p$p_�<Y�           Z�E<|��H�>�V3          �VՈ#����}m}��j�           Ъ.�ف�ݭ{]�           ZU"�}v$p����/W3          �V�E=;p���W�          ��-b���gG���#�           �
�v��|��H���?�vg���j6          РGQ�><�GD���>��9           ���q���������          @�wxl�X_]�           Z՝'p��X��z�           Ъ���Ώ�����G�;          �V������cl���ﵮ          �Y5�ǝ��mƱ�          �����=<�ñ����龟Mg���          @�E�?8�ñ�{D�d��w׷          �F}q҇������l          �a��#�k          @��'}91p�}��G�3          �V������{����z�           Ъ�"/���8��          ��(Q����p'�^K��3	          �����������î�Ov&;׳	          ���z{�)�{D��d���n          �a_�����}�W�          �v��O�zj�~�֭?_�           ��v���>�h��?]�           �u�܇>N��           ����/�/��Y��^�$           �||zڅS�?��&;���          @�N}�=��="b:���j�           а���b�5[           hW���g�w����          @�j�����{w>��9           4��{?�O�f           �*��xp֥3�_���v��?��M           4�aį�g]:3p�����y|�=           ��F|�̽��������          �U]��e�-�߸���\n           ��.p���'���           Z�E����.����          �Qu=�?Y��R����x0,�r�M           ��F<z��Y��R��/�n1ٙ<��,           Z�E�eٻK�����.6          �vu����t�yc��          @�����~t��          @��(W��_l           �*���ɲ����c+�6����          @��z�.{y���뺲���o.�	          ��?�����������          @��r���
�o�~�Ϸ          �Vը:����?�����          �U]����ZϷ          ��Ԉ�����c�^�����g��K��]�V�q���"�ɥ!I�Ig��3�a�t���t&��B&��MHjH�@��8�6��&cc|�ecC ;Nl�b���V{;�>0&c��=��������[���=���G�'��ͺ�?�'�,��gח          @�I'#n^[�7��GD,�-|{��           �k�G��ź�}�ڃ��          ��RD�~�>4:|�z�          ���h|m�߬{��Rߺ/          ��4���c��h��o��+++���          ����x<>�ޏ�=p[Jks3sϬ�;           zC���F�[��="bee��F�          ��Q<���64p��F�          �������-[�ܿ��           �~��ֺ���z<�Xk46�-           ]���x��F>������tavzvC          �����GD,_�pb��          Н��o�7<p��F�          �;բ8��o7h�-�m�[           �S#�ֿ�2�����m�{           �����#��x��c)��M�<���          �:5���+K�6�=           ]�D375p޿��f�          �{4�q�������h�{           �F�[i怦�G���K��͜          @Wx��M5s@S��Rcvj��f�           ��5{FS���j	g           ��jQ<��M��f�           �ӥ��=�����}M��          �hK���Z��4=p��xr���b��           Щ�O,5{J���R�P��z��           Щ�}e����="b��mw�q           ��h����]ۿX�9           t��X���sJ��-Ń��F���           �E�Ӌ��2�*e�~t,-�L�<]�Y           t�Z���;�$��ջ�:          �NѸ���J���^�Y           t�v|�=�}���           �K���ZY��6p�'{��ٹ���          ��'"�X*�����e�          @[�J���:p�=4��2�          ���S�a��w��vW��          ж)�|��K��ǖ/,/�y&           m�z�7U恥�SJ�ٙ�o�y&           �➲�,u��c���*�L           �N�ܷ���Ų�          ��4��J�g�>p�k��E��(�\           ��w��#��>�����4_��?U��           ���*N-}�}�;*9          �v�9���ݷWq.           ��"u���o5�n�5U�          @Vgf�ēU\����h������*�           �ŗ�:���{DD�WU�          @E��:�������mU�          @�H�7p_Z�{WW�֪:          ��*"���OVu~e�c������Tu>           ��"�M��W6p���߲�U�          @�h|���+�����*�          �uVb�KU�_��}�`ܷ���Z�           ���.ƣ����ҁ��)-�N�~��;           �^��b�wT:p��ؾc�mU�          @���T���w����U�          @�)��������=�����J��           P�"�ѹ81Q�=�܏��R�����           ��"�؊{*�GDl߹�3��          ��Hӊ{Z2p߱c��          ��-m��[qQK�G����B�w          P��=��ɅV�Ւ�{J�8?���V�          @y��;[uWK�Cc#ڪ�           (G#����Z�Q4E��          �ig⑓���e�7�险�'[u           M�3"Z��y��}�6�E+�          `�Rw���v����           ذ��_h�-�s(������;�)�.          ��*"����ZygK�oKimn�~+�2�����          @v)��V�������Ѝ����w          zL�V���{�����(Z}-           �n~>���K[>p�f$����=��{          �d��r�/m��="���gs�          �%�=ǥY�{>��^           ^U�����,��Cq����J��          xE/ƣ�r\�e�~eJK���          ��K�>���,����{>��n           .&ݞ��l��Q��(�\�          �������\�g��qo:3;5�D��          x��s��u{��{D��-��4��           ��"����g��ܵ��s�          ��,o�m_��u�~՞�����T�           "RwOĽs9��#"�/~>w           q{���ѱ�r7           ���}�4w--.-��           �a����'rGd�Ki�>3{o�          �^�"n�������}���n           �U)�[s7D����������h��           �A�f��sGD�����@����y<w          @�)">���������v~2w          @�)�qk����}�͟��           �cf�vw���������|}�T�          ��Q|6��J����=""��M�           zE�[s7�X[ܷ����           =bikl�3wċ�����`zxnfn"w          @�KwNĽs�+^����k���          ����.x�����s}�          �.�ZD���/�v��F���ٹ��           ݪ���|<2����n�������           �*E��^N[܇��\��          �K��zKӖ��������L�          �n�"�5'���x9m9pO)+K����          �m7�n����GD��>w          @�Y�X���Ӷ��{⫋���;           �ȗ����Ӷ��R����-�;           �Eqs�WҶ���=�C��          �K4��x%m=p�z0�9��0��          ��}>N���J�z��Rj,/.ߖ�          ��7�nx5m=p������           n���grG�����i �Z�_���           �T)�/-��;^M��SJ����?��          Щ��ݘ��R���="bpp�#�           :�r��[rG\���_5�����=��          ��^���rG\���GD��n           �4Eč�.U���v}�(��           �dnw��#.U�܏�'f�f���          �9�[Nǉ�+.U��#"�l��H�          �N��vc��訁����7�E�          �0Q��sG�GG܏�J��'��          ��R��'Vrw�GG�#"v�a�          �vWDqc��꼁{_�ͫ����;           �U�xf.�7w�zu��������s�_��          Ю��OED#w�zu��="bxl�}�           �U�S�6�#�>�����           �8>}=w�Ft���HJ�K�n��          �nR�n�ݰQ9p���P�          �6�RD�#6�c�W�=���;           ���sqb"w�Fu��=�T�j飹;           �GqC�ft��="b��,�"w          @�����sG4���G�ӳS�S'sw           �"���R�ft��="b���{s7           ��r4���#��liq����          @��]���Ѭ��>�.�LM.w          @F��(C��#"F���'w          @&k�Q�d�2t����Hz`fb�t�          ��+�\����(CW�#"RJ��           �jE�>���,]3p�=�G��F#w          @M����rG��k�W�K�M��x0w          @�7D<����,]3p���7���           �҈�>wC��j�>=�w������           -��B<|2wD��j��S)�.]X�1w          @����.([W�#"�ޟ�          �b��Su����P����̓�;           *t�T<P�Q���GDlٶ�ws7           T�c��Е��ږ���rw           T��sq���U�ʁ�������_��           (_�XD�+�Е��������           %[.b���U�ځ������&���          �,Eħ����U�ځ{DD��-��n           (O�ù����}���'���sw           ��o���ݹ#����+SZ��[�)w          @�R��"wG��z�12��w����          �o1b��#�����{ӷ&Ύ?��          �	7�㾩�U���{DĮݻ;w          �F�(>���zb���֛�/��           ؀��x������#)-����$w          �z���*=1p��98z]QE�          �u����_�V陁����������           �tŧ��z�V陁{D��=����          �R5��P�Vꩁ�S�7�27S���          �����ȣ�+Z���oKimme�sw           ��"���=5p���7���˫�;           ^���(n��j=7p�`����-w          ���>qb%wG����="bwE�;          ��,����9��������ę��sw           |�⦅x��9���="b���;s7           �T����ݐK��߲�-�����           /�@=z0wD.=;pO)5֖Wޗ�          �)��}�=�����F޷�����           "����sG����ޓf&όߖ�           E|8��;r��{D��e�QE�          �������ȭ����M�>w��c�;          �^�nZ�GO�ȭ���C{~-w          лR���nh�q����f�f'rw           ���r=��]��#"�T����          �����.h�ߵop�K��sw           =�;s��gsG���r8��f���          �"��ED#wG�0p���#�����          h��m���1p�kFҩ���}!w          �><���h'�/���o/�"w          ��VV��������%����;����          @7K7-��grW����cp���           t����ڑ������w�1~f�t�          �_����+ڑ��El��{g�          ����]���]�_D��>Q�����           ������_�hW��S)�.�_|o�          �{�H�ED���]���ѽc��8~)w          �����M�#ڙ��+8:��3s���          t���/��hg�bl߾w���4rw           mzsl�h�vg��*�ޗ��<7y{�          �s��LĽs�;ڝ��%�76�_��          ra-j��	�/�ѽ�[�g���          t���q�l�N`�~����R�          ��E��~�Na�~��<����=���          @�H���׾���S�����]�9w          �Ij��]�I����.�y��g�>��          hEĝ�8~<wG'1p_��[�ߞ�          ����]�i����`�3�g�O��           �Y�o>�;���    IDATwE�1p߀�T{G�          �}�h�F�Nd�o}���M���           �O�H=�3wG'2p߀�Rc��ޕ�          h?)�FD����o���?2=1=��          h+ߘ����T����֖�ޝ�          h)�oFD#wG�2po7������|�Z�oS_�          �ۓ��ys�Nf�ބc)��_X����Ʈ�ݹ          hk��w���d�M�{຅��To��;          �"����O���t�M:v �����`���{�@�          �T#����r�Ng�^����7.,,�e�r��x�         ��uf>�|<wD70p/��é>51���Tk���         �~)һ#�[����Kr����z~����Tg�w          �ϙz�,wD�0p/ɑ�4?39���Tg��         ��(��-������D�|�B}�+�]jd���	          ��3���#���{�������������          �����g�^�7�\�����;(��;          �s����3p/�����������|{���N          �M^o���{����7�ӳ^q�2���-[���           ���|�~,wG72p���������{rwP�᱑�	          dֈ���'�rwt#�����׾{fbz>w�ڻ4w          y��Z�9������u�;(�ޱ��          Ȩ��^o���{����331=�����7p         �a�0�����+t,�������Ay�         zY��^o���{�������'grwP��Fs'          �Ƿ�b�'sGt;���-����w��_{(w          �q�j�ng���W�����T��w谁;         @:9'>�;�����RZ[���_rwм]��c����          �P��h����-��W�}��g���A��         �S��C���+�[$�Tl�����4;         @�("~-wC/1po���j���z�[�;hΡ�]�;         �("_���K�[,�m��F��;�&|��         zA-�]�z��{���k�?8qv��l����          �.E�x=N<�������SO[���6����;���r'          P��D��͹;z��{�}{��;w�޹=w7<:�v�O         ЭR�G��������-������*�9w�I)šÇrg          P�Z<�p{�ƻŏl˜�S�[h���۶sۖ�4���ȝ          @Rl��Y���?���5�-��b���п��A9�x��s'          P�����_��~e$~lW��d��"Ϟ>��͛�7���?re�          J���=����F�ʐӓ�[���k�����swP��y�         ����E�����jeO�2po�g��������g�EF����@�          J�^����X~{sz��u��)�=��_��|���	          ��U^o��)~io��X��z��{Ş�Ω?���wѿ�A����s'          P�[.��X��U��:�
=0~���v�?��A5�x��;         @�K�)6]���=�3�W���+4�����ռ�ޥ�         :�%����-��RU��9~��n޲��������������5��ȝ      �Z��h�J�   �Ц�)�sg�&Ŧ�Ŷ�~�RD�g�h�u^p����ɏ�w�m;���Çrg          �A�������Z��Qv�3p���KW��؏��zG�]�;         �H�96:�."��@���r��0p���鉏�j~���ț�ʝ          ������f��{E��K��٥��.�����Uo�;         @�y~ܞ�:�+��0p/�䙩�z��w\q��زmk�          .Y-R��qP-��Q�A�#K��_~�������A�l��?t�rg          p�j�%�}��E???�R#"�K5qz��)���N�8r���	          \�}�bS�G��X��{��K����C�ޜ���;r��	          \��_o/ݿ��{y�K2yv��z��7]u�r'          �*R�GD_G��X��*�E�%x��±�{���A#�Fbߡ��          \D��Zl���{9�K0{n�^o�mW�:w         @t��8Ŗ����+���zEg�����'�7��{m��:��?�;         �r���)R����"�/쉟���\�����SO��`��������4w         @����������-��/b��[qQ7��n�c3�����D�����������          �L���	�)6��"�G��6���	������j���P�ě�-�          *�y�Z�^o�x���+��K-���o�c��e��F6w��-o�6w         @e:���Y�S����򋻄���~��{�6����=��zm��A     ���޽�Zv�g�޵��g�[��r��o�66����m|s��@�I�� �\�	t�H�uOZݙLZ��iF����e4Ҩ[%ݚ!!9����Fp��r\�r՞e�ou�^{����IȖ����q���,=�   ��4[���~��7Jz��o���6|���{����9�.�Nݝ/}M�          c1K��~Jժ��{r�F� 3K�}���#�hi�7;�P&���\;         @�N��K�'�����Ye����r����E�޵g�O���tRp         ��,moo�<U���/��kWj�5
�[��~�W�˽�9�NW^����k?�         Э�٨ϖ��)��O����!f��������]�����5X]�eoyc�          ����%˵#����>ۓ�@�}��;�~q�6p��n����          :5E[�_RI?e��������1K��OpZ}�����럩���w�;oN)�v         �N�(�O{��t�.)_�����E���o�C+�+��s0�N}�iy��Ԏ         ЉY���d9�t.(&��-יִcV(�����KKK�������Ԏ          Љ��v�W�N}	�d���f���Ix�ۇrm��f�̎[�}[�          ����x;��۟3L޲+�\W;�,Pp?	��|�Wjg`��s�9��k�          �4opo�O�8����kg�
�����3o�}ꮳk�`����[jG          II�����k�؂�ݹ���SL�i�ڦ�������M7�}s�          #)Y��%5YNRj�؊r<���!����������O=c�e�s0�.�⒜~��c          l[I�v���Lq��3����xN��L��e���|�7K���:�"�����[k�          ضi-�7YɌmo��0�gk��f
�/���g�~��Ɍ����v         �m)iR�֎�%K)3\�&�ؙ�w��1�f�Ov̾���Z�kg��ǅ��&]vQ�          [6��ۛ4Y�bT%�d��J��E����S�캿v����g�          [V�T;�4�'������}��9�������w�}ayu0}�Hfҝ�;K}�         0[���^�N]��jg���E(�����K���O�����ܽ�ko��v         ��v�L>]U���:6����:��M�U7����d}s}G�̗�����          NڴmJo����v��]�37�\;ĴQp��?����?��yCv���v         ��ҤW;�i��pߝ��L����ϼc���Ϊ�������vϝ�c          ���2U��&�IJ����Sr�%�CL�rp��T;�����v         �WT�˴ʛ���3��3i?S;�4Qp����W�>}��s0�.������j�          xY%���U�,�1v%�j#��R;ǴPp�������30�~��Ԏ          �J�&K�c$IJ�S��\V{9���)��t�;���=1�S?�ݥ^�����v�c���w瑿}�v      xI�r(�s�v   *h��6�c$i�f�v�	~�@N;?�_��NR�"<�������_Png�^����}�c          ���~�I�&+�#LX9sg�~�v�i���?���z?W;���?��E��         Ӯ����J�)�Ys����cXh�'�����v���ű�sG���wԎ         �<%K�_/n�L���+���-7�NQ[�+�����ԗkg`�|�SL�,��         �"e
��M���K̇������n�~���M{����9X<�\xn�|�[k�          H�����Kz)�U�0޻3���v����������X\���#          $IJ�Rwszyv{��k�9���!jZ���thx��g���뵵�����a>|�������Վ      �s,�r<Gk�   `�zYO������ْ=I;�����õ�԰�����Wn��RJ~��v         `��������r���ٙ|�v�Z�����p�?��v���o��\X;         ��j�ۓ�&�ϟV���NP�B܏����v�o��M��C�j�          X͂y�~���
ʛv���NQ�B^O}奔W;<��{��9�[;         ��Jڔ�*��V�?ݎ'������+��Ɂ�U�O����9�9M��?���1         �To{{I�A��gƏ���g�1iWp�ۏ�v�Qo��μ��k�          HI�Tڠޤ��xU�Zz&�|�v�I[�����3v�ټ�v�QM���_���1         �R�O�:�b{�b��~2�j�v�IZ�����?��څ���?v��y��WՎ         ,�&�U�-�T9y&�j3�b���=�^��d��r>��O��l         `�J��L~1x�RJډ�;�J�P�)���c�޾����vx9��卹�=o�         �su���j[�g�ͻsۥ�CL����}��[;�����CY^Ԏ         ̱����l2HR&~�<8����aRb��7��^][��KS|#�z�;�s������z�(      ,�a�d��c   0&M��-�ONI?M�R��dw.��C�/Gk����~�5m�����ɇ̞��Ԏ         ̡&�>�(��n��s��!&a��7�K��¬�g>�����_}�v         `Δ4).�7YIbW����'jg���/�_��ػ�7�7k瀭��޻r�Mo�         �#���^���v�gΫ�\�37^Y;Ǹ�}���c��T;l�/���.��^�         ���L���L�P?�i?V;ø���?><w�����4`&�ؽ�cǎ������      �@�9�a�׎  @ǚ,O�p�f%��{�Jr�j.���_���e\�������ϗF�������y�_;         0�&Yno�Ϝ��e�X�_;�8�m��k���`u�j�Q-/�����iڹ��         cV�KIoB�5),�/���jg��m��}䞵����9��^�����Վ         ̨�noWn�7��-o�b\���āC_�����/~2�_|A�         ��)iҤ?�������?Z;ø�����?6������{�k��Ͼ�9�̱�Q      �c�r(�s�v   :�f%MV&pR�6��ӊ�y���g>��?T;H��r������r;���W_�in�         :VR�d0�����>1�Ϥwo����е���~�*���ԛ�{`��x����Q��7ߩ     �95̑s�v   :�d�&��6�di����ʞ���];E��n��ӏ{����Z�0.M�����W��sG�(         �+I�,O�&e%z^�Sr�%�Ctm�
�����`�N?��|�7�v         `���SҎ��&+9Q�gҎ��H�]�;Q�|dx����?-M�a�]�������?|�v      ��0G2���1   Q���1��n����X��e��pN�g�w��?��j����?���m��Y�����򷼱v         `�4Y{�MI�g��Nߙ��k���\܏?���3�$��z���ײy���Q         �)�d0����$�L� ]������^��k��s���~���������          S��f�����d9sTE�uw���g�ѕ�����_��j����3_y�v         `
�Y�	���ْޱ���!�2+���[ÕՕ�_�K�^�,P�믾,���˟���     �7̑s�v   ���M�����d5%e�g���_�V�]���r������9���~�s�ꆫk�          *i�:��M��S�\�3��X;E�����C�X;L��R/_�7��W����Q         �	+�di���)�m>��d�]���'��x^s|�����Y�+{��7���������Q      �A�r(�s�v   ����1ܛ�Y�l�1|b5;^���o߯�d3���о��Rn��;����O~�g}s�v         `ƽ���`l��J��T�xO�����p8,�����9`]x�k���7���/+         `:�Y��~�vl������0��.����ܲ��~J�0������ʿ�Gi{~�         ������6M��2���8%��U;�(f��~`jg�iw��7�W�寥ig��         ��6�c�\�d0�ٌGi���j��̮u��}�Y��n�43�3����9��3�������pX;      Sn�#�x�   ��&���ЛR��lƧ$g�_���sl�̮t���c��z��K��;~�]y��)���Q         ��$MV�4��U��������!�kf�����`�����g��k�          :P2HI;��el[ᙔ�õlW�W����W�W���XE[��k.���j����jG     `Js$��  ��QR��FN�q�V�Ք�ݣM�dx����g�wf�?�g��{���=X�F��遟�P>�֎         lS�Ռ����Vx&���+w�N�3Yp��я�� ������j�          ����&�c�ܦ�e.u��N�3�x��_��2�{�s�<x˭������o���Q      �"��03�s  ��P��YO�|�uI���c+<u�W���p����Y�b�6�����E)%_��_ʵ�_W;
         pJ�S���Af�Z��(�`�g�[;�V��U����� ��˯��_�믾�v         �e�4i����&Ki�P����<P;�V��;����-����������w<���ߪ     �ʎ�P��h�   ��^6R���̒&MV3c�bNޱ�i��^��Gj9Y3��}���?U;̫�ݛ����Y�ܨ         �M�;/�'I� ��s����}�Cl���o8lW6V�_;̳�.:?_�W����֎         <��M����6�Dgp�3|�v������E��m+����9`޽��k�<T;         �����Z�޲^�4���L�r�fn<�v��53��{�}�vX�}���         ^����:�YR�d�әL�Ҥ�@�'k&
�������|'b,    IDAT�������s��7׎         ��R�:�[���7�3݆>P;�ɚ�������_^�LP�k�����_wA�(         �pJ��Y��~J���2���r�j�83Qp?��O�� �hmc-�����l��Q;
         ,�6���[�K;������N���>8ܽc��kk�Eu�������+)ūH         `�,����̒��A�3�-%��L}!t��G�:vO�k�>'̳���<�s�         �^I������R����X�v��kj�x%S_?x��Gkg �O~�ӹ��WԎ         s����Z�^�]�OI�ә̦6�﫝�L�c_�?ܙ������a�����~"��     �1:�C9���c   ,�6�i2�tfI/MV:��L���$��R��8~���)���8�������J���         ��di�����Lf�y;r�յC���n�>����jg ��o��|��         �FII��1���t>���&����r����g�7v���͵s /��/}*W�xM�         0���t\�-駤��L��0�dz�|�ڂ��r�K�^[;�BM�������N�         fZ��4�w:���&˝�d����[�T;�K�ڂ����D��K;�S�˿��2��         �T+i�f��%%�Ng2�﫝�L���ח����4������ͣ�y4��7��v      :4̑s�v  ��VR�f=��:o�Ք�݁��8�p����b���=R������j� ^����_���S;         ̔&+)�.�d���<s����ze�/f*��������3X]ɗ~��         ��4YJ�A�3Kz)�w:�y7��v�3u�h|���Օ��o�m3uـw��g���Cy�k߬     �s$��  `.�4�eG����&mV:�ɼ+�u8��k��QS�r��;�����R�����?��_wA�         0�J�6k鶈^�(��-傝����)~����w��3 [�_��˿���z��         �Tj���n�@7YN��J03c���	~T[;��ڷ������i�v�r'�3���#���z�(      �`�#�x�   s�I/m�;�Y��&˝�d��:����C���z\ci9o_ZZ���`�~����W\R;         L�����r{�*�Ӂr�f�vA�?l�
�O<�ă�3 �i{m��_L�N��         �i���im��� I�p&����{kg�am� ���p���t�ݶ���3n�������p�(      l�0G2���1   �B�A�:��f%STf�W��m�ϙ��KsC�_����ǿ������j�         �jJ�g��]�\N��t&��\��N���9SSp�C��� tgmc-���C�c         @%%m֓�g��d��y𬶗޻j�x���Ӕ�֎ t�m�#��~]�         0qM�R�v:�� ]�����v��L���Ǉo(�7k� �����[��u��O�     ��t,�r<Gk�   �YM��f�É%MVS�h�5s���O}$���j������O�W;0g_pN>�Ѓ�c         �D��i����&������9zg�ɔ�?}�����ɇ̫_{^�         0V%%m֓��f�(�/u6^����N�LA������:u�kj� Ƨ����~�)��_�         0mڬ���l^I��~g���3��W;D�����O��h��ܻ�7��w�Z;         �E�A�e�&MV:����ޙ��ST/�?q���� LƧ��g�_�$         󥤗6��K���;��rw�U�����Sw]S309g�wV����֎         �))i���ԕ$m�3ᕕ䝵3T-�o�嶥��R��d}�s�����1         �m�R:���Ӥ��<؊ar���ښ��t��j�L�����/�t�         0�6+)�w6���&˝̓�hҼ������2XY����@=�|��s��Ԏ         ��d)MV:��d��<ض�k^����\����Y�|����R>�w?U;         lKI�6k�K���;�mxӞ\�Q��j�C�{��Zg�����s�[��         ��D}-]�pKI����hJ���o�uz����g��W�l`:|��O�        0;���d��y˝΃n����U
�����s��g��ҫސ��uk�         pR���d�ټ��r;�ꝩ�5�r���]�6I�3���4M��I         �I)i�f��y'��:�L�r�fn~S����J<z�������/�-ﾭv         xI%%m��]�(�3�ʉ-�7��p8l��W��������>f�;         S��ZJ�筤Ҟj؊�k:�o�7����ڠ��30�zM���)�v�_|An}��j�         �h2H�~��,��]��;N���/��С�N�L�Xi�֓=�ɒ��x~����        0UJzi�ݦ�&��,u6Ƭ,���7O�M���G�?�3�������d����{u�0�lq        `��4�e��ymJ���a��1�3'Zp������{v�v�g2Y%ɫV�s֒�����{؈��/|�w         �+Iڬ���m�&+�N��1L�̄/܉6I��y[i����5�y�ɞ��k6�sλ����^[�        ���jJ�+?*�3�JrƮ�v�$Ϝh������yL�J�\��қڗ����N�G>o�;         �4�ɠ�y+)���B���;'y�D�-�����<����O.�x��K��ᇝw���靷Ԏ        �*i�f��yM�n��J��<ob�?�7|���ڮI��d�6H�ZK��xkƺ�3'��jG         `����YOr�ȓ���ہ�7��;�{��L��~��'u��$9g-9}��o�k�ќ�K��4��卵c         � J�6�)i;�ئɠ�YP��<}��X���C���I��x�%9o#�����z%Y���ܻ��>T;         ��jg��K��Y�dL�a��:k"�?��pes��u�s��&n$k��}~}��c�������מW;         s�I��m�%MVrb'<̓�|���rs��Sm�qk����Ѷ��w�p�i����Ԏ        �+i�f��y'�����Kw�m�N⤉|���w���8����O�[Oz#^1����b��'ޕ�Sv֎        �*)i�����7YN�[�a��3�O✉܇%wN����Ar�Z�tp�nK2p��$-���S;         s�$i���Q�����~'�`zo��)c/���'���ص��q��x��r�]�X�v��ޏ} ��~�        Н&�)��X�K��Nf�4+)���W���܏�-���� t���ۻ���~&�kש�s�}o�        �9�d9M�*H�΂�w���vɸ{������;�3�VIr�z�{L��&��s��O�_;         s���6��j�d%Z�,�a��:�3�^po����t�I���d���n��%��������%W^Z;         3��I��tSH/)�(��`��lܿqhx������y�iKr�F�1�r�svL���{>rO�         ̨��6�)Ug۬���d̘[���z��~���J�d�,�5���6�o����qϝY�ܨ        ��d5%ݔ��v���<v�8k�}����?��t��&n$�	�k���d-�rǽwՎ        ��i3H��Nf5YN�R'�`v�u���Zp7�s>��7���'�:I%Ɇ�;[��=3        ��k��&��ꥤ��,�m�qN[������k��q�gt�&9c����(��U�y�ks�Uo�        �PҦ�zG�z)t2f]InL���c�6����5��-U.�'ɺ�;�`�;         ���<[n/�j�d��,�k����5|l��}�<~ϸf3�i(�'I�$+m�̞��3;wԎ        ��*Iڬ����bI��(���Sn��U�W�W��l���l�}�r��9;��r���`9w�{W�         L�&k)YyNI�-�OI�����qM�7�O�_����k�پ^�\�>=��$������v         �P��4Y�dV�JG[�a.�5�o,���Ru>z����1���5������gWڤ����ҫސs.<�v         �H�^ڬu4k��^'�`N���ޫ�1x,���|�8�=m9QnLY��9�����sg�         L��6m6:��d9%ʍ�J���8��c)�����\��Ir���w�����^;         S����z�������G�$7�cn�����������l]Ir�z�:�o�XWpgξ��\|�%�c         PQI�f=%�o.i�d0z(X�'�u����{;̏u=��9k5�1��^IV�x�<��{�        ��������d�&+́���3���록�������g�ug�$��k�8y;�̓mx�=w�i;��        0�:ڸޤ�JN�����]O�Zڦ�l�)�ɩ3�����4���s��\y�U�c         0aM��f��IE�FP�����N��o�cs���]�dkv��Wuq����6i�n`n����         ���6m�;��4Y��E��8��t�'o-M��\��Rr���>Cd�;�q˻nM�_;         PҤ�F�hK����=,����#7��˙���?v��.�q�V�䜵��j�=ɦ�;۰���+���v         Ƭ���zJ��&���:H�47v9�ӂ��#G��r'�m�sדv���I��4�}�����n        �)IڬuRJ/YN���Е�tZ����{�a��g�E]���4I^���;}T���$�bn���OG         ̭&�)�w0����9��\���j����K��v�Z�6G��� ���W���^~q�         �A��4�<���IIx��sé]��~�ɧn�j'�A�s�����6]׍�#         б&Ki�6�޳%�2z(�G��4o�jXg�����Y����䴕�)��+󵑞ɹA�        `���i����V���x�k���Y�}mc�f���mr����f7�l+=�q�_�3�=�v         :P�<[n�-٤Un��+N��?~lx�����.f��$箝�t>�v,�N�����kG         `D%%m�S�v0g%�^ڛ��{]��[����^�Yk��h�멷�$�9����r+        �e%I����ړ-)Y�r;L����]��[{���o�b/o�r��_;�dl.��I����VWj�         `����d�aI���v����]��f�{i�M��6y��v7�j'`������WԎ        �6�YI���s�R�v�؊a��(���_;vm���0���$笝��Xn���؆�n��v         ��I?MF�\���^������v�ʦmT�������E�9�FXHW�xM�         lA�^ڬ�<�d�F�jz�Zn;}�!#ӏ<�T'M{^����-z�X���Yt������c         pJڴ�yN��4Q<���y�ͣ�������w�:��o�3F���Z�%=�`����?ve�         �������e�9M�)Y�m�0e�'ou���ᕵ�+F���$g�&�h��g�;�q��W׎         ��()i���v�9M�R��Q*`T%�Qg�F��=:�x��6j^�A�6ҟ�|��'�?];�檛F~�         cR��YK�ƚ��������;`��G{�����;ƻ��KN]��b:��l�g���9�Sj�         �E4YKI�%�4�D��"�6s����~h��7��y^�$9s���9%��R�̚RJ�����1         �mVҌ�u��M�M�0���f�Ϗ��'�w�(��N[IV��)��Noa.��#         �C�,���ަɪE�0�F�R<R�}m}��Q>���d�2�����HW*���7��v         �դ�6k#�(i���So�\=��]~��p�����Q���ZM���ͥ�	�5����/�k�         Xx%����I�����v�We����?x��\S��DW���^��k��2[�_���K.�        `����e#��KJڬ�(�ì�8%7^��o��~��7o��<_�$�j��n��di�W+���+/�        `a�4iG,��`s�!̒c)Wo�����?���7o��<ߙ+I�CE��w��bw        �*Nl]�H��^�de�@��~r�����5�����M�퓢��V]��        0q?(��#Mi��a����'���x���Ս��=�8su�o,�A�,�򻎅s��.�`u�v        ��Q��YKIo�)mV��
�@eW$7o�F����3Ky�v>����'+�[b�;[ѴM.���1         F�Ք�R�+i2�r;̺��+�/��'�Up?�������w�v�٣��V]|奵#         ,�6+ϖӷ�$i2q�;0-�)Wl�s�*�?�ԑ�������d��-�7���5�]t~�         s��r���0��dE��Jy�v>������`[����۷o�-�l���ޝ=IvVb?�ws��4�I-AjF��	;��c���y���y�x<�-K�%���/�p ��+�kI?d5����2�����@�u3��*3+p��ϵ�         ��j�u�ǰ�k�r����������y2f���_�w��s_�|�         k���.�|��.��W�J)�y.���N���5�x�^x�l_�i        `���Pn��k����g�z�3��}��ߜ�><f�}>�Zq�>�'�k        `��t�e'��G�g����BKgz��3�o�������a�$y�z�\\\�-�M�/|�u        ��QR�]��^2Tn����z�3�{�ޙ[��\$C��s�+ɶ�5Nɂ;        �|<*���WP?����
X^e���tZv����Y��������6NI�        ��J�Q���k���Y���y\�L�~�?�^U�a���{�S���Aҝ��&l���[G         Xi�(�׌��a������ݳ��L����3O�3��u��S�\�>�)��WZG         XY%I�����f����B��$��,w8S���7��ߞ-I2�m��qM��SMƙlOZ�         XI5[)X^����`SM3�˳��{����LǓ$yq8;{���f'�I^x�F�         +��$5�s߿(����Y�>S�}�3��������兲��i�xE�        �,��S3:��K����ɟ����i���;����#m�ä�o_�k����ɴu��w        �ӫ�f|����ہG�Tp?���^Ϳ*��j�AMr�k���j��o��e��        p:5�t�����ہ'\����S�=�����ÿ<_��uu8+_�x׼r��(�        ��f�.[��l�}8�D�:�Kw��Sׯo����t�8�K�������x�         �7+�o����ہ�d��L��J���]2�N�9J���y��
�         Ǫ�_h��Zn���̿�>ޙ|�\i6�^�/�5����;���        ��JzG���\���Xn��0�??����������G�,]Iv�N_�q����A�$,���         O*���N�[n/���)�L�,���IǞj���4�⢡6��������q�
�         �0�r{Un��    IDATN��^ϗ>}�#OUp���g�Y�z�n�Z��o����X�        �����SUI�R3Rn�d?�T��S�*����.gsl��Q�:����d��:�h0Tp        H������e=�lj2��{����� /�Z'�3�0��        �Q��(���p~����/f3�k��5����l�>�?���:        @3���ݹ��\�4�_��k��M��+�v�_<���:H�g�+I�Z�`��Z��`        l���.��,��Ԍ�ہ)�~�4ǝXp��?�]��}
W�������xZ�        �<�r�NJz��l��<���r}'_�q�Q'׻��\�q���w��_�m'�����         .����c�v`nz)_<�����7�8����u���0=Pp        6�|��������'sb������v>q�WM�;h��'��gK��Ⱦ�;        �!f���s��;�v`�<������v�I��N��X���[G         X�������]3I�ہ�&/���n�:�8�����u}�8��$9<<�t:m        `�.Vn��2I9�^
pN�/�t�s_�~��������d�<W��R�j������         �P%I�����b;�"�$��s���}:��O�g�\Z_vם�A��w        `}���۩9�*lIMUn.E\I���x�+�Ç�_�o��s�<'9q��{��{��;88l        `!-����^2IQn.I��������?�7�^&�dصN�i�`�}��﷎         ��r�y�r]j&))s�p�i�_x�ן[p?8����^���D'�6L��ߍvh�        XC�9��%]���v��M��/�����7��(Iv��SpZ]I����h��#         �����L���P�?~�ן[p�ޝ�4�8�c���������\}��q��        ��������-���xlE���O�'#��c\�N�YMzɨk��V��:        �\���^38�� ��sɗz�}�؂{W�?���j��~���u�������#         \����)&�ہ�zWr��}�؂����c�����J���nc=��a�         r�����v`�tt�W�-������z1aV��A��W-�5����=w        `u���>J��#�l�^p����0��+�V�u
.���V6�w        `E���^R3NI!� .���_9�]���ńYmW�pVW�&;ޯ7·��       ��s�r{�QJ,�˩fz��������YmW\�c-��N�e��~�         gr���(�Kl�������n��Ε�EZM��L�ޯ��^2�Z��2=�g�        X%�+���r{�����Vp���l�����J���z��Y,�        ��$��*���L�ہU�µ���d?��~l#~�]�N�<]�V���[p        �ܾ۬}�r{�����B��4���۟�J�����b�qVO�&�^��SIr�I��{
�        ��z\n?[����.[G� �J�3GٟYp�����Xl��s���0���)>��        ,����\��~j�J�h��{֭�\�b��EFYE����R�$W��n���n        �)�r�Vʹ�������y�n��z�Yl��ҫ�V�u
��Q�\�[��j        �-����^3L�(IYL0�K1��n}f�}<�Xl�ղ����F]2q�ڻ}S�        X����3ݯft�B<�r��n�}:����xg�V��k����7ﴎ         �������� �j�r����s^�z�3��7QW�-��kow��}ׯ�{7��t�c         nVn�9g�]�X%y9�wO�T?U�=,���DZ�����Xq_g��4wn�K�q��;        ���r���%%5�'`�+y�Tw��{�O_N�հ�J��0��fXK�n����A��=?�        ��*��{�r{=�<=U�X%���mO���ֻz9q�_M��j�+��A�,­�o}��5�Ԙ�        .Ǭܾs���.5�<��	�F�g���W����}�r�,���E�Msc��+_?�o�y궒AjF�         ��|��^J&�h�]����Z��/#�*ص�q�5���}�ܺy뙷��S3��        �"�t�{�r�l�S�	�'ܻ^���ɲ�J��^���Q�s���c�V�K��        �YI�^vR��j�f��a���Mq�|��۞z�o�o\N���Kz�Oa��d��:�t�����e�g�$        �YI/��������qJ���t�iܷ�l�\N��v�{�F{Ɋ�Zy���NqTM�$9å�         �4+����+�%5���`Y}��>Qp�����~�+d�m�mқ��zx���)��΁�2N�A        8������%55�Ü�������������A>s�y�ӸK��*kˊ��x����g��F�q         N���.�9K��d��l�;���?��=}���&���J��~2��a-���Y
�35�T%w        �j�δ�ޥf�r���Y��S����ܻs�/7�r��N�����;ӂ�c%�Ԍr��        ��-��NI?5��%��_p����/\n��ӯ��j7G�f�����y����}�Tr        �V3J��3�ht�G�����?�i�Е�+��$7��Spwo�ˇ�>��c��R3�/�        ��2N��)�.��d��L ��09����Oe�m�['`�\&��V�{�7��)�.��        ����h4�4Jj�)QPx��.�w�����Y.5�V�u
�M-�V�W�{oϧ��$%%]&)�B        ��$鲕�ѩ�Q3II��X +m��H�'
������Y.;�Y��tc�{cU�;���fgS�8�        6�l s�ݡ�hP��|(�+����d�u�q�ˎ�p��$��Sp�\p�����;        l�G�����Jz�2N��N���ק�a4��
ﶂ;�qc4����ݷ�]�c�J��=>        �ެܾ��ӕg��Q4� Nk�b�ޣ?}Tp��^^,es_L'���D)�cP��}
�jz�o/��Kz����0
        k����nJz'��f��a��΢����O�+�]^z��b�z;����ǎU��o�Z�s�tG%wg�        ��(鎖ۻS_3>��; �������6��fܧ��	X��\��R���X=*���LM        `y�t靲�>[y���ir�ѿTp����mg9��o��U���������y������,        XU%�����o�K�$9��; �V3}z��έ;�o�fI��O��s
V�W�;o�>�����5�Ԍ.�y       ���駗��f����I��T�yxz�}����m�,��$Z�`UXq_o���f�]�O�I|�        �j��;u�}���v��L�Up/��m�,�{
�����4N���Os�"        ���Q�l��Ȓ�Qj�1~	0?�L_|���.{�ލg�9�9��F�p��~�v�Ij�LRҵ        <C��ѐ�IJj�)�/<����Zp����Yw�Z'`�;+����߾�:�l       `ٔ$]�R3>ű�.i����h4��&���;���������˰����/M        �TR�e��}�^j&�X���+/>���^m�[�6a�����	X%Vܗ�ۿ]���L�����:
        l�Y�}'%'��J��} .�'�_���d0����Y��['`�Xq_N�yk	�IR�K�q�3:       �R��t�M�ɕɚ�)���9:��&I��M�,w�j�%���)x��~���-�t��I��u        �%�Q����NI��T� �M�j�t%9*���j�8K��~r8m��U��u���/�l�D�K�S�	        X��^z�M9�M\M��S-�0_����+u�\igy&��u
V�Ȋ��y㿾�:�)�Ԍ\�        ���^v���W�K���� X����~���	��['`Yq_.����gJ�Ǉc        ���a�S����x �S���Q���w_jg��Up���/�7Wf����^�LN�        p�.�t�:�qj�Qnh�\I�
�>��J�0���~2m��d�}y���o��pN55��t��        �J*I�l�������.[)�]N0 N�x����×�fY.���Ã�)XE�.�:h�����y���[Ǹ�rTr��        gQRR�}���<]J&9�Q���o�Ͳ|��N��zy�B5���7��Ã��1.�f��Q|G       ��JJ�줞0,Y�;���X&%��|t���z�0�H������I'��P����#�MI��RI>L       �qJ�t�MI���S2��XN�����������:Ͳ�����<J�O@ͼ�7[G��ه�I��!       �SJz�e'%�s������@;�L�<�up����w��:в�?L�N������f~��_��� 5%[)�        K���^v��G��LN\w����99zE���n�eIݳ���dŽ�_�e�=)IjF�q�        ��e'�fͳ���e���< ˡ��ྣ��Lw-�s]I^�N�y��i~�_���P%��L���N       `}u���s���lFy^�e����g���:���0��lt��~�ܽ}�u��+�J�]�(        piJ�.[�?���qj�QnX)��[ܟi�0y`ŝ�V�/ݯ~��.MII�$%��Q        `�JJ��׏Suj VTy������&�ǹ��:��aү�Sl�_��׭#\����m
        멤��NJ��9��.��t���9*IJ���J).�qw.���%�\�_�ts�?�d�.㸤        릤K��箲�R3���*+y5�۸n�n�N����'��!Xyׇ��I���W?�̂�̣3P]2        ��P�O/����ԌR3�r;�껕�[u<�α����S���/���a���߶��XM��g�       �*���N�/���l���� X�^��:[�Xz��['`\$c+��O��]>��a�K��f���        ��.�t�:��%�t�<w���S��:��>ɝ��	X/�`�B����na��R3�K/       �*JJ�l����U� 5��� �����:��~��ɴu��N?��N��^��/ZGX:%��e�\>        ��6+��fp�]ƩF�`=���:+��d�0��u
�ŧ&�����z�K���f�r�        h��K�ݔ� Z�e+9�� ����v�������k��u1z����)���fxt�&g�       �<Jz�e7%ݱ_�ي���+9ܪ��Ӹ��:��qR}֚�޻�w�|�u��7��?��        ,��Az�ɳ�,�G�] 6�a�]��Q�+��^r8m��uѯ��-�����#���rM        ,��Q�l�Y����.�.? ͔��:��~*�I��N�:yi��j�������u�3���{         �kV^�J��1_�R�����` 4W��:�Xp?�;{��Nj��ܙ�����VR� 5�<�O        0_�r���Ì�>�$�, ��0ٮÑ��i)�3oׇ��I�s��s+��$%.)        ��t鲛��3�Z3>���f()�:y38����a�����q������y�o����jJ����        .���^vS��"hI��IJz��L�9��X��,��N����'�>�]�/~�_sx8mc�$5�Ԍ�O        �K�0]v�NJI/5����ұ�~w�Y�W&���׿�z�k����I�        .��8]������8�x�,�����	XG�.�:h�bu��;?ma��t�JI�u        VPII/�G�'��LtS xJ��ǣ�9V��a��A�����Iq"�������fg��,Y        Nk6�����W?Kz�2II�  �n�2�Ñ�����:�hP�~�������/�lc���e����       ����wS�{�k5ãEwc� <�4ց����z�:��Q����L~��g:�����љ�O��        IR3H/;)O)���L��� W�a������~r�O�Ԓ�4n�b����?ia��ԌS��(        >��8]���:{I��޵	���k�����	��J�ׇ��g�S��k
dp�K��        l���.[�yzٳf��Q=E N�����^�����U+�2�N����u��Tҥd˙�        ����Nj�O�^�yr� N0��SN<wi����[�X~o���|�ޭ�16֣_D��       ��W�K�ݔ����p" 1�΂���&�N�:{u��œ�����@��Aj�)�c       6B� �줤>q�P��*�Z���yݱ��jrc�:�r���:GJz��$O��       �z�2N��||����f��A�zpA]�:�9�[
�,�K����cYp_65]Ʃ�       �����������R2I�." �0��vڳ�uo?ٟ�N�:�%ye|�q��������k�<C���\�/        려K�ݣ���j���Xm`N�)�v
��6ͬ��tu�Lz�S,�~�G9�?h�c�tG%w߼        ����^v>��^R��!�D��9*��Z:���[{��	^����|��#p���qj���        p5�t�M�xH�����O�`~JW�j��"n�͖�a��]rMG����UQ2H�8%�o        VAI�e�.[���f��Q�u�@��N��"�{��S�	^'�υI�����������ܝ8s       `ɕ�t�=*�?���$%�(��`�v���E��k��MЕ�q�����=�?h�3+���f��        ,��.]vS���m��%w]C .EW��7���@��K��0�����������A�����       �����ݔ�NGIR3L�8��<�ZK�`xQ��S�	J�OMZ�h���A�\X�����V       �JI�e�.�yTd/�)� 40M���
��pۊ;�d��\��ύ��4?�����8�       ����.;�}��Q�]���W��V�sqK��K��qR7�����cn����1���^�LRҵ�       �1J�t�MI��[jƩ�*��Z��������N�����ưu�6���h������fC��       .Q� ��~4HXҥf��^�d ��y���:���Q2�����|E�}��R3v�+       ��2N���h��fxTn�� `L�ޑ�����	�$�$�NZ��\��4����Z�`�Jz�       ����^�S3>��u4Ms�'�C�9���N[�`����+���W?�U�����cp)JjƩ����        �OI�.���Kz�2II�8 <�@�}����o��M��8�6����/�u.Y��%�        .���^v?*�׌�V�7�t����>o��Z'`��j�Ҩu���*�o����-��       8�.�t�ɬ�ޥ�VJ��c��(��ۭ���u
6��d��W:<8������1h�$���8���        �UR����R{R2H�I�A �����՜L�{��S�iJ�OOZ�X����ܾy�u��f��^�         K��K�ݔ���LR3l N�Xp_�[{���ƽ����W��:K��f|�5w       �Gj�e7%]Jz�2II�: ��T�}n�%��!�H���ޚ�}�yR� ե���s    IDAT        R�t���vfっԌc<��S�`�0���:��+ɧ&�S����~~�����*���2Z       �ƚ�'vR3JIw���o �˂����k��Muu�l�Z������r����1Xb�5�q���      �R�K/�)�f��I�@ V����|�u6٫����з���X%��l�d���        x��a��&�R3Iɠu$ ��Eyx���o��M5�G�S��k���i�ԌS�F?         SR�e+]�R�?�߮u, ��E�`�u6ً�d�?��w+?���Z�`���       XG%5]vR3��`i ����_���i�l�Z�W'�S\�k���I�<jj&��/r       ���駗+���ZG��>Pp_�������)�d;��ʠu��y��:+�d��Ioy       �j�2N�ݏ�ۍ���������k��M��qҭ���o�ͷ[G`�.ϵu��       �Jjz�I���l�d��.��D�}�n>L��C���5ye�:����g��;o��:kĚ;       �*Jz鲛.۩�Xm`���;L��N���>L���S�ݷ��[�#��J�t�8�       XZ5��s-]��:�� l��
���^��|z�������y�u�VI�0]�)��      �%QR�e;�\K�8%]�H p�,�_���i�l�AM^�Nqz<�w���c��z���d/q        ���U鯦����j; J��2�&��[����(��I��������c�JjF��/�       @5���B��Zm`�M3Up�,��Z'�Yu�3[�Q���_�]�l��~j�R�k       �%%]��ϋ��D� ��*�_���i��d�%/�Z�8���?
�\�����њ;       ����r-��`� �Xp�D���]+�,����p��d��c���?���+駳�       ,H� ���.;�� �R)�>Tp�D7�Y%�g&�S���园#@�z��>L\        �������JJ�� ��)��/���i�03�%/[�x�o���;ˣdp��ė=        �^IM?/���1� �6�����%:�&w�[���^'�%{�w�^~����O(��Xs       Υf�A^Mͤu Xj�L�.Y�u��|�:<VK��}f������=t&�i��>��       �JIM/W3��� p
5���~�n�%���)ౝ~ru�:�c�W�lNP��       '�駟��˕�Q `eLS-�_�i��[��Ozu�����{xx�o��ߵ��R28�l���      ��+��J?�� g`����
�,��$���N����?˻o��:�ZIMg�       8Rҥ�k�FJ�� ��-��O�[��O�:Hv�m3|�?}�m 8��A�LR�k       h��f�~^J/;�� ���2Upo�+�,�OOfk�|�?}�ݓÅ�~Q��       �e�ھ�~^L͠u Xi�䎂{#�+���z5yu����Ƿ���͓�ܔ���w��        TRR3H/��˵����E�Ђ{+$�Z���]$W�H������RX����њ;       �nJ�Ԍ�ύt�j �� C��>��Βzu2[s�L_���~�O�`��e�       �DIM� ]���)鷎 k�0�;
���0�N[����J����=��[w��o���.գ5�Q��:       pN%���˕�r5�� ��{��;lC�ɝ��)��v�����<�7��7��燁�V�O�VJz��        gRR3H�(�\O�%.G��&��o�����u8ޫ��	�_��__���()�[s      ��h��f+�\7l Tr��5R���a��:<[W��,��ӽ��������$�dJ�鬹      ��*�G��Az��^vc� m:Mܛ�&���:o��\.����o��w��������       �GI/%������+� �@�}Y���ux�O����^-��?|e1+���.��ZG      ���h�}ve�I�����u, �S����~��u
8^-ɧ�����������VN9����/�       p�Jj�G��]z��.;IJ�` �aܗ�M+�,��^��p���_�^�����>(���.5���d       X���$�f�^^8��� ��Sp_*�?L��C�	^'�9�j|������H���;       ,T�h�=�鲕^����@K
��d�0���:<_-�g��+=�N����ksx$XO%55cg�      ��}|�����k��: l�����y�A�p�I/yat����k?�;o�s���VR28�%��:       ������j{I�0�\OI�u0  I�T�}��ڛ-�ò{e����=���_�O�5]Ʃe>�P       ��R�;��z���^v�˕���2Qp_:�$<l�NVJ�[��=�/�ǯ�/l��~�l�I       ���fx��^R�K/�S3n x���RzO��1�fK�����_�?��w�cv���IJ.x)       X[%5����YM��$�\���`IMg{�
����Aro�u
8��d�����������)�R3��ٻ�/7��L���V��[S�%Q�BJ������s&��fs��$�x��q��z���g/�VR;�&�Q�A�Z�4	���~���j�QO5��O�~       n;��>J����f��i����� ��+�-+�9���o��o/&l��a�L�.      `˕��S2��"{�(���> ��.�4Qp_Io$G]�)��j������_�:���/�RM�qjv��       l��6%���+)is*m�DM ��Ԃ���&y׊;k�� 97z��~��\h�f%m�L��      �-RS3J�����i�?� �Ç��
�+ꪂ;k���d���q���^|�j%5�ԌS��<       ��f��Q��5��~J�� ���w�0�~�w
xp�$'I��c^�ի��O��L��J��Lf����o&       ���k��$���l��� xh���zx��p2�M��=���/�M������+��8w�R       먤�f��aՌ2���� �zRp_o$G����'v��]z�����^n`���njvS��      ��Jڔ��4w|����9U8 Xw
�ka�䝛}���{f�ԏuh�|�������@@��_�k&ޱ      ��(���d��1�V3L����/ 07�����r�w8�aM��c����d:uK�_I�(5�;��       ����f0[m�w|<i2I��)�o �A��ƍ���a�)�����w�D�|��0�'�4����^��x       X��fVlo?��6m��d�O0 `����՛}'����8��ʫW���i�q�OQ2H�IJ��0       ,TM�hv��cmMv3ȹ�����M��V�>H���?VMS����_�F�S�İ�JjF��}       =(��f��Wڎ��l���;�������4�;V�YS�6��o����(iR3��0pR       ��;�V=L>e��f�A�ݕ ����ڹr�wx8��8��~���;p%��L��      ��)�����_m/is&m�|�� �M��vn%��N�G?�E�}�3)�4������ԌS�\       `nJj�ZlO��aڜ��} �]���U+����f��8��\�Q��p|+���ā7�       ����A�����5����Sis� l��r{��V޹�ܜ���;�n�'���$�SO��do��D��*�f����(       ������l����jǫ����-��ྶ�$o��;<����~��K)yҶM���GQRR���ݔ��      ����R2ʧU�J�&��j��� ����ڕ�d���q�
���|�#�<�y��'{J�KI����q�|g=       �4�&w�Sx� m��d��` �
�~�����4y�V�)���~�f���?���O����������a�Lf��      �$��ͮ%�k��\�]�� �v�,���+}'�������]����ǳ;-1�8%5�4'n      ��Jj���z-���� |
����ar���pw]�?������K)y���i?�`s4i2N�(��      `[Դ�b��ٛ�3�� |*��pՊ;+��;���������h��XR"`Yj�i2��j      �MVRg��A�6�V�d�si�w��  �n��Rp_So$���}��w����t�ϟ^p`�JjF���^��      `=���|߽��d7��d��p ���,�o�i�K�j�$�{_~��?��g2ڱ������njv�]�       �$)igw������j��49׋�{�������ؕ�������ֵ���~���Z����R�_f`S���ٛݖ��u      �uTҤd4[c����W� �W>����nN��n��>���ɉ?gww��.<��4��8~�05�{��      ��RRS3���^7�� <�.G������{�F�	�C]������>��'�f���9'V���4'i��      �]��R2����Zm ���s�0�~�w
8�ڕ�����П�̳����h����դ�njv��      �j)iS3J�s�n�� ����7ӕ�}'�c�����k-y��Si?�`;���d<{��       }:�+�(%�����v `J�����x� �����T�.�������<;;�<���sH����Qj�)���       �PS3L�(���Ym �ɂ���\��N�~��;y��+sy�3g���g��\��8^+�      ,MI� 5����Zm �O�}c]�q��}��W�~����3�g��;���CI�����Ļ�      �������ڬ�v `Q�L?�1�q�%�Xq�'G]�����\�����/=������뢤d�&�Ԍ�      �1��=J� R�� ,�����A�	�V����y�������A��^x2�x�/l���a�LR�/       ��>L�(R�� ,ڧ��'
���Q�ޭ�S������]�s��ɧ�/���uQS���qJ���       ��������`�[���� K��޼�w�������z��<����N-��z(iR3N�n��      ���65���]�f�si��� ��)�o����G}�`���������Yq��d��]����6MƳ1N�       ��x<l��A�j����s�� X��S?�ཱྀ���L��Z�q����KO�VEVඒ�aj&)�6       ����>̃V�ji�o� X�N�}{�}3����0W��|��^��vwG��ܓK;�JJjv�     ��u|�t�z�b��j�$mι�
 �D�}�\=�;�����W9:<\�1���c��]�1��PRgE�qJ���       ,�q��d'I�]`?^m?�&��� ���O������r#9��75��|����q/\|<���^����fVt�Iq�<      `C���%'X_/)isj��n8 �S�΂�v�&yˊ;t��(������إ�<��Si[�hwSR2H�dvBG�      �ǣ_��r�k�5ô�O�QA �w+�'
��̓djŝ���-]��7�p���KO��U�^JJ�i2Iɰ�0       ��Ί�Ü��UR��tڜ�� ���]�D�}�N�wn���M�ǿ��#d��8�yj���Z(��f�r���      ���f8�{���^5;d?5;�� ��,�o�7n��_?<�w��̏��O}�H�<����=w����(��ٝ�r��       `���R3LN��^�d��is:�� ���྽�����3g���;�G<����������6MƳ�/�      �Ur��>J�&)'��&�����B� ̇��V{�F�	�4�{_�;�G�Z���iۓ�[�v%%�Y����      ���f��~�b{I�A��d�ğ �|�]�D�k\;L>8�;���;��������	�a�.?�R���TI����;      �r��Ԍf��'�t�$M&���v!�  歳�����N����w~�w��������������E�=��      ���b���u�f�6��d2�p  �ł;y�0�~�w
�]����_��{�l�?v���Z+���ĺ      �����C�KjڜN��)i� `��ޞ(�o�7o���u�ڛ�巿|����̳Od�Ը��ګ��M��B      �\���f����Y��A�S�3�p  K2��z{��U޾�Xq����~�w�RJ�s/<����20MjƩ�x�      <������!�$]�d��is:j_ �z�w��+�-��A�	XW�.������c<�����/���w`C���w�%      �`JJ�Ԍ������8��d8�t  ����O�����ɭ{O����o���7��;Ɖ�ǣ<���}� 6��ɧ&��	(o�      >]M��QJy�k�5���O���~ �Uӥ��+�o�i�+V�y_������PΞ;�'>s����))��D�      ��2+�'�<�Ē�6���\�C.� �.�|̕V�9��i������c<���y<��L��l����NN      믤�ۇy�ZV�N�O���� ��.�Ă;gŝ���_��k�]�;�#y2���X%5#Ew      �B���aJFy�:VI�AΥ��Gz ��v�r{��ֺr#9���$I��o��5M���N���,���xVt      6ם��桟�$i2� �R2�[: �Ut��~o��[ʊ;��Q�?���c.vv�y���)Ų2�hǷ����;      0G���#ۓ�f�6��dw� ���}���޴���ן��Û�}ǘ�S��y���}� �DI���٢����      �VS3x����$��tڜu- �2�//+�o�i�\���}|��w���̓�9����ViR3N�n�D      �\%%%���9����n9���G �f�L���-���Ȋ;wqpk������;�B\|��L�v��l��6MƩG�      V]��b{I��<ҳմ�\��z�� XO]����Yq�~��O7��w@�Z���3��l��fVt�M�r      V�q��f�̡�^R�f/m�S��  l�.�Iը"o�H6���#�������Pm��/�i�(�QҦΊ�^�     @����|��IR��A���� ����^M*r����;S�j>�q��}�}�X���a^��tJq�/�/�'�Ew      �ɇ����G����\ڜ�k�  �:wN�u+�|���#,�ީq�y���c [�v�}���x�      ���b{I���?{N  n+9��#����4�z�w
V��ޗ���T�;�'>s�� I�����>J�r      ��v�}8�b{�����Ԍ��|  ���;����Ȋ;I�~� ��ß�c�~���?�w��)�f<+���      l��.�ϧ:U�f�sisڀ �=t�oQY���:ꬸs����}G�����x��w�;�Y��x�}^�      �MJ�;����VR�d�A�͞ ��9^o�w��Sp�Ӽa�}�uI��?�e�1zSk����p���c���ͬ�n�      ���b�0�J��f?M&1R � �� w>Ɋ;W޾����_��W�A�K/=���#XE]tWt     �OZT���� g��lJ��=/ ���r� �*
�|:+�����i�V���0�_z:�(��J�      >nq���&��?{n  N�A�;w>����%������c��S��y��'��p��      ��b{�����4�$�� <�Z�Vp�o�7�|���㕾c�����O��;�Pt     `�,��^�f�sis:E�
 ��t��^ܹ��.�b�}���o�C�V҅�O��ٽ�c < Ew      6�b��%m�2�~Js}n �mt\n����q#9���%gA4    IDAT�]�?����;��z��'��;�;�	(�     �yYlO���r>5�?7 ��:z��w�m�%oZq����^^��}�XYMSs��۾� ��ǋ�^�     �~_ld���9��� �n���)�sWn$���o�o}�G}GXy�A��/_H���	���E�qjv�e       ����]h������9��w  ��=p�=
���4�7�N��M���K}�X��(/\~:��. k��d�&Ew      Vև��ASlO��f���f  ,�у>�$)M�ו������XG���N��v��kc��8�>�d�1 �q�}���$M�q      �z��wf��Ō����|��Z�1  ��K����w�y o���E���~�w��sn�T���X�1 ���$�Ew/     X������)��4is&mΦ� X����ۓ$�rs���y� �a�}#M������c���<��ǟ8�w��9.�OR3vB     �%��؞�Y\����$��ώ ��LO��&G{
�<�ׯ���E��+o孫��cm]��DΞ;�w��*iR3��۾�      �q�ؾ�Eۏ���6��d���  ���3�h,��޹�\;Lƾk6�׿��}GX{Ͻ�d���{���0W%MJv��(]N|�       �SI��Ix�哚A��2� л��k��wN�}'`��]����c��RJ^��tvv���L�     xe��^2ʢ��%5mN��9׶  zםx�}�鞂;'�����þS0/��͛y���������ҋ2���\�E��4�Kɰ�8      ���b�pI����$��O��B� ����%�N�9%���ɽz��j���������Q��6�^z&M�G+��JjFi���Q�O     ����Ѭ��,�x5��9�&��v �J�N�]��;'w�(y�f�)xTG�.��}��ggg�K/^H�~a�AI�0M&��      �Ql&Y|-��� ���L���  �L��?���Sp硼z#��q_k���7r��}��H���<��S)E��-�Ew     �-R�^l/�is:m�S2X��  xX'_p/�w�ͣ�-+�k���{}G�hg���������d�E��IjvR�p�     �����.��^�d�AΧfg�� ��<̂�4ł;���ɑ��t4���?��cl��?�'���;@JJ�+���      6H��wf��˩����4�K�Q `L���h\�M���a[vɕ��	o�];���7s��A�1������\��n�Q zQ2H�A����t9�;      ���I�ܺQ� MN�,��  <�.G��#�<�7�'�N~� z����]�����>�S��}� �UI���Ԍ�|     X+55�Ԍ��r{I�6����K  k�a�%E��G3M�ƍ�SpG]�g��}��*��<���G}G���{�IJ�q�H     ��TRS3��^�d�A�S���� 0o��ݥSp��]9H�.,�o~{5�޻�w���45�^���h�w�QS3J�IjF)�     `�R2J�,�I��r>M&1� �κtYp��;��������?�;���\����n�𡒒ajƩ�Qt     �II;�^3L�|ͦf�6����ҏ ��u�t��%E���x�V��a�)��i�|�}��[m8<.�J� UR2��wS��     ��Jj�b� �^M�i3�ٴ9�� �F9z���w�����^�巯������w��7r�i?�>���AƩ;�	     � %uVl%i��b{IM��i�?[� `�t�PpO��v%ss�0y�f�)���|�G}G`fww�K/=�Z�{� `��4���$%�%�V     �<���aJo���&�r>5;K=6  ��e��],�3_�^O�f�WR��O��W���&���p�BJQ�����Qj&����     ����hVl_�tK�&��|�L��b=  �Ui�=
����ir��|���|/o�z��|̩��<�)%w�RS2��wRz8�
     �>JJ��u�a�~jB5��9�&�z�  ��t��Ѷ�-�� ��Hn=ʝX��~�}G�.Μ����>�w�5RR2H�85㔴}     X!%5��b� }���2ȹ�9c� `�<�z{�N����v�7�N���$���_�;���t.\|�� k��v����(�     [�Ί�;I��Ul/i��tڜ�� �&�#�3�b!�$��d�pWo}���굾cp�?q6�n��W��`�Ԕ�K��V���<�͎      �AI3�w粤��$5���  �o�G}��w���}'����?�������g����JJJ�i���Q�>�     �%%mjvR2L��DJJ��3�y�v ���=�{I�,�{���o%{�6ջ?��/���p�孫��`���2M���r�w$     �GTS�$i��^��$5����  I�ܞ$]�xu�B�r=���宾{=����}����}�ɜ>3�;�8�9>�:Nɰ�S�      'WRS3����M����QڜO�S��  �N��<��z��B�8J���b����~�wB)%�_z:{��}G��E�Qj&����     +����F�(ǫ���f�sis&e�  �Z�sXp��;�����Ќ{o����U�xH���p���G}G�05%�Y�}��W     `Ŕ����d���BzM�AΦ�ٔ�� �ʚK����0�K޸�w�����ן���<������3�����n���8%m߁     ��VS3H�άD����I��i�?+� ���2M2�El�,Ǜ7�syS'�(�o��mr��g2*^,N���4ٛ��-}     �DI��QjFɊ���e����;  kanEaw���}'�>�G_�;s2�y�s�*�,\I�(M�f'k�\     ���fG��ո&QR�d�AK͸�8  ��n~�f5^�޿��{�����ͣ��{��w�h8ls��3(�,C� M&����Z
     ��Jjj�b� �SlO��f��i�w� ��sy�΂;����d���b;��g��;0����������i2�-�8�     �����QJFIڬ����QڜO�SY��=  릛ۂ{Qpg����}��_��������F�\��3J� KWS3J�^jvR��     Xi5%��>̪��kFd?mθ� �#�O�}F���{�Frk>w!�.��]��g��;��3̥�.�m�d X���d��q��S�G     ��jj�b� �Wlf�s�b��  <�y���4��y>!��Q��v����׿����������r�g�4�u2`�4�ٝ����J�     ������v��`q�f�AΦ��Y�  ��\��k��;=x� �������I�X��x�˟���г���a�LR��6�     �%������aVm�=IJڴ9�6�f `��t�k)��ө�;����7��uI���_�;K4[rX�Ob��dl�     6TIM� %;���w�ג&mNg����� �5���$��i7�1�7���ܙ��o_�k/��w�l2�ɥ/���;i�������l�Ū;     ��;��GIھ}���6�2�y�v  n���Ird��^�z=9��7�ۏ~���#Г��n.��;��))�f75�=�     |��k����A�ռ�vIM�ɬؾ�w  ���sd���u�k7�N�Y��O��wz4����-�����fVt��N��y     ���y�;��W��q��b{�IV5'  ���Ѽ�rZ�Sw�u� �>��l�kG����K�1�٩�c%w�WRg���즤�;     ������k�ɝ���� ��Q��Wяj��N������B?�ٯ�����]r/�	��VRҦf�&�ىr?�    `َ��Õ_kOn�w�Zl �gXoO�i�v������탾S��������r��8�_zJ�`m�Ԍ�d/%;V�    `�Jj��Z�(Y�s�-��JY�uy  �Âv֧��)��^���n|hG�.�����s��^�{�I%w�5s|��q����    ���^k�%$+^/�b;  +iQ��t���<��a��v=�0�;�z���Wr�歾c��Ξ;��K~���뼋`�4�i���V�.�     �p����wP]��xIR����R;  +�x�}!5����N�YW�s�d���d�����I�Xa��O��������JJ��5��Ls�.����     �Vgc2�SDPl `=,l�q�N�΂;+��kɋ��a��tI���_�;+��SI��֟Uw     ���[kO�{%;i2�e �յ��ʴ�Y17����Ϗ�N�>��u-o��f�1XgϝJ�5��o�UrX{V�    ��o�=Ql `=u9\��dZ�S׮'�|g>����}G`��>3���N�� �9�Ԍ�d���+    `���׌R3ʺ��kFis>mN+� �6���3��%7k������au�+��N�>�����;k��~A�`㔔R3I��l���z     6OIM� 5�����i��AΧ��v  ��B��uV����έ��[}�X}�����c��N�+�l�;W�GN�    ��JJJ��y��k��s��$��b{c� �5���yIn�N������t1w0����o���;uz��/=����JJ���Zu    `��S���A�m��v�������  l�E�ϻ�v�.�����7�N�ھ����57���嗞IӬ�I  N�|d�}�	t     VXM������;��� �f:J����rP��ӛ<<�7����i�|���;`���K/^Pr��o�:���GY��     6Q��X���6�x��$i��� �F�.p�=I�t���}lV�4�o���b5�q������}�`CL�vsɒ;��)Ί�㔴}    `˔���������b�cirJ� ����p��_���iwc�G�9x�0y˽>�'?�E��0��N.�b�։�mt�������v��y    �uPR��J���Kߡ�'��ί ���OW/����H����ʵ�p�'�̗��;}G`�ǣ\z�%w�-v��s���d<[�    �Gw�Z{2�:����v  �J�i�K�<F�Y�Sw��Q��r�����p���?��5����.f0h��@�ԌRs*5�n�
    �C�)�֞�.��3�y�v  ���P��:=���6޾���������t�b��v����g�Qr ��e�����͖u��    ���W�=�2JY���v�}2+��eݿ  8�.��8�A�v�K8���ד�^w��[?�;[@��OSRR2L�qj�)f��v     ����AJvg�׿^Rg����d�M��  ��tKXp�Rj���st�(y�F�)��%����f�1�;;ü����������&��줤�;     KVRgw�� ��Kj����'1� �6[F�=IJr�����r4���o$7���d%���ʕ�c�EF�A^�ܳ�}G`e��R�Xu/l     6������ ��l^Ҥͩr>5�(� @��p)�))�2h�]��`�^�v�d����_~�w��p����]����( ��۫�w�ݝ�    �%55��]=�I�l�9��6mNϊ�ٔ�  �aY�.��i�YK���}��Ƿ����#���6/}�b&{�}G`-�;��{��Mِ��    l���65����;�[3H�3d?5;}� �4Ͳf����p���R�������5풿�����-�45�_z&�N����)������>JI�w,     ����QJIjߡ��v��͹Ը�5  �Ͳ�ۓ���_ǧ�o-�0g�$/�w��z��{�~mK��Y��\z�BΜ��;
 k���d��q��g��u�W    �UPRS3��ڇٴR{�Ԍ2�9�v  x@]��v�i�A={�w�����[[�����?}G�$I)%�_z*��O���v���d��ݔ�Qv    X����G���-Ijv2�~ڜ�-�  ��-��^3����\߬_I�F�\O��`��8�	_����� �SJɳ�?���y������Z+)ig�.]���RA   �N]�����ir�о��KJjvR3NI�w  X;�ݍ�'�R�ok��n��c�Bu�+גg��N�X�G]��7?�;|�O��y��7���F()��s��r�in%�   ����æ:�{��ln�=�����d7��� �"-{��(僶�ڑ	w6�;��wo%�7�.b/��V�G�]���<��Zk^���}G`�Ԕ�d�.�t���V:�X    ��R����.���4�f7��� �r.�hM�m��@7�M��d|:i7�w���g}G�{z������׿|��( l��0��we��t��w,   ��"2��K�M���]Ҥ�$5�l��  �ѥ�r���r��� y�Y�aaq��+ד�㾓,�W��w�� �u��3���W��j���o ���II�.�$��r+ݒ�1   �ٜ�u�m��$)ig��;}G ���Gc��A����N���A�ޭ�S�ߍ[G������@�����N��q����_���M��Ԍfo    x4.!ú()���]0�lC��f�6g2Ⱦr;  ,H�������R�7��:d��|-9ڰsn��͕�#���>3ɥ/�ij�Q �%%�Ԍ�d��QJ��   ����a���ߕ�wR2H��|hIR��A���\jF}G �֥����o�$�~���e��4y�z�)��~`����wj�˟���������S3��g�m��   0��JJ�ٹ�Q�%����W��6���tJھ# ���2���$��tnݼ�aU`H�$�-��#���/�m�ࡌǣ�����d�%5%�4��{�в;   �=�t���R�`��>L�=�R%5M�2�cir*e��v  �[��>�v2+��<��A	`�^��m�����4����;<���a.�bF�A�Q �r%55�ԌS3�]Rv   �(w����Ajvg�1�$��XKSҦ��r>M�٦�  VE���[���� ��4yu�O���W�� �l4���]��x�w ȇ��͖�ǳ[ںH   �e�`}Xj�I�(ǥ��R3H�3d?5;q�  �2Mo���,�����$W��n�����Ï�w�`.�6/}�ٜ:=�;
 |�q�}75{��G�w�   �C�aY>�Ծ]�f�AΥ͹�� ����ޞzg�}zx�v/)`I~s-9Z㡉o|�{}G�����ҋrn�T�Q �J�2��o������   ��:wX�K�-�'��9N����_��7�4�����ȅ��M"��J%�IU�3������\�5�ƀߘo|1��x�3g���}z��T��Z�DR�H�{F<���"���d2r�~ �df�$R̈���a�@��$I�$��
�G�[(׳��וL!��nK�pmK���9?���U�!�T���\�9�`i�U��H�t�@�V�#���6�\�[�$I�$�4�R�)EaR�8�*�mRZ�c�_�$I|���{H��M!��כ0]��!����қ�G�����9�4����U�"I�g�w�7��$I�$i��<$����%�Hh���`�$I�4����ʲ�P�����������5�=��+����R�R_]�<K�����yn@P�4�z�\�awI�$I�4�lp�N�P��e��Q�(�$I�����#a����ip�X��aq�jW=������e�#H}7{a�4Mypo�,�$i�v�V=�$I�$IҩDr��K'b��c�@�	���F�$IҰ�2�������M"��7���]����"����W=�t.������:�z��Q$I:�"��"e��	�k�%I�$I��Hu-m�0)B�u����RjLRg��)��$IҐ�~����=H��M��H���*t��$���b�!C��jr���4'\�P�4슰{�/�����$I�$I�>��eȥAHH��ڃ��]	5jLSg��6�$I��S���?��D�+�F:g�kUO�y���G��]�Y����iw&�E�B�'    IDAT������!�e�]�$I�$�*�!���P�M�JhP�5.��ZJ�$IfU_�)2�	��w���mx�U���˿���G�*Q��ܺs��NգH��c�@��	���%I�$I����D�4�Z �Ң�5f	ԫI�$IR��g/�����U��HYX��j������z�2I��/����zI��"�!a���%I�$IRu"pט��Oj?B ��u�I�"�V=�$I���U��*�+(��n������]�L���#<Y-������_�z�R!����+_�U=�$I}�vo��!�]�v�$I�$I�'��y3�_�!�v���Р�u�Hh៑$I�4� ��~��� ���V'&����$Uc��7a�Y�$zp�Y�#H���9�4����U�"I�9(�-ڏ"��H�ܑ��$I�$I�H��R�	�H1�}��Oj�\y���H�$Ir9�Ix����^����
`�]cii:5���~��?U=�4P.]��Ѩ���"yn�$i\��7��P�ݣ˅K�$I��3�ѴjO)�7��)����M�$IҘ�ca7���|������a�����5j�ſ����zi���N��k�i��;K�4��qڤtHh�'�$I�$I��n0NfK�����$a�@�?-�A�Y�̑��?+I�$i��1����G�	�n����;K�a��׫�������Ϗ�CH�Smn�p�f�^�(�$Ul�}�<QW�O�$I�$�4"Y�z�4�		�2��$Pg_$B�(֏lQ�"5fIhT=�$I��J�AYE���<���E�7`u .BYXtA�S&&�����VգH�4 �:	��ٽe�]�$I�$��`4�I'�?�h5�^ %�C�9R��c��$I����7������"�'k��jg���T;�4j��[w���ũ�G�$i��r��V���&� v�$I�$I�ٮz����"�>a���Ԙ-���s�$I��p�kp߽��j?�di�le��_�����SuO.�7��Js���«�Ǒ$i R)�,�����b�$I�$i@p��Je��d[�p�@�DY��V=�$I���(??�_����j��ϛM���L���;����������ru�z�ƓGω��%$I`�hh 9�l_��ߡ�$I�$������48��XɾP�N*)WyL���$I�$%��@ ���x7��lՖ���OOנU��9/Y~������>�4��gh4�<��@��U�#I�H$��\�]ݷ=�-I�$IҘ��]� |h7�~4Ii���$I�$�s��n���^a��y5�H�)��d���Ky�����$�PS�mn}�F���;K��}�	M&Ii��,��$I�$IҨ��d��F ��P'a�@����cR'HI�Pg�3��%I�$S,��C8,��l�1��'�څW������_��	��j5���Z�fգH�4�R:�[�lϒ$I�$I�'ݪ�И(Z�w�&4(B��цRB��ԙ#��H�$I:�H��>Z��g;����/!t7V׷�I\��a�/P������=�4���������dգH�4􊓎ڤL��"� x�Q�$I�����=@��5�I���$�,��b�V�{ߦ�5fI��z$I�$IC*���^���;�|�׸���z��H�-�B~G��2��o�����1�$����ʥ˳U�"I�	��:��Ih���$I�$��h�"���([ڛ-���"�F�)�̓2銋�$I��(9����[��Im�'�[o��:�463XZ�/��}��˫loyQ�׮_��l���1�A#IR� %��� r"��]�-I�$I���lW=�F@ �2tm��W���rU��� I�$I�T��)O��w��_ߜ�<Ґx�	�u����9>xֿ�Kc���Y&&<��@��U�#I҈J$��.�����%I�$ID9[ā:����cAE��P{o�����V�$IR?���@��{BY�K�;�4\���V�9����۸4榦����:����$�[`�$\��	�.�,I�$IҀ��������Hh��z�z�{! 	Mj�Rg����J�$I�X6�����{�$�wi�d��oQ�_��O}ڲ$�V���n�j7�E���R��l��&e��vy�t�$I�$U'�+�IG)Z��e��I��ql�B %�C�yj̐Шz$I�$I#��܊nG�;�?��,��Y���ow;�����R���5nݹ��t��Q$IS�v�t�ݽ�'F%I�$I:?9[��;����7wC���m�$I��4������Of�/��|Ǒ�ӳu�Ԋ�^y��������!��4M���5^�|�u��H�4�v�"�����t�H^�h�$I�$���V�#h �r������(~� ���vI�$I���2���z��8;�y���d���Z���<~��7�t,!��6O�����%�ܖI��W��R�Yܻ�t��\"M�$I��!�ٮzUd/оjW? �$�E�Q�8�$I��\N� �{�d��z੻S��l尰7:�����no6$�D.\��Ѩ���"�ۃwe�$I�8�� �Q�^gD�D2�˳%I�$I:���<������
��K�$IL�y�{J����{Qu1,oll�iy^o�f[���ߛI:��d��?ܠ�nV=�$I:B�t���$�M�$I�z<)+I�$I҉����XBB��&	Ͳ9�����
@B��ԙ#���vI�$I�#��rgs�����=������oi�-���޳��w�J�F����`fv��Q$Iұ��$m��vy��2I�$I�>%�M$�z�\R+i�0AB�"О౒�K�Qc�:��1CB��$I�$�#�.�n�죀����sG9�x������6k=�I��$I����ʗsU�"I�N$ )�	mR:$��v����$I�$I(9���\�nK{����-�\��EZ�g/I�$i�E���(��P;x����p�\ƑF�fkp�s�ǿx��ہ$�ɕ�sLL4x�`�<�+�$I�'����99] +�[���$I�$i<E�A>���$M�)�t��$�Hh�0��vI�$I�"���'£��}p������#���[Щ�������R��t&��h4<�����n��H��3I,]�#݁݁�$I�$�"�^�=TB�V�SW%��0AB�%I�$�����C�?���1�����#���5X?E>��x��Y$�]����7hw&�E�$�TJ�AB��)���II�$I҈�٬z}B(W�K��a�&�:�1��UHhPc�:�Ln�$I�4�r���H�8��_]����#��x�
�	�/��W��<�ή^�q���\���zI����MRڤL�M\\�[�$I�4J"[D���B�^/���1�ګHI���<5fI8�ޒ$I�4P��m0⣃����l5�.�tz[<]���ݿ����|��CI:�7��Bs���ӗU�#I��*��M '����A I�$I���بz�H�&p/�ť$L����$I�4:r���r�G��C����!��-xU��c\��~}��-�a�ŕ��ZM�_$��I�4vN:4�D��{F$��$I�$�H�H��1�҇av탦h�/���K�$I]Y�|R��G��A�����nwM�Ig��k�8N�����#�g�g:���:ͦ��$��P��n��"e��v���K�K�$I�Wn{��)��Hh�m�M��9��"��Ҧ�5.����:�$I�FU,W-`�����?ڋ!ĵw���g&itE��*t?S����ҹ�#�wZ�&����T��Q$IR��#�iՃI�$I�P�B�U�#��@{���HhRc�:�Lz�F�$I�X�lW=��|��G\&�������H�a+��k��ϟ~w�|���S�Z�w��17?S�(�$i���ۤL�{R[�$I�t�r6�L�Nd'�^'�Y��hT	5jLQ�5fHhT=�$I�$����Gx|���n���~
|�׉�1���j0�<�����w I=B���/�L�x��y�)I�tPJ(C���ߺ�p��$I�$i$䶷�YB H`�M�,��0Q6���.I�$i|�;��hp?4��gݿ �s_'�����Rh����p���JR�\��f����ݧlmu�G�$�P��wN��w����%I�$IꝜ́?�=x����Y�mi�$I�$(���C��'����wi�D��*t?\Y�$�b�FA���Ώ7��jW=�$Ia��=�M�T��Y�.I�$I�YDr6�b$j$��pt�\�������Р�4u�1m�]�$I�vE`��!>+����ō/~��q����U�9�w���o�HR��j)�ݾ���+�/��zI�4d�@{
e轐��a�$I�$�r6lo?�N3�^C����@Z^��*�%I�$IE���@$�����i����iIg��/7`~������j��s!��6O�����%��_��$�,������]"9�%I�$I���}����HHh���Cc�$I��}"ݪG8��v��{~?����=��z�˝�[Z�v�x��?�s)i\�8Es���{ln�R/�$i8�2�N��^�ܻe�=�*Ǔ$I�$��mo�GC Ͳ��Y�8�$I�4DbY�6�6����þph�=���{���ߙ���ǫЍ���s��H�v���n05ݮzI�4�	�	-R:$t�&��V=�$I�$���ޞHI����MMu��b���(�A�i�\�ƌ�vI�$I:����>���#��޽_��4Ҹ���Ờ�??�zI}V��|{���\�zI�4��{��&)�2�^ރ'�%I�$i,�r{{��~0�ޠX�ܶ�aHI�Pg��$L�ߧ$I�$�N>4�x隷Ԏ�����=����#�{�����+f/LU=��>!��y��&�,��ybA�$�d7�^�Y�.'����D�$I�FǨ�����&`=���	&���$I�$�E����'���������H<���G�hN4h�\VO���h5�w�͍��Ǒ$Ic)�0މDr��v/�K�$I��Ѱ��a������"��,C���Ǒ$I���S܇C�#��Q_����؟q$<��c�<���Y6W�H:���w~����dգH�$;�	-�$L��"�(C�$I���Y{{fO��<7):�vB���
Mj�Pg��)��$I��q����Q_;2�>=5����#	�ɽ' lnn���1o����Iӄo������E�$�#�ly/�mR�Hi��,�ߏ<� I�$I�P�����'��f���r?�����GMB��ԹD����,I�$I�S������"���Q_H���,j����ݧ��[Yci�5W���p"I��+i��<���J�$i���}��s"�Ȉ�ZF�$I��T�mV=ƮPvv�}�8(�'�0��$I�t�"�U�p"M�{�G|��=�.�w����(�4b��}����_��ͻ���T��w~��D�Y�(�$I'�vOXwH�$����66I�$I:O9k���n;{���8�ήQHI�Pg�Hh�߻$I�$���,(/_�+G}�{�+��/{?���.K��}t�����ت`"IUj6����:���E�$�B��� �U�;$�4�D�$I�$�Kd���B�X�ٛ���Mu������̑�q�_�$I�*t��z�ާ��ɀ�����O}]��,<xJ���J�,˹w�,�+�JR��4��o�r�����I�4�����$�I�*C�E˻'�%I�$�72�������#��=�=.���6u.R碡vI�$I(ݪ8�@<}�=���ގ#	��ݧG~msc�G��qI�dn~��?ܠ٬W=�$IR������O�7��I�$I҉�l�x���v��}��)�@BJ�:ʦ��r^�$I�4("]"�V�����~2�>;w��vI ��~zq���y������4h��&w~��셩�G�$I�P��7Ih���	-�����$I�$.'g��O��[$4�vv��C��L�9H�$I�Qd��N�O���'/���4�O��N#	��}���,>}I��dz�sI4i����Wy����/dI�4	E�b�E�6�x��#I�$I�-c�x�}�@���J�����_ ���o�]�$I��G$ҭz��lp�d�=l��辫�s��pxx�;?ޤ��QW�.��n7ypo����{!"I��{���2b�V��*�M�$I��钳y�WÁ@�av��Ni���f��H�$I�NaH��Ii|2���u���/³��kG�tJ����X�˲��w�s�	�q֙l��/n25ݮzI���h��"�M�$)mͲ����$I��ѕ�Z~���	�}�Ͳ�;��#�$LPc�:��1m�]�$I��ؐ�_�+���'� �o��z7����^?{}���o���?�Ҹ��R��u�+_�U=�$IҀ�	u��"�>IB���Ҫ��$I��3R"]�n�=��a�Ϟ��
$���s�P�$I�t@�;r֫C:�b���1N�O��C�sw�\���ٓq$��/���d��o^��՞���4��aB���9&'[<����v��$I�\(C�龾�X�Ɉd��YUJ�$I����bf�}�K�=�8ͫ1��"���_�$I�A9[d��P�,�!mo�g�ǹ���=�DR�񽧧z��ӗ�[Y��4����T��?ܠ3٪zI��!vP&�Hh�M���%I�$��P�$��)W���!��Y�d5J'6�ϓ2e�]�$I:RN�
 �l)��L$2���ϟ��g���_��_z3�$��S�c�<�����^q#�����|��+�E�$i5-R:�L��.��e(^�$I��&����E�=)��f�or��G�:��6��_))m�\4�.I�$�@��r��B^/+֐(�ۇ��5�g�?�v��t�'/J�zg�����f<�����o�$F+�qB��k�t:<z�D���$I��) �G���@g���&��<p$I�$��);�H�	����HN��^��!V4�O��0�.I�$�Bq��G�G�tY��LSI'��"����?Os���51'�������6y�p�G�H3��|���iw&�E�$i��ݶ��)�$t��ŝ�Ŵ�1%I�$��P^�(���$L��[��B�6����ŵc-�FJ�:sԙ#�c�]�$I:�H��wG~=g���s�H:���kh��[+���ܝ>p��C�޾z�73IZ<C���7������L#iT45nݹ�ܼW�J�$������v|o�0Q�K�$I�a��s����������JPg��E�f��a�P��$u�q���)I�$�^���g/�Xu?L����=�����T;Ζ�/�4����g��[��<��'�z��&��=ٞ��$��7��3��ɣg�m>�$I�	��ˇ�zy٦�ɀX��$I�4X�H	��}�YZ�O'��r�ϩ�¾� �����$I�4�2��l����
���{��ɇ��⟎s�c��u��O��x�q$���s�����91F��]��7��h�d��F�Źiڝ	�_d}ͫI%I�KR�b��bzψ��}���$I��I�2SJ� �����ዡ]r\�P�ڛ$e��P�$I��9[d����H�e�\���$9��y�@��q�w�#3.N���Ƒ��p���˲��w�2lJ���D�;?����٪G�$I�g龖�6)R:$�Hh�� ���$I��U��^+_{O��&aj��w�A�60����/4<	)-��R�5�I��Ќ$I��/��VǊdtY��<��E��ጒ��^�jp��v���Y��zp��������u�<�%iO�k�/39����gt�C�4�$IҘ	�m���[$���$I��g�tZ��w�\�3+�T��@Z^��$P�zI�$i�tyw�ձ����Hi�x*�4�0�+�e��'[���Fó�-�!��ne���_�Ս�}پ��63;I�3��K�[Y�zI�$�Q�9|�D"������$IҨ*B�\��x���0�����H����f�=*I�$�嬓�y�md�')W���}{;�UV�t�;��ο�޿_~��l3I�W��勷�|�oۗ4�������k�/{��$I�H**C�Hh��!e���	u���R�$I&;-��W    IDAT��Mi��yj�B��hܨz�B�g֤�4.Q�	m��$IRE"]2��d[]V�Y�*ꮺU�qVw�/Ǻ��X� �߽<5;���g���p������F��N_�G��ty�hs������_�'I���
e������N��^�{$�U0�$I��ctُ/��R�:�@JB�@��:xQ�$I�4 "]��=�ZN�25f�u��٪z���;�=�}4(�Ώ�QI�[|�����yx���Q��LR�t:���&���E�$I���3�]6�w�ϛef�j%I��[E�=�(_��G���$���p$�H�P�u�H�"���N�$I���x��b��m2��t����i ����=������|�q$lml���۾?O�����S�][�$-M���*7��B�x�]�$I;��l}o��"-�FE�}�@�@�"�.I�$��kˉ݋*�+��E��ݶ�q��I�F�c��ws��4���ER:徑$I��A��A֧���u��t�"�Ğ�GP��x�{�w��8��G���%b<�`67��w�[w�"����vqn�vg���X߬zI�$�@  �!}�ȉ��@�y+�$I����İT"�]�'����!�O %�A�IB��%I�������񮼠��\�L������������c��U:����|���y��9�o~q��+i�LL4����������4!I��Q���Q�)R݋�{�*�����S�$Ig��=����n��'O���򵳪�\m�Q�\�U�$I���tY�{�u,���E�V�%S#Q,������{�c�������������N7�4�.��s�z��D�ɥ˳��ܒ�K��]���T�G��2O�H�$鬊xH ��lO������w�K�$�*�C�;'��%g���+R|����&S$I����H�\�k�)>e�\�O�+�U���3����3'Za��������3IZ|�T��.<yA�Ygz�S��K.3��|���yx����U�#I����6Ĵ�l���=���}���%I��n�"�t7�ďV��y��d�T=�XI�h�M���Ǒ$I��#9�d�o�%c��hv�\�W�$��E��w'����y7�G���t
��ο� ��������:�V��$�F�ƭ;_�l�5K��G�$Icg�1�`�*R����}�^�$I{v.(�	�o�\e��G�
+���@��'4pEI�$i�m��\<��@���z+�ͨ@���_�r�?�ǉ&����j� Y������A��/RI�B���9:��,��=WJ�$i�a�⿇���4����k�$I%;��v.��}嬑��2��hio�д�]�$IU^<�d,S�^>�ފ#u� s���(�>a�W�Ѹ@:wU�67��w�[w�"�J:���6���&�>c����Ǒ$I�>a'ܵ�ٞ������H$��H�$I={����{a�O=J�/�%�c��H�Iʦv[�%I�����Jg��}���J��h�d�J{;@��D��1�_=�ؘhO4N6�4�V޼����T= s�3\��E�cHB�_����3�|t^8I�$I�H$�hz���5�H��q�a��hdO8x�FQ��r\9�,�eK{ÖvI�$iL�l��m�c�1CB��14"r��sV#��;~=w����=���o�^�q����%��gO�U=®W/��h5�ty��Q$��s�t&[<z������Ǒ$I�z(H���젝�����^�$I��>n^�h�x�X5�~
�t7�^F��$I��Y$#c��1>��B�by�A:�H>J�v����	� �k?ܥx��y�#|`����:�3��G�4d��:��|ų��<[|M��YJ�$i$Dg��@^6�!��x�$��@ ���|l�V�l��V�C!v�쁆I�$I�D2Vn�X�U�Bգh�mW=@��?�ޙj�'�ߜ�q�8{�t��1F�[�;��t&�GҐ	!p��S�=Xbsc��$I��������m�������K���R����{v�uz�.+U1�je��AB�$I�$&�=���s��X%��Y�V$g��X��ۓ>���K_^��N�i�Z� �#�.p��4'��@��t&��Ǜ,>}���o�G�$I`Hw�9�Et����{��sv�$IR��o[/>O�[wn3T����|����d7����=I�$I���A�z�c|R�j�"U��Q4��^�qY��t�]��B��tLKO/�������O����4��$�$	\�~��I=Xb{�[�H�$I�P�	������=�X��&xI�>VD����{K�+g����Ǩ\�S���ҪG�$I�4D"]2�U=Ʊd��p�C�uu�3�Ze�'}Љr��+au��[kZ�x��Y�#isc�{yJ���tzS�m���Mff'�E�$IIE�=!�����&	-R�$L�2IB��|�@��(��$��a=P�mAL��*v�߇����	�2D[+���T���dC�臄)�\��%j̐�2�.I�$�"]����%���}A�N�#��[���o��q'opޭ��������4�������c��:�/���W�E���R���K^�Z�ɣg��p�PH�$I�#�؋ �έ����ǒ$��P�fR||x�����GJ�n����6�'��'U�$IR/tyG$�z���$g��VգhH�8>�"��4�;U�=	p��!�r^.��z��z��O�|ym��Q$��s�t&[<z������Ǒ$I���� <ek�ᑣH,C�{ܶ��$�"�>x�?�'��fI�*�}پ6�ih/VVp�I�$I���F�F�c�J��ru9W�ҧp�E���=��Np��k��?O�XiܼX|I��t�/��Ѩ1i��Q$�f�έ;_����^��I�$i���=��Io��D�X5�JҨ�kV/>�k[�k\/�rx��(��I��WR�T'�nHC�$IR�E��x_���d,S�ѧ�lo�Iα����=ۧy�4~�?}^�'�����3��U�"iȅ���E&��<����/$I��Ѵ�>�
6���k��Kҹ8:�{��O��%},���R�=Hv���K�$I:_9]V��HqN��5R:U���Gu�X�{~�5^��ݷ�/�L����8y��Y�#�H�������u:���Ǒ4:�	��x��'/x�r��q$I�$U�` ~����Ax���G��~�C�N+������#>�$v�I}��B�}�2\��uB�&I�$IU(��Y�c�D�jy��X�X>�����o����<�Tw��W���0�W�}�4.��W�;@�G�]��7h4N�τ$�Jӄ�7�`z�����vGc�C�$IR��3o>�,�����E+��!���g�L�(;*��Ӣ~x���� �?2V���������%I�$�g�m��8��P�"�ч"����x�Ǟ��D$�[����ϟ_�`{��ݟ�p����j.5)�7ff'�L�x���o�W=�$I��T���O��~������vn=�$_<&�/��tv�%J��d�q@=qA����&g��1>ɆvI�$I�.g�l���N#���J�dգh����<��ק}���n~�o��봏��Ű�67��w�[w�"����Z�7�}��7�x��m�$I�������s����;��ć_+���+i0|؎w?O��^�z�ξ���q��ey�~���e�݆vI�$I���/W=F�d���g��Gр�G���u�G���EV��2��Ы�ϟo�`��:�/���W�E҈��0Eg�œG�ms�$I�4��/x��{���C��{�����xd���0�4�B�q7��a+:쏝T��x��N"i|uy�����}���+I�$iXD�����]�Q�"MR�p,�O�&�߼;�����7~�zv��lCu��w���7����\��k�U�!iD��.I�$I����	��x@~�c�߿�h����G���N��<^ ��}�{+|G�������4r��R���@����A�̪4�$I�4��,��Y��"�E�T�c�bk���~��_���>�L��-�Y�����}�mH�lcmc$�� ϗ^S�׸ty��Q$���6������Z�8�$I�4B���r��O�`�=��佯|�?*<fg��M6?��-������������4���o�������=��`�������?��+IU�t��)�^��\+��u`�]�$I��X�p;@�:�f�_���e��� �x��)�p����ɳ�G詅'/h4j��NV=��T�����5^�Z����d��.�#I�$I#��0�Y�����A�YK�IE���풨b���@{���$I�4jr���BČ�p?o<�lW=B_�g����o����<^uϞ<�z���1���"��U�"i�]����_|��T��Q$I�$I�$�2���l{���	jLQ�"u.Qc��N��g�A�$I�h�dd,W=F%"9�C��==�0����y���y��{�Vih�Z�;@�G�]`ss���T�F�ƭ;_�Ս�$�'l$I�$I�$��2�ϴ�"�ޢ�4u�3G�4	-���$I��!�L�ۺX�/c�8�M��Xd�����B�g�����eX{���˳lCe/G��c{�˽����=�WI����Y��%I�$I�$�H��w'zL !�IJ�:�4�TڧH� ��iZI�$IL]ލA���uY�1���|�/j�;��3��)�����Og݆4�^,�f�`ss��??%��G�4��:��|���_��.I�$I�$i D��|�a��v��ԙ��)�㝒$I��W�9U�1"kU��s2��D��Y�q�{���ϺiT�\݀;���&w~B�{���������]�$I�$IR�C�v�)j����*�V�$I�Od���U�1P2Vm����^���n���/�]��g݆4�^.�v�`mu���ѐ�����]�$I�$IR�r6��8��}�����$I�t�HF���H+U��>�lf=��I���8s��3�o�����ۑF�˥WU�p.V�Wy�`��1$������x�vg��Q$I�$I�$��@�vvI�$I:�H��ı���\N�����P�D��ho_~ϯ�p֍�9�~;��7��>9�v�Q���e���\i���;��~c���11����׹zm�6wI�$I�$I��{<R�$I�N��2���1Z�*;�GQd���� g�&>s�`su���b;�(y���G����/����7U�!i�����E����LN��G�$I�$I�$I�$I��xO�V�c�H$�]�c�Ƥ����w��N�}1���b;�(y�8�m�O^����4�K�f�[w����/HӞ���$I�$I�$I�$IR�l��V�C#g��ͪ�P����̟N���j��^lG%/��3����s޾�*2I�on~������NV=�$I�$I�$I�$I�؋l��R�C'�=�C=2F����/{�����ե���z���}^.�o�=�ȣK��Uw��_�^����o�R��U�#I�$I�$I�$I�4�"9]��i�B$��~DD��O{;X�7��PO� o^��m��%���K���Ry�w��5�J�T��S��/�an~��Q$I�$I�$I�$I��L$�-q|��=��J$�z�Qd�2�׫�,��h6�m��%���K���#�r�������Y^CҀIӄ�7���[�h4jU�#I�$I�$I�$I�4���ӭz����wU��3�t��"�0x�/o\5�.��rр;@��q�/O���Ŋ��L�t��_|��+�E�$I�$I�$I�$i�e���Wku��l�g9����.�^��_^�w�k۽ڞ4�^pߵ���ݟ��e�t%��A�$�/��s���4'U�#I�$I�$I�$I�4rr6�X�z�����]åc�������?�jc=���K���j{Ұ{�������&w~B���VR�:�-���&W��#�P�8�$I�$I�$I�$I#!�%c��1FN$#g��1tB9[U�p�"��&�{p�nm�u/�'�ՕU�W��r����-�!wI�J����s�����D��H�$I�$I�$I�$�HN��D����h��6��ɪ���^n��������{�=iX�X|Y�key�G��C� h�����:׮_&Ils�$I�$I�$I�$I:�H�[�쾉�2�a��]�����[�i��k�%�r/���{�d��S޼~�U�!I ��ty�;?���g��~�����N-,V�ŝ��Rd�l6�łY;��	r�@�� ri����0;1�x�cE��k��	��#ِ��&�h4�����������y�\�{<���:�w��KW�Z缇d�E����={�K�        ��f�R�Y:�ﵲ�ڏsh%��󴹒�����с��L7V�=~�`'_z�������<���t���޽+.������H        }���T�,�10ZY)��稲U:��o$__����������w�5�׸��b=x�G�Jg ��#G����:��t
       @ת��Vvt��稲�z0�=�N5�W���ӯ���Cǎ��N�&��'�_ԃ{O���|��0::�ӳ�y��S۽�t       @W���f�Kg$WܻW=��f�H�;��;>p߳gϯ��kB��{��tBO��I�>Y(��C�NN���3�>q8�F�t       @qu�ie�t����L5�C�n6����N��;��;>p�7�4�-/,-���B/y����eݽ�8�s�����P#������읜(�       PL�*�,�N]:e����}�z{���|���O����=I�����b��\鄞t���Y�7r����h�x�TN�Ngdd�t       @��ie!u��!�N+U6Jg��ޞ$�юm��}��}����b��|鄞T�u>x�a�WK� |�C����9|d�       ��if)���x���+�.�w�A���\�������v�.�ŕlm�oV����w뾑;�Ն��2s�X.\�����9        m��J���v�:�+�]�5����d�w�W5n/<[Xl�kC��{<W:���u��߽����) �i���\�|:'g�24�(�       �㪬�[�n��j\q/��V鄒�Y�w���2pO���s�h�kC7{���}'T��K�0�[���ѩ�xe6��&J�        �*�if�t�����z{�Ư���6p�`�Ϸ뵡�ͻ�cZ�*�޸��5mt���ќ�p*��8�]�FJ�        ��:�ie�t��u�r�z{�T�ڮ�n��}�ȑ_j�kC7s�}g}4r__7rzþ�{r��l�NH��(�       �����B��!|�:-W܋����~�]/޶�����O�-}8sO�K'��f��wo����`?���ᡜ��ʅK�3�gw�       ��P}8n7o���wޠ_oO�/W�;����m�'��������Ѝ�{�����y���lm�O@���˅�39q�h��\s       �]��,�N�t/�N�ຣ�A�ޞ:�_m��u�~������ׇn����	}kk��[��d{{��` zK���Ա��|�l�W:       �S�ifq������j鄁Qe�tBq������m��>��u�#*,.�����vn^�k����ё����o�����9        ?��eW�{X����.����4=������v�A[�?2�x<��ٓv�t��G����[7���18@��;9���O���T�����       �ie%�l���5��^:���I��[ȷ��m_U-/��f���Eժ�0�X:c l�o�ݛ��jU�S ^Z���ѩ�tu6��+�       �*�ie�t;��F��Ե�����&��v�A���NN}����b��|*��Y[����w\rz���HN�N���g2�gw�       `�T�L3˥3�!u��%�6�Sg�tDWJ����m�gr���u]��}��=�+�0p��6s��]#w��ML���K�szv:##ås       �Pg;�,��`�UY/�З�_ow 9���l�v�ߤ����s�={����n0����#w�_:�/�����ԁ4��9       @���L3��~q���J���}Ǐ�����|g��o���{������=t�g.��%�    IDAT�c�􋑑᜜�ʅK�3�gw�       ���i��9W�wV�����$I�tdޑ�����O'�Js��,#w��LL���K�szv:##ås       �>P��p�n��Ϫl���ΨSg�tD�h��g�x��܏l���֖����{yF�@�9tx_._;��S�h4J�        =�N+����F鄾Pgۧ�k����N�QG�g�66�>x�v'�J�{d����6s�;�?���rrf*o^>�={�K�        =�N3���,B���:U�KGt��|�#��td��$C���N��2�d�t�X7r����X.\����ٵk�t       �#�YJ���tP�Vj�����k�*��E�_��;ul�~�ԉ/u꽠��������WN���L;�F�Q:       �b�,��f�
p��u�������νW��u��ݥ�ťN��������l�o��;w���u��2<<�������88Y:       �B�������|�^���Iu��������}�Soֱ�{�,<���N�tR�����J�>���Vn^�k������̞;�7�<���c�s       �.Qe-���Π�:u�l���Au*��@��r'߯���G}������l!u�i�ne������t�LN�Ngdd�t       PP��4�`+]q�eTٌ��?h(���_�L���V��g��4�d�t�������kg35}(�F�t       �aU6��R��Dm���Z�]o����l��N�aG�7��<x�~'�:e��|�^��;0���r��\�:�'K�        Rg+�,�3�=u>�H΋��U:������~$DG�I�����N�'t�����	� #w`P���f������+�       �Q��4����/�N+u�
?��t�;>p��x��t�=�柸��K�܁A�wr"������錎���       vX�f�YHm��'������9�T�(ѕ��r�߳��k����K�~�w�-�N�%�����}�|�l�ON��(�       �:-�v>SW�?O�V��tF7z��o�A�ߴ��F�Q={���~_h��'�裑�֖�;0���>~8���f����s       ���|�>��0���:�g�= �ꯤ����ܓd��ɟ-��N�O�K'��67�r�����.��1cc�9{�D�x�Tv����       ^R�������|�:[)�S�	u�q�����WJ�o����Ƀ�X׾H�/OK'������Ν��{
,{''r�ʙ������H�       ��T^no��G�I�l���B������g%޸����c�Gs���xoh��{�����ꪏbϡ��r���L�8���F�       �S��΂q;/�6��!�����N�����r��.2pO��T꽡�,�N`�ZU޽q7�+�S :nh����s��l�,�       ��:�,�N�t=����Rg�tD�J�R�˘>s����v���f�V�Jg�CZ�*�n���S`0���f���y�L�NN��       �|4n�ryE�A�����?K럔z�b�������VJ�?������aUU�ݛ����)`pML��7O���S�=>V:       �q;;����:-�����^ʷo�z�b�F�Q�=���R�;i��|�ڠ�����=[*�P�侉\�r&�g�3::R:       L�f������[�~>�WJ�y��{������;e��B�ڤ�����Q����C����9~�H���~	       �q�V�������E=��>�?������/oll��O�s���}4r���3��P#Ǧ�򵳙�>�F�Q:	       �T�f����q� _/�_S�oi%�͒E����w~�d섅g.���w������3 ����pN�<��W������9       �w���w�L������tFWk$_M��]����=Iv��t�������������ݻ2{�x.\:�={�K�       @_hfq�GȴW���ȻN�z�h|�tA���s��^]Uu�x.����r���� ]eϞݹpq&�/�����9       г\n��z��z!�*�Z:����G'O�}t�t������铅|�ރԵ�s ��侉\�|:3g�ett�t       ��V�Se�t`���u���.����\ɷ���(>pO����r�x��K'P���r������Fٟ������#�o9      �����V�Kg0 ���^{p�42��.��������:�����J޻u?Ue��qCC��>������ԁ4��I       ЕZYN� ��S�E�:۩�*��i��#��.<��/��j�������wo�3r�##�993��W�d����s       ��<���N�UpŽ�`���	��ۋ�ƻ�;�.�'����WK7��hn7���V:��V��r���4����4�w����'r���L�(�       ��SR= ��:�I��=�;��']4p?5{�J7��X�[L]��M��������V�t
@W۳gw�_8�g�g�x�       (��%�v�����7��S�������V�P��#]3p�~d���W�7Jw��Z�[*�@���ʍ�og}}�t
@�۳w<.����S�+�       ��RZ1���:I�������w���>X�7��t�G�f���F���g�]�^�³��	t���fn�s'�+��x��&r��̞;�����9       �V�,�2n�K��*��uZ����:��7]�4@�ܓ���Q�^�✁;?�ժr���,-��N�N���ٜ��ή]#�s       `���m�s�^��f�^��_W܏l����Ʀ�%�)�.��)���{����S�F ^T��ȡ��r���̜9��QCw       �C3���t�*�$U�U���U:��<[���,���j�~�lc��݇�(�/����R�u�|�(�͗N�)�F#�����kgs��wշ�       ����.Jӝ���mj��_�?N��,���n)�w�޿Y�^���R�z���Or���� =gh��cӇr���LM��P�t       ��:�,����l�N�1U��ԥ3z�/�����8�77�|. =�w^ԓ�����Ե?<^���pN�<������ԁ4��       t;���U���T}5�������u�;�X{t��7Kw��Z0p�%�=[�{���^���HN�L��9|d��;       ]�q��-ݯN+uz�6u�a��V'�8��z鎏뺁{�L���d�xQKs���ܼ~'�f�C Pʮ]#�9s,��Ɂ���s       ���if������ϫ4S�Y:����t�'�ʁ���Ǿ���e�IOX�[*�@Z[�ȍw�dk�� �c��]�=w��      �.Q}8n�./��ͺ����dmO��\��t����N4��y����"���Ϋ�����wngc���|���c�=w<.�ξ�{J�       0��T�6n�G���*��S���9Ci��G��j�Oҕ�$��3�7K7��������Z�z��V37߹��Ս�) }aϞ�9��ICw       :�N�f�S�Y:^I�*uZ�3^Z�VO��K��/�n�4];p?~�������8]mi��v^_��ʭ�w���a	��b�      @��i}8n�q0|��?}��f鄞T'k{������k6��~���Y���3��λ7�e~n�t
@_1t      ���4����6p���k�%��(�Y-��i�v��$�?Y�>ˢ�;;���|�ރ<~4_:��|o�~q��      ��|ܾ�:U���7p�*�г�4�\��t�����#_jn7��O�ZZX*�@��I��{Z:�/��;�����ɉ�9       ��:�^n7q�Ti&�Kg��*���^Q�����?-��Y�z���6�}���;��,�������w��z��^�g�x�x��       �������=2���W��T������+��������I2>1�S���,�/�N��-�/���;i6[�S ����       ��*[�����'��zZ���n�<]?p�:q�ﵚ-�!@WZ^0p���V7r�������o z��_t7t      ��T�L˸�>����l�����auO�_)�y�~�~uc���P�>���R����vn�};�+�S ���;       ���z�Y4m��u���N���=�N~�Q��Z���t��=I�������,��N�4��ܺq7�+�S �GC�7�<�={�K�       PP+�i�V��P�N�f�OTe3IU:��5R�\����݇�����͏�0�\p�������>ȓ��S ��ɉ\�8�g�o���9       tX++i��Î��+�uZ]��c旳�+�#^DO�Ϟml<���Jw��-�{*�Ϊ�:��<ν;�K� �={�s�x�LޗF�Q:	      �6ke)���΀��!y�:��#�@��ɿ�*]�"zb��$����r��8�)��ㅼw�~��.�0P���rzv:��������       }�N3�ie�tQu����v�Jg��:���/�g���L|ueie�t|�e�)hqa%7��I��n�N�̙c�|�l�N�А�;      @���B*ע`���U�U��ǝp%g�tċꙁ��7����t|dkc3[�=�I���Ս�x�v66�Z(a׮������kg35}��      ��թ�����^%t��A��ԥ#�×�/��5ݞ�'��������%�����۹�Ν����bFGGr��\y�\�O��pO}�      0����|�4K�@W膯�:�]���R�\醗�S˛?~j���O��Kw@�,�/�N��i6[�y�n��<xP���p��Ε�����TFGGJ'      �9�4?���qch����:u�
7�[���x=5pO���s��t$.��}���=���J� ����:�����      t�:[�۫�)�UJ_N����r�4����/���o���_,� ��t�������R�u���74��ѩ���ٜ�����h�$       >Te3�,���|\��������G��ϗnxY=7p���q�ѽGJw�҂�t�gO���{i�<���Fޗ���f�����U:	      `�UYK3����ʌ��T�(���N���o�Q鎗�s�$�X]��K7���t�奵ܺq7��e?*�t��d._�����+�      0pZYM3+�3��������V����g(��[��U������ٿVW��(jy�78t��Ս�x�v��7K� �1N���39�T&�M��       u�YL+��C�'t~�^��V�߳�5[i�\�Wѓ�+G�}�N���􊭭fn�};�� �J��&r�©\�r&��K��(�      Ї��۫8	/��vG߭�F�o |u5�xX:�U���=I��F��������	�ª��{����g�S ���c9=;����fj�P��{�[u      ��R��v�S�/�N����{5S�Ց�u�����gW3���~qkk˯d�YZp�������|�ރTU]:�O�k�HN�<�+o��ə�����N      �YuZif>u��S�'u�k�r�}�-�d�/��xU=;p�p�������(���ZY\)� �d~n9�n����o�����P�Nȕ�����t�v�*�      �S�l��9W��5tb�^e���1x�/%__/]�zv��$G��������	��VW�s���Y[�@�k49tx_._�͹7Nfb���I       ]��懗���)���=p����b���^G�t�����7��9��t��?{�?���R�x-CC��9{<��-��KX]Yϣ�sYZ\-�      �u��������2��jӫ�ie-Iզ�X7���7��}§�/�7�z���ϗ�`0�.��N��VUu��A=�+��Kسw<��8������ԁ��s�       ;��e�v�A�^e3��;�N���'=~�=I�h�>�ժ���>=fcm#��\:v��#�s��T����`�lo7���b�<�O��/~      � ���҇�Y`'��p��׬�J��۠����ƻ�C^Gϯ¯l|���{�Jw0XV�VK'��{�t17��M��*��K���ù�ֹ���ʮ]#��       :�N�f�ۡM�qŽ�Ǝ�&IR�z��ۓ>�'I���+�,+K>�����o����V� ^���P�N��kg3s�Xv���N      h�:�43��\๝���H���c若vB_��8���k�t�c\p��mnn��۷����9@�j49|d.]9�g�o���I       ;��V��Om(m���:�T�ޱ����e�˥#vB_���������}�t�c���>�jUy���<z8W:�״g�xνq2����ѩj�N      xmU6��B�ԥS���i��+U�ء��5~�i~k�t�N苁{��:��K708�u]��������Ե� ����ќ����/��ə���5R:	      �����f�Lۡcv�{���'.��ϔ�)}3p����GϜ�#VWJ'@�<{������ܩ�� (ixx(G���9�����;^:	      ��if)�8P
�T�����i�����I�/��~�t�N雁{�,�/�����%w���zn�};�� ��F#���Ʌ�3y��:�/�F�t      �����B�l����z���n��?���[������s��l��O�ke�������x�v���J� ��&&�rzv:����Ա�&       =�N+ۙO���)0����Ye3I�s)|\���ϖ��I}�\y�X�ѽ��a��ߪ�;�ժr���ܿ��t
 m�k�HN�:��_8��3�2�{W�$      `�U�J3s�y=x]��5X����)��Kk���;���I299�J7���t���ݛ��jy��5r���\�:��Ne��=��      �Te=�,�N]:^�J��T���>����;���G.�����jei�t�����o����V� �hr�Dνq2����#�34�(�      �V��̲i;t�W��^e+�#�m�p9��Z:b�����j������_(�As�����ʍ�ogq�C �n||,3g���[�r�䑌���N      �R�f��z���ԩ��x�N+uO퀿�|�U��w���'�����Ǫ���h�i���w�~��{Z:�α�C����̞;��}��      �>Q����}x��6/~ŽN�����$�i����З��4n���������<~8�wo�K��#�A�h4r��d�_8�7/���#�34�(�      ��:�if�%�@��������vd�W��R�}�tE;���=IZۭ�T����j��hiq5�߾��O�����̜9��_8��3S-�      ��*���b��}���N˧0tH#C?S��]������Ȯ��&�/�B��:����(��'�����t��[:�B������bVR�u�      �K���V�Jg /`8���g�u�����@�O&���}�h�^p���F���~�t�gcmø>G�U�[�s����) 2�o"������LM���p�$      ��Tif��zH�9ܫl�w����q{���$9i��U-Y��ZY\)� =��ù�w�~Z~/Xcc�9q�H��u.�g��{|�t      PX�V�3�*[�S��P��w`u�������V'��W�v�������έ�o��.��N�������o��Ɔ�� ���FޗKW����gr��4��Y      @�U�L3s�{	�F��u[��fGKY#�_]��^/��N}=pO��ё�P����b�/msc+7޾���� @211�ӳӹ���?y$�v��N      :���4��:u��<��������O���ΪR�d�v����ʏ�����y�dv��\���    IDAT�.��V��{�������S ���#96}(���͹7Nfr�D�$      �-�4��VL���}���l�N�P�@z���B�v�����7����|��Ǫ��Z?��{����� �5��ۿ'�/�ʥ��9:u CC��Y      ���J3�^xz]���+_�����ۥ+ڭ��Ir�����l�LvĲ�;��Ņ��x�N67���Y ^��ݻrrf*W�p>'g��{|�t      ���l8nw���G��T�Hb��A�P�~�tD'�����ƃ��n�a�����J��뛹���,/��N���ԁ\�r&.����}��     @���f�?v��u}M��N���;�����{�#:a �I�klן/�@Xu�vL��ʭws���Ե'� �d{�����t�~�|f������      н괲�f��u��T�N+u6K���O�.蔁���?v��=~�T��޷��;���r�ƽlo�8* >���Pٟ������gr��~W�     ��ԩ��BZ�(���G�v�t����J�N��{�Ѩ�=����>ܡ=V��r������^:�011��3Ǿw�}����      PR��43�*ۥS�6���:���N~*�������=I������ֶ�Fx-��>���ܼ~7�ΕN�G|t���W�     ��*�if!u��)@[U��U:bmW�~�tD'���G&��޼�[�;�m+��Vu]����y����Z����s�      :�N3Kif9.�B��?��tuZ�|y-ߺ_���j��$�S�l�z���J��+������Y:��;      �_�V�3�*�S��������GZ:j(�_+��i7p���<�;�߿w�t�ke��:ess;7޾�gOK� У\u     ��We3�̥N�t
���i}￫�;�N������Jwt��ܓd{s�'J7лV�VK'�@��:w>x���?LU���W�;      �VV�̢�+�*U��Fg4��R����\t�Z]���ZX���x�zK]���G�#[(d|b,��Ndll�t
 }�ժ�0���gKY]Y/�      ]�N3K��Y:�:��?6h�d��ꀧ˙�I��Q:�����l4�o?�������u�v(h}m3׿�A�K� �>��~��L.]����������     ��S����������q�sv��S�8nO�{���R}����httt G���'��俸��3�$G��ĩ�i4��2 ڠ��,�����,.�����     ��Ve#�,�����>������P�:�3pZ�i���o�_:���w�ؾ�����ݯ�����N >���Bn^����f� �H���侉̞;�+o��ə����r      Q�V��4n�T���g��i��uܞ��=I&�3��-��IеVW���}�奵�) ���ё�:�KW����grt�@FF�Kg     @��i����� (�:�����{����J������߹{�Ν��5w�6�f+�޼����N��ML����T��u.��gr�D�$      h�*�if.U��S�"����������h%��/JG�4R:������H���7l�y"�Q]�yx�Y�V7r�����[ ���P#N����lm53?��������.�      ��N+�ie�tPL�*���k�������~X���?5���?�y!�.�CW[Z\���~�����) �]�Frl�P._;��N���5Jg     �K�S���vh���i��=�����������û�n�z�ƪ�;t�����x�v>xV:�2�o"g���/��̙cٳw�t      ��:[ifΰ\��$��Ӵ�O>�wVKG�6��$��c������~U2��W�K' /���<��,�޼�f�U:�2<<��G���ř\�r&S�ftt�t      |�VV����/<j�S+u쬺�v3#�tD70pO���;7?�Z�������K�W��}��%�@獏��ĩ����s�pq&�����P�t      $���BZ�#�@*���5�/��w�N	~����?S����>�ƚ��k����u�n�NȉSG��y Jسw<{�����T�W2�l)�Kk�k�     @g��N3���I��i&y�w��u�C#��tC�p��C��ٽ߾����;�n�.�C�z�x!7޹���f� ��P#N��'s孳993�={�Kg     0 ����y�v IR��:��<���|��#�����iT���t�m}��z���F���,-�x- ��ѩ�pq&���f������C�      �yu�4��fV�]>T��v����.�&���?��g�ᝇOJwн6ܡ�5���{�^��y���W6 ���ݻ2}�p��u..������5      ^_��43�*[�S��Q�2n�&7��{�T:��XL|����O�n�{m���N vȓ�����ln�F��g�xf���/����ٷO�F�,      zP+���B�T�S�.��r���E������?�п{��?�[+�AwZ_u�����f�����-�N�24�ȁ��9���\�¹̜9�={�Kg     ����|ZY-�t�f�JG������)�m�?�O6ͻ�����t��UܡߴZU>x�An��0UU���O422��G���ř\�:���366Z:     �.Te3�̥�O�>�J�f�~��|��x�c|��'x�I=���6?�wb�t���������7Kg m2�{Wf����X� x!+�k��[���rZ-�V     0�ZYu��u�l&y�#�C�p&_?��fFέ�w��6.��KG�7��R���Q:h�͍��x�v�<^(� /d��Df�˵9��N���}��<     �AS��f�ہOUg;;1ng'�_2n�d#����̙�����OGFG\��{�W�K' mVUu��y���̜9���@�k4��7��}��:+�kY�~ٽ��?(      �Y������p�T��i���c�������~��O�u���?����;�..���X\X���~��� �[��ٷON�N�ڏ���sǳo��4��     �/uZYN3K���g�R�Y:��OV�o���V.��=�'�۪��54�9 ��\�,� t��V37�����96}�t ����F�́��i6[^u_���Z�4      ^C����.2��N���C0]����\���9��9~�o^?{�������������*��wr"�g��k�g� �}�f+�+�{���J      zL����b�
|�:[myf(��䎿�ਿ����7KWt3��?�pc�ϖn�;l�m�N 
ZY^�;�~��K� �k��#�s��L��u.'g��g�x�,      >C�V��OӸx!M��Х��/�n�v.�������'fOM����|�*�t�'3s�X��='@������r�-esc�t      ���V�R��/�J���M�g���Z�/盗�T�C��H�^����������;��嬭�������W��Fsl�P�M���V�3�l)��ۥ�      T�VV��z��gԩ��v��y]�_�q��rz��w����'s��;(k}���׶���y�n�����  �g��]�>~8���ͅK�3u�`v��4     @��if��g���#;3�?�JU�ZR��V�7��x��1�50,�p!������L2�d�$!7��s37�L&!L62�8�%B��` �-l�n��v�j��Sg{�����I]��Ω��u������uT�z��h�r;�%���D�k�i�#�Cd�Ex��%Gy��p�w �e����3ڵ�Z��u  V��PY6��5�_���ݢ��*��]�        �-����U�:
�LIe)�w�?���酯���*'+��p'hp���P�����cs��  ��N/�_���;        @�Y%�S����<��12�]����
J�p"+(�/��ص�.�9�NФ��쌱:t������� ���̲���]���'5�j�u,        �L2j)ь���<��2\;��wǜ�ς�"Qp_��^x�o�f��{T��]! �_����m�U�4\G ��J���N���Wn�5�_J�        `ѬRՔ�*�n;�%���\?�X�(��!�����8�5����']��&w ��$��<~H��1<p ����>��         �`)֌R�� �(�D�q��}8��N�%}�d��k.��f��Ӄ�����
� �h�DE�z��/Y�����8  8q��vr��$U����lM�jS�r        �*�T�j� Ӓ��;�X�)��Cd�K��K���zt��]�@絚���ta+��t��%> @���+hl|D�^�Q��p�.�2���!y��:        @�X%�5K��22�۳�U}��YÂ�2�۴��à���@�=$"� d��VG��Q��-S����/  ���c�#,�       ��a�T��x5����%�&��X��:DQ�^���8ul�v��::+�(��0�ZS;����ɚ�(  t�g.�_�e�����U�ȡ0        �V��*����"Y�1p�����:G�X����_��h_��::#jQpp���h��ê�յ��u*8k �3�����!���Z�f��J���\]!��       @���&K�@X%�J]��"x��q�!�h�-�_�Cv=��ۮs�s�(v@���ִs�>�kM�Q  �Z��ihՀ6l����nѕ�\���,��        p^VF�*JT���M���2f��+zh�u��b����y[���}�Q�Q�7 �E�����'F�q�|���  p.%�4�~\I��Zihn��Z�)kyR        tV����w���\'�2�/��y�%;v=���="a��
�9Qa� �%��+hl|D�^�Q��t�.�l���GT(�c.        p�(Q��v mgK\W2��woM~�u�,c�����c�}Jy��|�r�0f� �e�}O#�C��V�FK�JC�ٚB��        :�(\Xm7�� ȝH�ڒF�\g�:Z��M�����۵�u���w pjͽQ\G  �<��Ъm�8����DW]�E�7NhhՀ�h         ��RՔ�B��
Hd�����n]�_w"�Xpo���Z�-�cm7�"�tȩ5����h��q�� ��+��U�Ӻ�1EQ��\]����@�r�>        pa�"��Rl�BR�]�O��ΐ4�����s�e�]q��X9���o���w���ǔJ�h˔K��  �+�X�kMU��U���u$        �)V��J���#�HR�w�*��a�1��tMӷ�?iÂ{�$Q��Ƙ�}�u��(�\G ЃZA��;�� @������!��I�Z�H���굦�5��       ��Y�JT�U�:
��_n�u�,�������-�6��};�]qÕW�΁��3��U?�:�ƚ;  ��$�굦jզ����uw         ���S���>DÂ����F,��Q�?o��.+��E�� zܩ5�u�Ǵnj�5w  VH__A��k��aYk����*su��u<        ��Q�TUY�Q �^���v����E3����ޭ�]�k�u������N>�: H��ʺh˔��~�Q  �)I��Zi�Zi�Vm(My       �|c�@'u�����=XӃ���{۰��f�j��Lj����I8�{4-�ھ_�֏k�Ԙ�8  􌾾���G46>"k����*ew��       ��P�j���#��u,�'�z{���>��Gp틮��u��/�*3�1 �y�V�-S*����  ���0V��Te��z�)cx�       �l2J�`�@YYE�9PÂ�3�޾Xp_A+��4I�}�Q�F&��7 ��Q�s�>mشVkW�� @�*��*�F5>1*c�jՆjզjՆ�0v        ,�� \����d��+�����������ƛ\�@����S��t �ixdP�/�R?g�  �&a�.��kM��       ��X���(t@�Id���,�O�nM�/v"�h�����lŏ�����M����W�6�s�>Mm���I�� ��RQ���5�v���
�H�jC�ZS�Z k�y        W�Z��<_�ӲWn��<��u�!�Xp_A����o��/t����W��&��Z5���S���:
  8c�굦*suժEQ�:        =�*]Xm�\GГ���'{�kXp��z��b�}�f��8�c�=�I]G �%i��ھ_�ScZ75&��\  ���=��idtH���굦jզjՆ��8N       @�JUg��#va��kPV�޾�h�����������~�u\�W�}�� U(�-S,��  ��Z� �T�6T�4Ԩ�#       �iV��j{�:
�f�*�}D���5M��u�<c�}������xg���a�����R ���ڽ�֮[���Ys  #<���`I��%��S���Zw���uD        2�*USF��8eg�����\g�;�m�w�<�^����΁��W��  mQ*��-S*��  .P����z ��\        ��*V���R�Q ��$w���w�Ś�Q�)����(�����9P�aV�<�\� ��"��q@��ڰi�
�u$  �L%�4�n���
�H�jC�Z��;        �JUW��u ������'�w]���;�#_x�K7�v�k]����>v�|��\�����拧4<2�:
  h3c��fK�z�z��z-���       ��(T�����(  ��(�����zx��S5M������{�|���&&֎*�΂�}�fI�BɝO#�|Y�fX�.�T_�7  ���F=P��T��P�]G       ��R�d��� ��](����M��S+sC]os�Pp�|��+~��]�����%�SA��|�q ���>��8����Q  @��Q�Ѣ�       ���R5ds�� �"Y��c�U��?\���s�WPp��=����pin�ڱ��,X����;�ŗ�<Ҧ�֩���u  �AI��^k�Vm��h�Px       d�U����� ����.�d�=��_U�{\�LPw�o�������΁7+��� �"���vnۧ��Q  @���zͰ6_�NW]s����Rm�t��'F9�       �RV��u�r;�.���ދ<y���Y�Ow؃�g=R]�i��:���xꗯ��4 ��#��|��6  �V+R��T��Qǉ�H       �f*UMV�u 8#���1���[������� �������o{��h�HF�� �bjզvlݫ�GN�Z�:  p�\������r�z]{å���Ktі)�O��<��_       @gX%�(Q�r;�.e��}���c��k�w����]t���Y�xgZp?�׀<�n ����|�:P`  gE���u�z=P+��"       ���R5d�@�ne���>��C�U�piMߛq�װ���yv�����:�ǨŉP ��l��k�:xL��d  x���>�֦�&u�5���.�]�I�ScZ5 ��=       `y�bŚQ�:�v ]��@�����Pnw�W���};�\~��\���k�}����ė�^P*�q�FF�\G  a�U�l�^T�5ը�       ��Q��R�� �yYE�J]��Yp?<���z��:H/�s��=���/_v��e�./���%w y���<~H#�C�t�:���  ���{Z5��UZ75&k�� R��QT�6���Y        �����b;�L��{���;��K��Z��}�ˏ����.s��w��y���i`�� @��}O�֏kr�qh  ,��Va�.��kMEQ�:       �ì�3_�    IDAT��(r �*��kV,��i�:�>^�t��U�f���$N��W�S�F�|E���:
 t�1V��Pe��M���`�u$  �A��\�W�ܯ�QIR�5���l�T�
[���        ��TM5�l�!��b�!�~���3�]�ß�~�/y������b�O�U���
���5>1��֪P�]G  9��F� T}a�Q���u,       �2
��&+���%f�n�w,'����4�b��'��0�l�����.�K8���
�%\G���9QQ�����q  �H��khՀ�VH���
�X�Fk���h���S       �*Q��BA ���(�\��u�Bu���g��_����׹΁�[��<O��QrУFF���u���L  �45��Fp����;       t�TM5h�$����:�����4�f�!@��k���O��[;|tx�M�.����|��Ӡ<�� �(��495�uSc�<��  ��Xy      ��b*U���� ���*�U�:�S9-��V��u=��uPp�*���������_t�g�܂���
_r zYy������P�u  ���8Q��l.��끌a#       V�U�TuE�� ��͗��1��i��5M��u̣m�E�nm_��ʆ-]g��]X�]��'_mJ �5�v��o�P�໎   i~���l��lj6C�-^`      ���JՔQCL� ȶDF��]!�� �e���y}��i�������a��?t��g��(����( �ԉ�s��յ~���G\�  ��y*/�if�$)M�ZA�f3T�l���
B�A       c�ZJU��q .PJ�=���r{wa��}�k[�^u�5��s��.t��_ey*�����[5<�MM�\�w  ��Ԩ�h����[J��u,       �:V�R�)��	#�H�>��l��x�t���+���i,�w��;����_�y�໎�`Ԓ/Qr I�ZS���׺��\�F���;  н
_�#�<��0����+��F cxr      @o�22j(U�:
 ����ܞkV�ϔۻ-�.u�g��؋^v˵�s�i�Zp���<�S�m' d]�T��͓r  ���a�F=�/�7C��w       9ge(UC�(�ܰ��de\�:9Zp�^���}�� x6ܻ��ǟ�������BYIV�|�K�  ���<~H#�CڸyR�w�   �T*�ˌ�H���
�X�F�t��h�Z^�      �}F�R�d��� mE�=�<y��ޝ(Ow����}_|��_�z�90���x��iH_� �,��irjL�����\# @�c����ZAD�      @fX�JU�Q�:
 ���U���s�ɂ��j�~��83ܻر͟>~�����k�<���-���4(Λ �ӌ�:�Ԍfg�ڸyR#�C�#  ���{Z5��U���ܥ�V+R��$<y
      ��X�jʨ!&; �UB�=�R#���8;�]�O?���x͏���t�+��~���|�/I 8��Am�<�r��u  ����DA3T��Z(���c�      ���j�ʸ� +b~���a�'����kz�߻N���M�嬵����7{�[F\g�u+Yp�$_}�T_� pf��ib��o\+��Z	  z['j���{K�f�V��       ��b���(v VP�un�2^p���MMvg��: ���<��;���_����`e%��W�u �J�Z?6��\]S&46��/  л��>�}<��45j���PA�� �
"Y�M�      ,�U�T�\G��ʰ��#�6���.��iF|�K����7����Vz��_%y�����,��͓*��f  ��1VA0_xo�B�=T�r�`       �b��)���� �FF��o�2����t�S�n��sc�=#�����+o�������(XaF�|�����s�U�ڹm�&֎jjÄ
�u$  ��������*?��q��Dj�"��P�V��ْ1<q      �:��R�e�P�^`e)��O�-�����{��y����ï~�s��N-����L� �X����q   �����Da+Rsa��T      @�E���u ��r;z�.��߫i�6q�!h�fH����:[=8�f��:V��QK��O7 �O':��N�T�q�Z�\G  ���T*U*52:t��ij����V*h��c^�      ��*Q���"�Q ��(��+�]�ܞ,�g̟}�w��ͯ�%�9zQg��y��k@��� Y�y�&֎jjÄ
��   +%M�ZA�f3<]~�-��      @6�j(U�: t�|�=u#�2����5M���X<
�c����{�.���L]��E�}���ŗ+ ,M�ا��j��2  :�Z{z�="��H���[k)�      ��*U ��,C� z�����{=������r���: ���<����i��|��(<��TMJ� �Dq�h���:q|N7Ojp��:  @�y��r�_�r�V�y���ZEQ��{�
[�Ҕ[      �b�R��N =�*��{��r{�Жͨ�>��]/z�-����K�-����'_e�e �36>��'T,r�  ����Q+�����¯      ��U�Tu���e��rl�-��i�Z龖� X^���o�������!��=�*�QK�\G�L:9S��lM�Sc�\7&��[(  @7(|��Ъg����Fa+
�W�[A�0�k-�M      �*Q���B�Q ���r{O�~�r{6��ʰ?���?���W��������)���Tv 2�T*jæ�]��u   ,��v~�=�1�     �yF�J� ] �Q�:D�da�ݓwoU��u,�VI�����C'�_���::�(�'O����r�a��O<�UÃڰi���  d��y(i`����N����P�V�(����     �K�R5eԔω�d(���$��5�!�|,�g����'~�'~���:G/��S|���u ȅ����8�b��   y���t�=c��      ���R�ee\G�.q���� ����V�����u,���/|����8�:G�u[�]�|���: ��{����1�>�   zI'j��(��     ��1����( �E��"�f�B���~R*\Q��f\��1S�[|�-W����J%ּ{�QKy�K .�1VG����Mm������H   �b��w��     �ne+U]F��( �e�µ���{����u���<iN��]_��y�knw�#Ϻq�����$��c @��ԆMk58Xr   ]�Z�(J����{|�m�8f-      +�*Q���B�Q �م�v�:H�u낻'}��Ko��N]g��a�9'v?��M��rÑ��|N{P��|ʣ� mS�5�k�~���h�Ɖ�.z  �7y��R��R�x�??S���{��     �dV���J�� ]�r{��F杔�����?��?}�[��\�ȫn^p�章�� ����&��4�nL���'   \8c�����(���<�     �S�R5eԔu ���N��wﮚ��)�4�r��o?q�W��ΑG�_p�(���*��Z�qB��t�t   �M'�Z�?�6JG���L     ����(��| ��|����N�{5��jj��� h�>��^;���ˮ���B_�u8a�*PA���
 �_�ڷ��f�q󤆆ʮ#   ���>�}g}̙�Fq�(�EQ��_��<     @fY����1 ,�vX���ܞ/4`s�>����u/��u���Ƃ�<O�_� ����G�~ㄊE�  ��<����8�_���୥     �M�.�S��Ű�e����s�i��J�u���|���X9���}����:2�q��o��JePr�vr���\]k׭��1�>�\   t�B�W�Яr���n�U���(Q��O��      :�(R�:%M X���&�'�(��-����?��=o���s�I�ܟVP��; tD�ا����q�  @>�.������8N���DI�*IR��     ��*V���b�Q  c��uт�j�~��h?�W9�w_x����4�:G^d��.y*�W�u ��r��o��5]�    �45�Z~?��g��(V��Q     ��/�7d�� D�ݵ.)���2W���q�A�~}�`�<p����Fyp�u8d�H���C�V�}{kh՜6lZ��!��   ����B�_�r�9��$�_|O�DQ�(I��I���}�P�     ��d���� �Rn�$���m���ł{ν����u?��?�:Gdu��O��Ur z���6n�T�Tt   ȜS+�i�>���ߧJJ��Zב     ��*�QS��Q  ��/x.ص.Xp������N]���a�=����x�/��Ė+.9�tr�*ZXr�� �T�4T�������6��X��   �X�V���8NN/�'Iz��S�     �A� ���r;��BƓ~�r{�������;~���_�#���}!���~���|q� \(|MN�i���>ߗ   ג���S���2|��2o�t�}�3�     ���R5eԤ�	 ��(t��r�ݓ�j��N>8:�fU���￵�%�}�E�sdY^
�����G� �)�4�a\c�#�    �=��3���̿�y�3�K���    �w�����"���]܏������Y���: :��o?���n�����QZt�Q(O�|]G��ǉ�?����a�FF�\G   ������T\�S+�
��+����¼�1�f��녷ijd��k     �m�3��0�=(��٬�_���(;�����ě����S�sdU��O�U�G� �[5<���jp��:
   ��8U~?]�_X�7��s�8oҧ��3~�
��/     �A� V��Uĵ�K�Xp�җ�~]G?(�a�����O��۫_tݏ^q���\gAw0jɗ'�K 8U�5�k�~�^3��'T*q�   ��
�
����G�(��6&    ��Pl��cds}�3�?���Y�+ Ȝ������_��/&1/\�iF���7 �`n��[�����J��u    96��     ��*UC�N(U��% ���Q$+�:����M?�::�s ������+~�U/t�#kn��u���W�%w �"���ɩ1��\#��!   ��j���y�u     2��v Xy��vQn�z��*h�SngM����N}@�ǂ{���o8~���x+�@V�@�HS�ÇNh�ֽ:9S��<I   �}��*;     ������5�b; �(+K��g��v���{�㎷�����9�]�$�@V�} �nE��;�����L�u    9�y�FW�r    �.�t�=Q]��% ����v��8��5�u�!�y�� p�C���C7����sd��c7���!�
�Tp p偒�֏i�����	   @NժM=��I�1     �2V��2j�� 1_ng�=[|UЊwWf$]U���@�>,���o�sߏUOVx$��J� НZA�}{k׎�ך��    ȰU���c�     �yV��uB����#(���<y�F��wQp�a�ߝ���/���t��h�4��� 8�f���w=�'v?�f3t   @y����!�1     p�Pl '�,�v���FU���p��{�������y���W]�@7:��N� �Y��Ԯ�����C
��    �f����,     ]�T�}�b; t��U,K�gJ������(�������ӽo	M�AЕ�K�<� ��W�4�s�~��sXa��    #�GU(�41    �wX���� ��/�[�WqV��iz��p�W.���o|�+����\�@��2jRr�����i��}:t��8q   @��<O�#C�c     ��R��)�	�jRk 'N����~P��3�!�wH��������Gv�s�[Qr�,�����9ml��:tBi��   �ٍ�Rp    ��������� ܠ܎�J|�_��c�A�wH��󝻃���W~%a�gee�  2��cGNjۣ{(�   8+
�    �<�J��J� ���UL���'=4�:�w��7�{�]_��Wv���,��S�A  K��Fǎ������葓2���    <��������     �ũb{��2jQl�.0_n�s�s�]S����A��r���z݁�0�s�� Y�$�:�[�j�DE��t   �y#��\G     ��X�J4w�� �V!]3��52o�����A��r��x�K��»��V 8�Pr��	 dQ%:���vl�G�   �$idt�u     ��(R�YŚ�Q�: �4+���������u���s ��/?|��x���������]G�:�<�ge  ��%��0���,6   ��Z����Q���    ��PF%��  �`���7敯�
n�_u�WtmE�ζ�/C~�J�}�K��c��qt
�dee��2 �q� ��'�Ҏm�57[s   ���ixd�u     ��ʨ�X3JT�� ]�(�v,����8
�8��}�wv��K�9���K����h���9L�   �Q#���	    Э����U�� �kYY�]2,Χjz�3�C�;y���y��������s��>v��]Η�y����(�4�~L�״�R    �\��z�O��    �3�
�.o]� ���U�!�᫨�.�O2k�_��Gڕ	�B�b�����������E0?P�  �Ew   ����48Tv     Y�JUS��jPn��ge�ây��I��Rp ��?������ֿ����|����~�2�*��>q� ȏ$I57[W�RW�اr��u$    +$�5��    �e�(U]�j�J\� ,ʩr�q� _������4��v�A��@�bxw|�[�^�^��u�n����x*h@���|*�4�~L��\Э�    t�z���w=�:    ��X�JՐQ�:
 `I�µ�r{��UTA��T�]�~���9�� �W>���?|��=a��R�r r��ڷ�vlۯ�ٚ�8    �hhՀ|�]    @g�J4�X��� s(�cY�I��A����O��G>����~�9�%V��; �Ew    <���Ѐ�    �\�2j)֌Ud� X2��X�/�4�a�!�L�`)����7�����wą��nv!�<�����  �V(ij��V�Y�-�    t�#�gt��1     �3?���)K! 2��*�Z��|UВ�!�D���8�R��/,�c)�?��{�uYrj�=q ��Xt   �axx�u    @�X�JUW�JT�	 �f(�c��Rn�R0��%ٹ�[G�6O���[o�޹�5V��;]��4�T�|q� �/IR���57WW__A偒�H    ��X��񣳲�\     .�U�T���*v p���b��$y*���� V�J]��
GB��4Œ��w����w�u�N����V�Z,�@9��k�U+�q    ,��yp    �QF��)֬�Z��  ��Ȱ܎婤�Q%L,	w,�����G傃%�2
(�@�i6Z���!�ض_'g�   2`�0w    �RX�kF�*2�\ ���U$Qnǲx�聃�S {
� �v����ra�䭯����\�Yq�Z���;]���D�|y\� ��$I��\]s'k�<���#   �,�<O'g��c     ����QS�*2
�8+ 䍑U,���� _���7��5M��C��3,�c��������ӽ�]�@6�N� zM�:t�?�WǏ��~   ���PY�ρT    ��Y%JUS�Jՠ� �ddɲ܎��*��8��e���a>��O�������e1
�- ��(JNݏ9�4�!   �-<��Ъ�1     ]�(R�9�:�T�5 �-����J����#�яJy    IDAT]�@v\@��=0}|��e����b���Vw��N�1r*�$y�s� ��1F�ZS3��ĉK*8�	   �����u    �sVF�Ud�.�� �+#��ut9O�*��?[��ow2�'��dt�����W����αRLj�������k���� �C|���Ĩ&��T,r 
   p�Zih��\�     8bedȨ)˂/ �#���>��WQ�鏎�]���G;�	��4&��k���+�}�#�X6�HV-q[ �1VǏ�iۣ{u`��a�:   Г�ʮ#     �����D'��A� zF*���>.���v��h��� ȇ;�y�ܷ�y��ny�_�߹	k��zc䞕�d創^ �� u�؜Z�H偒��x�
   t������)Mص    �^`*U}�Ԟ�� � �TV���O�*=��w���9	���_�|���߿���=�:��*�U�: ����ִc�>�y�����8   @�b�    r�ʨ�X'��"C� zPB����]�C ?(���>�_�����n�b��(�v7 ��Vڽ�v�<�Z��:   �{��    ��R��-��w\ ��DF���>c��V��� �
�h��鏟���|�m�:�3\�DVM��; ��@O�~R�wT��p   ȭ���     md*ќb�(U �k� ��(��=����5�u�9�/��?۶~�c×����t��,�b��]��u�de��W�$�u @��D�'k�T�*�T.���   �J__AǏ���w    ��2j)Qu�n��@  ǬbY%�c �<�$I;���)�I�A��XpǊ����ُ>����SE�2jrj pNA3��'��������9��   �<���`�u    �2X�JUS�JT�� �$YE���.�'����� (�cE�#����G�2sl�u䀕�QS�q ���0֡�Ǵ��=:rxFI��   ����    Yb)ќb�(U�� `�](��::�Ó�[U~�u�S�u ��޽�򣉫o{�K��<�u�b��]��u�ge��S�<e�� `�cU�:~lNQ�T�W_}  ��HS��ٺ�    �s�2
��"���" �9��b�?�m�����[�ì�bE���u����3_��W��΁��2j�@ �h�Z���j��ڷ簚��u$    s�\G     ��U�TU�:�DuY� x+�r;�+�
�!MǮ� �(�c�ݗ|��O��ɽ�	
mbN�'��  2�Z��ٚvm߯�;�Zi��   dFwD   ��be�R�Y�:�T-Yב  ]��*�8 �6����/�΁|�U	���ON3�X�ůy���B6�TXku�{�t�`�ʓ'�� `��(��ɚfOV%y(��<ױ   ��V�6E��    �KVFFM��ʨ�Z; �<��bQnG{��u��$j����6F�|�#��۟��gw�΁<�?���* `y�0֡�Ǵ���:rxFi��   ���\G    ��e+QE�N(U�b; `(���<�Y��$�\gA�QpG�|⃟x��o����2j�(t �aq���S3���:xLQ�!c   ���   ����ŚQ�Y^ ,��Q$��h3k��^����{�5-�;�}�}��9�`�fmoKD8���l������ѩ)R�ęX��c���&�f���m�&�!^2DD������_�}��Z�z�g���4��/��~����:u��>���>�}�z��po� ���4?��hg��|���=�Z5u�+c�;�LCϨ "e KF�4�b�t;}�׶rj�*�j%u,I�$i"D`c}'uI�$I�y��@����SG�$M���0u͠�����i�9���u�}���#��������ߔ:˕��>��%I{�����C�եZ�Po�RG�$I���Tʬ��JC�$I�fT$0��MA��o��$]��<uͤpz@�=�m�N��QJ@����n��'�t;u͞ݓ���1$I3���q�3<��	67���AdI�$ͧ,�<�)I�$I{,RP�&g�M������f�]�%��`�\�$�/ܕ�c����o�v��Yb�s�]|�$i/��N?�C�gmu���#I�$Inq��:�$I�$̀ݵ���lP�%�|[�tvGA-�kD��:���Ρ�SN@����/�n-_w���zS�<��,b��uǝ�c�E"#JT�,uI�)�@��acm�� �ިQ�xK-I���0䴚��1$I�$i*E�.M}"E�H�����k��M$���S�_3��gG���g?������|����<��(#�L��*$I{,�H�;`}m�n�O�R�^���%I�$�"[���1$I�$i���)h��m䒤�	�۵����z�S�|�����o��;o�����t��E$�y#'I�W͝�?z��<���!���$I�f��b=uI�$I�
�@A��uFl��$I�)���Di�����r6��:���Jj�{��:]z��o���R�yF.�O�Ȉ����$I�h�4w:ln4)�@�Q�\�<�$I�fG�T���H�$I�D
\k�$�@ ��N�'2����!~�)!۞J��>������r��̲,u��e�}���K��%I�.�@��c}u�~oH�V�V���%I�$��N��0OC�$I�&F$�R�$��㒤}�����~�'���f�$�oNJj"��G~�o������94�}_�&I:01F��Z<��I~��Mb�I�$M�F��:�$I�$M�����S�!:p*I�W���h�]�k�}X�˩�,�kBܝ�և�M����G���"C��1$Is��p��y��8�o2y�#I���T�WSG�$I��d"r��C`�:�$i.�QO���o�_p�S�� ʩH�[����ع�-���Z��e1F����1�gȨ Y�0��9R�v����6��z�F��-�$I��GQ�6[�cH�$I���)hɱ`(I:8#y�������Q��>M�4�(�<��/.V_��W���/N��R�gQ RP��.IJ ��U���m:��J�z��:�$I��ܲ�����)$I�$i�EF�4	�v�$I,�����W������I��J�HO���Co��|��:��AAA��EwI��h5�{�����mBp�E�$I��^�R*9 I�$iVE}Fl��IA��Z�$��E`h�]��υc��H��உs�{:��]�<s�?%� �q��������!gN�����8wv�<��
I�$M�ZݷI�$I�-���9�h��$I�[�HN�ˤ��Ր��.u�ʩHO�̅{N�v��m���\N�mc�;�LC�(2"�D�IRb!D:���t;}*�
�z5u,I�$�I�f�A߲�$I���	z4�K��H�RDr"!u͉H���~<ݧɓ�9,=�����'�_��z�������Xp��%���%Ib0���l���"���B�R)KK�$Is���i�Rǐ$I���R�&�/��ryI�$D�D�K: q�������Y���T�&Y��?�7���}��:��G`@`�:�$I_e�r��:�{�S'.��y��$IR:�F-uI�$I�"�mr��M``}P�4A
��v�������JDz&���gs������_�����>��o���R�Ȑ@�D#uI��JQ6�w�X�aa�����������$I�$��wI�$IS!���H��FF�F��7����)�gSN@z.'O�Xo}��n~�k_]�����1r�w&��J% ��
`iP�4yFy��v���&�QA�Q�\�M�$I��r���cH�$I��
)hS���ԑ$IzZ���(u͝p��@��:��l,�k*<���~be����7��)���y�P%��.I�P!:�k�[t�}*�
�z5u,I�$ͰR)cmu�]��$I�4"�-="E�H�$=���+��,h�7��D� �sq�Q�"���yß��wR�|�"]O�K��Bs��㏞����s��&E��K�$I���JI�$I�E}Fl��AAǢ�$i
D"C��,��L��ID��55����G?��w�|��P:P�@��+�$ISc�r��:���8�N\����$I��S�Yp�$I��F$��E�:#��ԑ$I�L��r�	�1�̯��!]�r� ҕ8�z���÷��֛+�ʁ}�#w�q�}=M�݂{F�?���)#��6�v��iS*�h,�Ȳ,u4I�$M�n�G��OC�$IҜ���(hQ8N&I�J��p�U)��t�=?��԰�����_�d���w��U/<��i�]_�{�r��n9P�4=Fy��v���&�QA�Q�\��N�$I�:���V��:�$I����)hS�!�c)P�4���G����eĝ��{�Sg����M���~�M����ک�h>E���rJ��R��X=�Ƀ�=��c�h�,%I�$������$I�$ͨ��Mr��%I�V#���J'�������HWʂ����n��;~��y�+�����t��:�$IW%���V��9̓�=���FE�X�$I�՚wI�$I{'2��=.�o;8&I�	�܃ZJ*0��3��:�t5ʩHW���}'֞-�z�^���b��uǝ��54�"�� KF���V�v����6�N�,˨7jd��7I�$=�,�X���:�$I��))�)hR�%�㺭$i6D '���R
�����I��a�]S��_�T�]�Λ�|���u,��E"#2Jd�C�4���6[M�QA�Q�\�'I���V*�X��I�{"I�$�
�����.I�-�ȐHHDs,#n�w�?�:�t�l�h��������G����A4�"��xQ@���0�X=�����GO���"�^�$I�%�����$I�fE$0`D��uF4	8$*I�E�`�]�#��a��{S���wM�u>ߺ냿���x�;%��$iִ�]�;��>��3���ԑ$I�4�u�$I��Y$��5.����$U�4��� �6��?�s棩sHת�:��V7�;�y*۹�ͷ��Xh���c�;���?W��  KF��=B���E�ӣTʨ7jd��<I��y�i��v��cH�$I� ��.M
zDL�$̓�o'ф(>7���o�4�,�kf;��/7_u��n�����%+�2�HAF�̒�$iF9�[m6כE�^�Q.��(I��y��h���cH�$IJ,R�QТ�K$Ƿ^K��E$�@�&D8���YO�D��5S���Ǯ?�u?���z��^���u�"0"�X��$�.W�%I���p����NC�$IR�@��6mK풤9���"u	�����_JD�+���������q�kn��~��n��N��	�(� �[I�h5���]��
G�[���fa��:�$I��I����$I�|��D���%Is,���!u	������O�sH{�w͜����3��{孯�ۇ�;�'����x�]���B��鳱���N�,�h4ꮺK�$͘k;�cH�$I�g�!
Z.�J��\ 0�7�hRDFr��7�f�mKͤs��yh�D|�����U�j���<�V��D��%Isg�4w:l��0T��>%I�f�څ��$I�$�HN�;.����RG�$i��S��.��ntS'���wͬ��ϟ���淼���gYp��@1.��`+I�/!D:�U���6Eh4j�J���$I�t�J�����%I��Y�QТ�;.�;*I�����&IF�)h_`�X�,�~�M�Y>������ǚ��HE

���%I�O�ހsgֹ��c{��[-b�!�$IҴɲ�rُ�%I��iv��e�&9�t�o��$IE���5iB$��9��:��_*�H��ɟo~��?��/��?�ݷ�ܧm���.%�|��$i��i�th�t�V+�n�����z�h�$I�L�j����$I�4M"�H���@�:�$I,���Yj�DFw8ug��~�Y����;}����Mo}��K+KW�g�����[���̒�$I@�n����;;mb�z�J��EI��I���f8�#I�$M�@`@A���!Ѳ�$I�"��Z�&�����_+��f�Rs�������S�K_��7|G�|���ܵ_.��/��$=i����V�����J%j�*Y���&I���h5;�{��1$I�$=����G��|>)I�����rh�](��h�}Do3ui�Yp��x����d�?z�+����ւ��W�%w�{�$]�����bs��hTP�W�T�1F�$iRt;}:�~��$I��"�H\jo[j�$�
Er"��P�(v��C}��I�D:Nk�ܝ��+���o������-�N#]*R�Rb�I����|���MV�o��X�����W,�K�$%V���$I��^ 0$�'��$I�:q\n�`�&R������:�tPJ�H��/|�~��G��!� ����RG�$i���ΜZ�{�q��9�;b��N�$)J�$I�}Fl��Έ��vI��Z 2�ܮ��5��/��!$�>h�7>�y�ܹ�ͷ���и��&��]wܹ�ɤ]�/ِ$�Y������[M�QA�^�d%I�t�F����f��$IҜ�)hXē$隅�!1�4����! O�D:H6?4�����O�^���^����s�5�ஃW ��2��#I��+�@��c}u�v�@�^�T�:*I����"����:�$I�4�,�K��F�E.����G��S'�����[�����[^�Џ��Oޘ:��t"9��@)uI��F�ե��R*e,�,r��q��2Yf�]�$i���~f!I�$��%�@���=YI����5�Cc�d��t����H)Xp��;��/�^��/y�㷿�]���HO't�X��K���B��ӡ�ӡ\.q��2�]��C��I�$��$I�^���%I�w�Hn�]�.FF�h��O�"�b�]s�×�����?o��%/��w��
'=5�"�H�u2���H�4��"���ds�I�V������y�h4j��I�$M5�$Iҵ��.I���}K
^u5�ſr��S�RrXs��}���{�����ڷ,Z~��O�����I_-2/�{C���U�N����6��m�"P�W-gI�$]�,�X��I���$I�t��m
Z.�J�t Fr,�k�/8��0.�Isʂ��[�����}�����T����59��
�%wI���hT�nuY��E���^�Q*y��$I�\�k;�Rǐ$I�&V� 2��c�]��"��Ò�dg`����I��,�KcǞ��������v��Ȳ�.4Yp�d��h���Ҭ$I{%�h�tX_ݢ�R*��ի<��P�$I_mcm����.I�$]j���/��	-�K�t��x��k��B��s��A�I�S��ܺ;����_�������O��H�4ҳ�
z���QMG���Bd{���V�J���#�\��C,-/��&I�4�Je�K�$I ����evI���r���
EA�?����A�Ia�]�D��������7����淽�7h�E}2%��H�4�F����6�w��*���?��F-u4I���Q.�1�$I��Wd8.���$I�## �"]���sN$ui���Az�n~������׽�}�=�: b��uǝ��IϤ 
2*@�:�$I3�(�v���m���E�^�Rv�T�$͹��6��0uI�$�DC=
Z��$I� ��r�4-§��o�W I���.=�����=y_�[�������-�K�t@F��v����6�NȨժ�J^�%I��i5;�z��1$I��}�[j/�R�"з�.I�ĉD��5Z��>��ð�:�4i,�K��ԙ/�a�|��}��1�2�
������K�t`����6�[t:}b�Zݲ�$I��Vw|�O�$I�%�������>�0'I��
�r{HD�����'R�&Q%u i�����O��E7������?�_�#]�@��@�z�(�$͕"͝͝�R���"G�[��u+��%I�L+�=h/I���)�	SǑ$I�� ��U4e���r���A�Ie�]zV������������H�+2$�h�a�N���vi������%I�L+�K�#H�$IW-2����8I�4-vW�}Ê�N�ې�OD�dN�Hϡ������>�i���h�`���H/    IDAT��A�$I���A��v���m�!Y�Q�W�2��$i���C�;��1$I����	�(hQ���B�X�$����V��A�+(�͐��S�Ҥ��+]���#��|�*d�J�E�2�HNFF�?��$%c�����b}ղ�$I����a>I�$ir��Rj�Ɂ�:�$I�ba���i�/8���WH�Ŷ�t�������epS�,ҕ�@��-�I�4	.-�o��0�(�v��$I�$���l��!I�$}�HAd@A������%I�f�!^�5��%:��t�S'���w�
9��:/z��HW. #2*Xr�$i���v�ln4Y_ۦ�R*��[v�$IS �Gln4Sǐ$I�����t�CP�$i�E"����4}2�v��]VI�E����)���΀���JF�R�@A��q�]�$M�Ѩ`s���F�Z���#��n�����$I��VV*�� I����%��x�=�$I�������^C�<��ݩ�H��	_�*��/)(}xA�,��ʨQ���I���ewI�4�z�?p"uI�$͉HqI�}HLH�$�@ �r��X��!g~!ui��j���a^�ʂ�g3XL�E�ZJ4�r I�t�Xv?tx����k�$IJg0�y�'Rǐ$I�����Q�8�$�@���vizE��8�xJC�b���i5���7<��`;XS+Q���ƒ$M��t;}�6�l����ɲ�Z�j�]�$�#k�Rǐ$I�L�r]
Z􈮷J�4'"��Cm���N�0��,]��5r�7��ק�"]�HdDFF�eA���B�����b}u�AH��Z�f�]�$�#��%I�t�"�Ȁ�-�q�-��&I�L��{�M�.<�g�0l�N"M+���5p�5n��^�:�t-.~@�[r�'I�4�q�쾽�fmu�N�O�P�W)���K����q��f��$I�B���m"E�X�$)�b\n�p���Z�{���A�iVI@���ʏ�к�)u�ZDr%�R�8�$��i�th�tȲ��^��u�T��((I����$I�t�"�!���w�Y%I�n_ew�Q�v�)����N"M;�<H{d�W�0#|1�oH�E�v%d���$i�dY��R�#׭Xv�$I{�/?J�kI�$�kE
"��:��MVI�t�0.�{�M3!DFp�_�"���Z��/+Q�3`%ui/d�(Q�˅$I���P��u��n�F��:�$I�R���c�"%I��+��%��"u I�4�
9x�M3"2����a�Ҭ��(�C��H�����fE�2@)uI���.��^fq��:�$I�"��s�<�5Ғ$I�ʕvI�t%vW��,I�#~g��_G �r� Ҭp�:7��/uioD"#J���.I�l�
ڭ�;lm6r���Z5u4I�4�6ֶ]p�$I�+�+�-
:���K���Ǉ�g�,�_��Z��I�Yb�]�C��e�-�I�E�+O�f��@���P�n���F���m��!1Fj�Y���$I�W�Xo2�`R�$i��(�P�"�'��{�$��x��/�yk΅��I�Yc�]�'C�~��ߚ�KSg��N㒻�6I��E�^o��V���-:�>!D��
�ox�$I���$�}��$I�l������w]i�$IWiD OB�cq5P���ܱ�I�Y���b��[����ݒ:��W"�d���$i�i�th�t XX�s��2�/��XO�N�$��^$I�fCd4.����J��k��v�i��n���!��K�D�U>u���
�~_ �-ui����QKC�$M�z�ʡ�K>����E7I���㏞��즎!I��+�[:���ԁ$I���s�_h��O��W��H�̶�t s���9�u��H{-�L���H��K�J�+��n��G�)�K�#I��}t�3O��E�$I�-R��CW�%I�>��ۥ����>'6ui��F��
G_��H�E�kd�SG�$I(�2�O��7�F��Y���g��n��!I���	/)���*I��K 0��A�}�6�ď�7��~��.�e��`��|�fRF�5��H��gS�W9tx�C��Y^Y ˼w�$i�?v��V��$I���R{�J�$I: a|�ᝇfU��>����@:N�Jhȹ�ܐoN�E��+d��%I�3(�@��gk������"�z�R�{I����V�~�:�$I�܊Dt)hQ���]O�$I�o���ίfY�������N"���r�sunxp4ui"#J��e�$鹄����l�Y_ݢ��B�R�P.{/!IҴ��n��Yp�$I:8���@o\h��-�K���	�{ʹx2#ˈ���H�:�4�Z��߭p�����"�@A��%��H��)B����jv�U��*�+�>���ʢ��$M�,�:-I���"���>$��*I��+ƫ�1ui�d�͌�{��;�:�4o|� %s��
�OAvK�$�~�(��@�%G�$]�R)ciy���{�QKI�$]����ln4Sǐ$I�)�b\f�-�G�c�$iBDr"��1�}{�����D�$�<�m(%������=uie�h���I��G.���Z���e��%IJ�ԉl�癩!I�4�"a\d�	��ԑ$I��"��W�OѬ�F��D�S��:�4�l H����(� �0ui����QOC�$���%IJ���U�׶Sǐ$I�2�@>.�	��J���V����h�E��I���$ui�Yp�&�a^q4�}XN�E�e�4�R� �$iF]��rh�r��I���wI��˳�ξ�Ҿ[l�$I�t�Ȉ�a<͉������?��RRܥ	��+ޔ�}pnRs �D��J� �$i�]��rh��E�&#I�~8sj��U�$IO)����q�ݎ�$I�&a|0/�"����|?P�N"ͻr� �v9�D������'��'{#e���$I�%Frڭ.�;lm6�����֪�JއH��ڭ.�N?uI���"�Ȁ@��6�q��~�$I�6�G�5?��9�>`�:�$��Dp��7�)u�``T�,�K��P�^w��V���-��E(�KT*��,I��j�ztڽ�1$I��r=m
�O�H�$M�8^m�"�p_���`�J�D�.��Kfȹ?�q��2���Y�����`��.I�t0.�����׶�Xߡ��S�j�B�\JQ����ju-�K��9qi��CA�@\��I�$]�0^m��F�$���[Gl�O�D�WTR������S+<�"��M�E:�� ((� ��%IRy>b{�����0C�^eye��C��Z��.Iҳ�2��$I�jw�'0�؇�K��5�ۥ��7G��s'Rg���|� M��V|
�[R'�V6.�{K�$M�,�h,�X9����"�+�$I�Ĺ�\8��:�$IҞ���%I���b{�:�t��0|w�3�ND���i�4�����|xY�,�A˨Q��:�$I��*�2����K,.z�"I�o�%I�4��B{N��.I��F1.�{���3��H�S�>uIOς�4�y�eJ��1u�e�)� J��H�$=�j����+�9tx�jշ�H����3묞�LC�$�DF��ڇ�%I�\ڽr�]s���>0�ԇR���,�KS����H�9���H/�D�Kb�$iz4�:����"K��J��-I�m�%I�$�D��%I� �ք�A�"?���Ϧ"����]�K��e%J����"��Q��{�$IӥT�XZ^`ye��CK,.�SG�$i�Yp�$I��+��|\h��%I��kD`�Ӝ����>�	��gKP�"�}c� l�hN�(Qw�]�$M�J�<.�/���H�^MI��kv����Rǐ$Is*2"�[h�$IzFa|�T�"%T�f��?�� M�ҔY��{��ʩ�H�d�(Q�˘$I��j���V-���@�QKI��+f�]�$��r�Ņ��B�$Iҳ*��LVk��O�9�`�:���cAV�2C�=T�E2xg�,R:�%*Xr�$I�.�@�?���a}m�����>E(�JT*��.I�|�f�N��:�$I�Q���]
Z����$I��I��[�b��;��K�D���)�4������1�7��"���ȼ�I��b�]�4��;��%I������-�K�$���O��3z��I�Dҕ�4����l����Y��vd��K��e�]�4ZM�$�jE"�K
�M
��QY�$IWnD �7�H�DF��gϧN"�����[���_~$u)���q�]�$i~T���X9�����F-u$I�:}r�����1$I�T��q�=/�J�$����UHD��C�?�:���cP�n�E�Ǘi� ��MFJ+�Q�D�pI��y��#��Zlo� �$I��I�Rh�-�K�$���vi,#ne��s�r�4�l�I3�����u��H� �LF��r�(�$I�Yx�$�%I�E�0^�-�F�#I�$Ͱ8��*R�&E���s�3��H�6ܥq=�s(g�i�h�,Ҥ�]s���!I�4Q��
�u��X^^`q�A���$�ڜ:q�����1$IR��C�U�$I&�W�C� ҄���������I$];�`K3d���>|G�,Ҥ�(S��RG�$I�H�r�ť�%��J%?.�$]�$͏�,����m�J�$��އ���C(~����HD�����4cxً*T����Y�ɑQ�FF-uI����e�F������Ej�J�X��	w��y67��cH��=������1u(I��9<d(}�"2���SJD�ޱ�.͠��� |}�,�$ɨ�Q's�]�$�T�������XOI�4a�;��V+uI�t�"�xI�=�
*I�4AF��3J����9���"ioYp�f�2��Ό��y��H�%�D�WH%I��V�\bq�𾴴[z/���A�����eg��:�$I�B_)��.�J�$M,Wۥg���>'&uI{ϧ��;�+_��VRg�&MF��J�$]�,�h,�X/�/�,R��Sǒ$��=M��MC�$=�xI���/�?%I�&����3��q�ǿ �L��'͸e��1��h��"M��x���$I�^k,ԟ,�/-/P��I�e�=r�v˂�$I�$�/Yi��$I�����qE� ҄*>����_m �*��X���c@5uie�(Q�ˢ$I���V+,,�Y\j���`q��ʻ$͐G:I��OC���������n�C�$i:r���^F����� �f�M>iN��G�(PJ�E�D�x���%I�L�^eiy������{��Q�$M��<A�;HC��9�E����֟$I������e��>O�S���|?�4'���oWx�2d��-�׈
���K�$�� g0�a�	@��=Yv_Xl���H��G�4B�R'I�~������vKO�$I�%���|��L2�\��]Xn���=i���"�_�sH��5wI���Q�VX��/--���@����4i���CK�$iD"#�K�=L&I�4���0�(ui���g�M��LD�����4��ʟ��_J�C�t�k���1$I�t�,˨7j,.�YZ�-�7�Ա$i�=p�1�C�J�t5.�v�ه��K�$͍�Ì�eȈՃ7����Y$�i�94��npC	x}�,�d+ƿJd�R��$I��hT��h�tX_�fmu��N�� '�H�R�T��M�҅���XI��K$�RТ�G`0^��z*I�4��%=��`��[���H�D����.ͩ�>S�:pk�,�d�Dr222/��$I)�H>�i���l�za����nwM8F*�
Y��$i�\8�I��$Iz���Ҁ�m
:�2{�R�$I�\
r�^P����\HD���ɮ4�V8z�өsH� �L���.I�4u�,�ި��Xga���勒�H�^��|Ԃ�$i���O�%I�$�ڽ?��!M���������Y$��S\I�!���?�:�42 �NF/��$I��һ$흿����$I:`�o���nY)�%I���tq���E��������I$��[I �
G�oS���k�$I��һ$]�"�|���1$I�W����'W7]g�$I��p�]�R�l�79�P�$�Ҫ� i"�7��2ǖ2x�0�4�tɨS��:�$I��H��~o@�7��&��F���R�r�Î�PE��$�HA�?.$�D��$I�"��KW�| �u�I��\p�t�����@�}��H��5wI���T�VXX����`q����wIsi0�y�'Rǐ$iOE#6,�K�$銹�.]�������ėSg�4,�Kz�o��p�?@�-ui�d@F��Z�(�$IJ$�2j�*KKu�4�T*���$i_u�y�D��$���1$I�45\m��F������H�E���.�i|K}��ޑ:�4m2�d4�\s�$I�X�\z�𾰸[~_X��e~,#i6t�=}�T��$�H�т�$I��U$2r�]�
q�;z��|�,�&�OR%=����~$�9uie�(QOC�$I*�2���u�u���K�J͝�;�:�$I�"�gD3uI�$M���Wۥ+�w"Ż�����Y$M�]l��oJ�E�F��K�$�JU�5�����U��%M��Ǐ�KC��}3b�@�:�$I�&����5jB|w��ID�d�騤ge�]�v�k�5��J�$�j\�������뮽K��;�:q!uI��M$'g+uI�$M�@dH$�"M�&���9�'��H�\6�$=�q���7��"M��%�%$I�$�j���b��B�F����n�]����6gN���!IҾ�C`�:�$I��r�]�M���ħS�4�,�K�,��ސ:�4�\s�$I�~*�K��U���'�׫��I�a�or��z��$�H��7:%I��V1.���A�iք�}N�q� �&��:I��|�R�������H�,�DF��5wI�$�����3묞�LC��}WЦ��:�$I�T$�)R��]�D��.'>�:�����{����;������-yfd0X�&�1�\l�lb��l �d�B(6�M*����fkd�IQ�J�F0���������`a�\����H�-�-Y��Fӗs���A��F�$ϥ���zU�$�U�̓�>��s���`�\�����g����-�����o��  `���Oܗ��;�: �@�$��	 �6f�3I<����.�wl��m,w�=;/=1��CI�t�Xv���7S2l�  �2|�����T|��� p$��d��3  8T5}Ɖ6�A0n���;pM���7M�%yi�X%�tيo�  ,��������]��Q66|`��]g���9C? ����Y�  �4}�q���.�;�s��C��cE\�g�Ϝe�$/i�����(%��!  pU.�777��5���(�͍lm�R�?��;u�'�ȅ�� pd��e��Zg  p������v80��o���l,'�0�e��{�`R��u���k�I��)  p�66�ٺa��h#�͍�p�f6�F���h���������k� Gj�s�  ˮf2B���p@.v)߱�3?�:X^��u��|�3���3I^ٺV�k�  ��RJF�����������>�	�䣿w&��u ��I&9�: �������z8�}�n>��C��f���s����$yU�X-]�J2h  Gf0�>���hs���Q�Ώ�`���o��l�` ��4��g�: ��VS3M���A*�C5�����_j�,?��朼���ה״n�US2J�Q|� `��R2��x��������(��y��j���߼�u 4Q3�$��  ���W�k�X)%��������˭[��`%����X��/�k[���)�R���;  |�RJF�aF��6»��k:������ ��,g���  |Nu>l����SR��̾e7��ϭ[���=�����9q[R��u	����tٌo�  p��n>z=6~�l\���q����j� �����3� ,��d�>�����>�L޸�{�k�`�X�����ٺ-ɷ�.��T�e��Q�  Xz]W����;\��ws�~�u 45�#�e�u  ��O�I��u���t�~�v>��C����9��`t<[�>ɷ�.�UU2H�VJ��)  ��66�ٺa�Y���͍^���~�bΜ��u 4�g���&    IDATR] X55��L[��*�������V��;p�^1<�?Q��n]��d�.���  Gk8dc4�����x�_7���P�{�B��l� hn����H�  2K�i\m��T�d�s�o�.V�p^1<�?Y��h]��K�͔�  ��(�d4f��?v�t~cc�׶�F�:?�cy������Zg ���+�T  m��LR3k+���;����h�`�y�8"oϝ?���k]��d#]6��<  ,����h>z�|?�ecc�
<�Sgȧ�}�u ,�>;��B� �5S�����:VZI�d��������-��|�R9����$�u���.���Z�   ש�J6F���h#�aF���]�w�V���}����3 `A�L򠫡  G�O�I�):p�$���]w�.փ�O�Q���#�xNN����1��j��%�e��$]�   ��}���8{���w��dc���c����h4L)����Ԁ S2ȍ�� ���ij��C`M�S%ݫvr��K���-���9�������.JF)��  ��`�ec�����|?�lW����#�[g �B��W� �,}�q��J�oÔW?����.֋w��&.�#��xn�I�ǭ[`ԌS3M���� `m�f}f;{��y�����p��|������l���:xR.��������  +��_m��8:�7vӿ6��|�`�8�
4u,'�jI�E��)��f��  ��`�e�1�p8�?�_�σ��ï����3�L< �h�S�{$ ���ί���!�N~m7��3�֓�;�܉��k�[�p�JJ6�e/  ��v�*�`8�`�ͯ�?6��4�n3S�?�,����;R�7�����e; ��ӧf���u����K;�1�w�u���I���o��c�uZRߖd�u����q��R���A�   `��Z3�L�����1���������~8��V�әq; <�.��2�_ �����}�:��/�$ߜܻ�:XoN!�xnycRޝd�u���k���   XF]W2<v!~0����_������:\��N;;{��G�n� ��8Ӝo� �Dj���C�>TG�$��ɝoJ2i��`���-��)�IrC�X?%]F)و�  �:x�0��k���0�sx��vN���� �Ц9��6 �
���M}�XW?��;�7~�;1��9�[_QR:���-��d+I�:  `�R7x���`>���.�����n���~}�?w!w�9�: Z�$��k� ��jj�����5V��n��P<:X ��B�)���S>��Z���*��(^.   �K�㻮�t��/]�/]�؅�'�������|���}�����p� ���$���Ʀ��%�?����:��,ր�u,������I�H�X_%]F)و�   ��c�R�n>����R���7�_���G�<n@�㩜���|��G��) ,'W� ��O�$5}�Xg}����;�a��'c�,�g�El���I�[`�ud+ɠu   Gl0�RJy�|)�`0�xo������JLs>}ƭ3  ���������2铿��3��u�S1p�3��/�2�P��n��d#]6�%    ��s� Xo5I�>����&�������! O�:X
���9K���|m����(%��!     K�w `=]���C��b�|�v����! �K�: �J��o��1����C�[��>{�e;5��1     Ka�g�N  8B55��ًq;�W�sI}�q;�,� ���|z2γo���O%���=��$���.    ��J��x +o�j;,����^����u��2p����q^��͜{^�[Z� Iҧf���7h     x*���m pHf��x8,��򉚼j7w�^���a�,���q���fn>��k[� �jf�����_t    �r�� ���ۧIj��1w�^��3w��Z�����Ϗrs-�+[� �����������A     �K���  d�~�1�H�GF�|������% ���Xj����<��IyC�d4,���O���    �J���s� Xr����f�:x���ws�{��C�[ ���;���9�ۛ������$��=��fI&I��A    �s� XV}j&�<IM}�n���d{�u���4V|�}5����!,���>;����     I�l��� ,���I������v�~|/w���_"Xj���x$���5�eI�m�|��Y�lϯ�$?    ����u ��If�a�������9���X�u �A�)/��}fJ�[��R�e��Q�    �f&y�T `���3Iҷ�BI��)k/��E���d���g�_X2�`I^Ժxj%]�l&�    ��>;��B� �'�S3�A<X|K�};��ݭC ��;��� /8����*��Z� O�d�.[��    X/5�<h< ,�i�L���!��(�����ws�[� �A� �ò����<�������{���'�&)��    X%%%}ƭC ��7K����(ɧK����̇[� w`��?���޻�s�Irk��s��f��KCw    ��V2L�ݸ�
 �ѧf��i����S5�W���o]p�,ǀ5�Ѻ�����]��o]|n�Wfٿ^Ե�    8D%%q� 8b55��L�v�J���^���>ٺ��kc/gy3��xRސX����+�$��;    �������  �¥�aǩ��4J�+;���|�|���PZ ��r�u}��o�\��Q����    ��f��Y.��  VVM�ϯ���r�n����I2m]pT�B��C��ϗt�Nr_���Ռ3��Ԍ�y    ���> �Cѧf���vX6}I�G�9��1n֌�� k림�K��L�'[� W�K�͔[�     �Y.d��� ���S3Mͬup�JʤO�;{9��Z� �`����y��%ӟN�׶n�^� %�)�N    �n5�L�@� `��ˆ�.���XR�w'g��:�k0`��s�γ��d�Uq��PM�$I���}v    X^%�+� �u�If�3Iҷ���}%�wr�Ϸh��X{���8/�m+瞓���=���/�[�     \��a���  ������`y���>��˙�j�К�;@��u/g?���w��:�@Ò�%�&���;    �rٿ�>Nuu �"����4�܁eT���������u�"����8g?����J��	K�ίL�t)�Z    \�A�춎  ��S�/=�Xj���u���P��E�B1��xF^��.�O%9Ѻ�>%��l�    Ke��X .WS3��2l�eWҽk'��;�'��Yz<����_�S�.�'[� קf�>�g'�<    ,�Anh�  ,��d�>{���Ò��_;9�]1f �,.�<�������?�䅭[��PR��.�x    ,��IH�u 2K�I��ae�R~�bμ�u��� Xd�|�<�'��0ɗ���,5��$%]�   ��T���LZ�  ����/���$&ݟ�ə��nXd� ��v����۶2~N�[[� �f�d����^    ���0}�[g  G�O�d�A7W�aU���Y���˩_o��謹 ��]�^�~`+7�O�8�+��f��YJ��Ew    �EQ��TJW[`=\z�ҰVMI�� ���ɩ�[� ,w������6��>Z�oN�Ѻ8(��;K2H�    `A��g�u p�.��I��1�+)�q'�7�s���- ��z�ϋ�&�ޟ�Z� �d�.����    ���\�LZg  �&���4.��J�]����������5�����.��$k���if�N����     �����	 ��ۿؾ�!6�WX5%eRR��vN�O�હ�pN�k�]3yoR_޺8,%%��     mL�@jf�3 ��֧f�����r�K���~_��e5h ����ɝqn|�([_R��l��Yj&)I��O    @%I�q� �����fǜau��Ou��s�?�nXfZ ����8g߻��m$���5�ᩙ�f��.%]�    `���g�u p�.]l�İV[I���͗o��[� ,;w�2ν�i��}�$oL2l����ijf))��    �ٿ�� X|��}E�vX%�;�$gεnX�u ��9�}Mҽ/�sZ� ��d��Q�ϵ     ��f�Il� <��f��Z�]������� ���ܔI��g�|y��h�ݷ\t    �4��g�: �,u�����+������9���! �����|~����3�Z� G�d�.���;    p��f��[g  ��If�3��Ͱ>J�`��s�Z� ��A� �U��O��yٻF9�����upT��G�'u)>O    ��A��ƀ Z���LR3k����3z�NN�z��Ue�p�>Z�9���<�lR�1N:���AXS2��     ���6 ��U���36l�5T��w+����=�[ V����)'_�'�%��up�JJ6�e/�    ��U3�$�� �54K�i��u�@I������ħ[ �K� G�|��k�˒�պ8j55��rq��B    �kW2H��� �Ff��K�q��a���II��vr��b�p$�8b���K��$��[�V�t�H2�b    �&}ƙ�|� Xq����Q;��r�d��vr�{[� ��A� �u3�=;�����l��$/l��PS3K2I��t�C    �j��g'��H 8����^�$w����|�WZ� �w�&��s��[��|��&�Zm��R3M��R     W�·w ��0l��t�u��+���j����
h�Dny}Myg�g�nZ+�2Jɨu    �jf��� ���L�Oa�\풷o���O|Q h��`���o�\��%I��u�ZM����N�4�B     O�d��� �}j��g��$�����Ν)�� M��� n�W>�f㶚��-�b(�R���a�    `A���4�� �%�b;�x%y���/\̩�o�@2h ���ܷ����c3�6���u��?X+))�    <A� }vZg ���4l��Ӕ��t�_��;~�u	 ���G�8ga37ߓ���uHri��4Cw    �r%��z �S�S3����1�B)�����Ns��[� ��: �'w</�ڤO�/l�,��AJF)�N    @�4�<�: P����O�/���NN��x���1pX`7�d�����l�,Cw    ��iΥϤu ,�v�i�R~�bμ�u On�: ��6�=?+_�t�Oʗ��M��Pn����k    4�g�: �S3M�$I�:X@%��Ky�v�|�u O��`�]̧'�}�fn�I�x��Y�   `ݕ�g�u 4b�|n%���R_��;oo���3�X"'r�7��w$yf�`q�R2Jɰu
    p��y(}�Zg ���a��u��j��};w����e`��dN�?QSޗ��[��f�    ��^�y�u �v������^N���! \9w�%�y�����I�s�[��g�    �f�Ϥ���C�χ��!�(ɧ������[� pu� �z۹<ν����;I^X�V�_��%))�Z    ��$��f�
�S3I�$�A.�
����R�~;w�A� ���;��쇷��H�$[�{�Ewi�>M��   �
*)��: �a;p�j��}'���I����1 \V����Kk�K��[�eҥ�FJF�C    �4�gRӷ� ��Чf��Y�`��d�t��NN���- \�V�^>���|��g�~Y�?պX5u����O=|�    VB?�t ���v�ڔ���m;��Ѻ��g��"���8go���;I^O� �X�_��􆗡;    ,��.}vZg �U0l�]I��d������- w�3��o湿��oJ�ٺX.�.�'5%���    ,����nX|���<���U�]o����i>�P� ����:����d�SI��u��JJ6�e/   `��r1�\l� O�&��g��o,�ݚ������h��s�`E�s�7��o�e�'���u��f�����    Ke���N� x�i�L]l�KI��d��ݜ~O� ��;�
���㽜��y�٤�>��ר·�IMICw    Xl����^M2K�Ijf�	�%�Ãt��Ω�[� px,� �����uI�-��n�_�FJF�;    ��fy$�l�� `��_k�F����to���Nҷ��p������fp[R��u�J��2�D    �⩙d�s�3 X;�������<<�����j]�ѰDX#�|��8��fƛI^ֺX}j&IfI���    �@J��B �F��i�I�����)wӽ����˭K 8:.���9��5ys�g�nVI�.�)�    ��r!��� `����/�����;���'��X3� k�y�Ww�~*�ߺX5]�l�d�:    �Z�$��k��J2lGI&5��s7��a� �0pXs��KOL2}k�ok���.]F��^z   @�|&5}� VF����-��()��2�����[� �Πu  m�䞽qξ{��g%yy��u�J��r�$IM2H1t   �#��3�i� ��,}&��)�u��Jʯ�l�b;���- �e]�����W��w&���-��*)��(>O    G��n�y�u K�f�>K\lOߥ{�vN��If�c h����9��zN��;j�[� ��d��Q��
   ����3�gZg �T���R3�k���*3��Gr��Z� �8�� x�q>}q/�[��$/�C��O�$��/).�   ��()�E >�>5�$�TہCV��^2|�vn�/�[ X,F� <��囓�I�պX}%��E�a�    X9�\�,;�3 XX������ ���t��I��S{�c X<� <�g���&�%yi�`=��$�2���    p0��e��Zg �pf�a�k���������~s� נu  �m7g�oe�D1r��,5���$���    �V%���n��B���^L�t�� G��f�5s�[� ������9�s[y|C�Q�"`=��W�>Ig�    ׬�f�B/�Z�4l��f�v�(�t����kǹ��- ,>! �����$�N��[��S2H�(%��)    �tf��Y.�� ����BF�@�5ÿ��;�Y� ��� \�q�~�<���xI��u�n����t�ÍOl   �*I��� �����\��\��UR���M��㽭[ X.�@ \���{��-ɍ�[�uեd�.�xi    �K�$�����j����T�v����nH��s9�P� �� ��X^��%ݻ�|E�`���S2JI�:    �4�ϴu �b�>���4�[��c'w�H� �נu  �m�O�?��u3�/LrK�`���=b�3t   �'����`u\��>I�,�������7��̻Z� ���8 ���s�g��;��.ɨu����q�)))^�   �ej�쵎 �]z?����ֺ��1ݫ.����% ,��: ��r<'�,�mI��u@���$�2���    ���Y&y�u �l6��n�,�������;�Y� V�s� �q�~f��e�񉒼�u���eL���    �OI�>;Ij� �X��{����k8�8��.�o�ɩ��.`�X� phN䖿XS~4ɱ�- �+�d��a�    8rӜO�q� >�>53�v`Au?���7%��H� V��; ��xn}~Rߕ�[� |�.]6R�/�   X�\�,[g �j����|��pv���vN���! ��A�  V�8�>0���:��DI^ں������$IMICw    V]I�g�u �S�����i\lSw� �����u	 ��z�#s,�|gI��$7�nx*%Ô�R|   ��U3���# H��k�F��ª%�w�d��]>)	��3p�H=+'��4yG�?Ӻ���e#Ɇ�    ��I��)hc6ʬ����+R��Ŝ~[���(    IDAT� և�� �ݜ}h��m+����t�� �ܥ�)�$5%]|>   �UQ31�hb6�<�����+�~+�z'�~�u ��B�f���+K��$�k�p%J)�d�:    ��,3��� k���Z�Q;��J2+�y;��Z�S� =w �:�������on�p�t�H�F��   `���4�� Xq��i�����()���o;��l� ֗5 �Dn��>�GKrc��+WR�C���u    \��Y&y�u����/���C �JI�K�����Z� ���X������L�[ �V� %��[�    ������� +����g������I������u $ɠu  \2ν����oev�$/m�pu��1�Ӕd~���I   X\5cׅ��l���$�5XJ��^��S��.�K,n XH�r˟+)?��٭[ �U����{�:    >�,2�N��%T���g�v`�Ւ�];�}_r�n� ���; �y����dR��u����0��p    F��Ls�u��S���YI�w�������- �d� ���S��y�Ol��v����[�Ҫ�xO���EwSw    ���X'��6M�d>lw�Xn%ݯ׌^����K� x*V5 ,���%5��%���- �d��QJ��S    X[5���:`A]��>KR[� \��LJ?��S�{|a`����R�˽��ȗ�u���%9ٺ������i���    4Q��� ����]kVKI�;�e'��ں �� K�Xn����cI>�u��)�]u�9T    ��4��g�:��K����+��t�����'��i W��������Է$���[ ���}#]��   ��4˅�b����|�>kp�Jʹ.���?|g� �ZNC��&���q�}�Vn>��I��� NM2M�8��b��t��    XM�����If�3I�t�� ��d�+%�Wm��u \� Xz�r�W�ԟL�U�[ K� %Ôl��x    J�q�9�:���$55S�ځW��~d;w���% p=\p`�s�}�<����O��%��VR���}�������   ���:�������A����l] �� ��rSN��Oޚ乭[ � ���    \�I�3�V�k��z)I_2x�v6�j����= p�` X9��U�)�xR��u�Q)�d#�Uw    ��$�/,�K��gI��1 G���-��vn���- p��XY�r�M%ys�g�n8:�t�H�0^�   p%�y(}�Zg \���O�̵v`u?������]�[� �A�x`�=3/�c�toM��) Gn���FJ�S    X`�<�Y�[g \�>I�Z;��Jr�K�7/��[[� �a�t`���S�s�m[��\�W&�n8:}j&����%]|�   ��6K�q��+��s����ٿ��>J�_*�x�v��ϭ[ �0Y� �6���/H�����- m��R2r�   �GՌ3��� O�O�,5��kl;���ݜ��C �(X� �6ƹ��qn~�VJ���t�� �ޥ���TW�   H���i� �����i��u@3%�GjF����m� GŒ��t"����$_ں��Ǯ�[�    ��8��N �k� �)�$���_��Z� �Qr�����������o���%yI|�Xku~g��{ҥ��   �V�/��-�$����\���e�vr�[�E k�j��w"�|CM��Inn��8�2L�F��   `�Ms.}&�3��Q�|ŵv�˕dV2x�v�?�ܵۺ Z�T�$�s��K�j��- �d�Ô�R< 
   `eM�p��P��ҵ�Y\jx��r� �����Ժ Z3p����7��_%���- ��K�0]6�t�c    8@�\�,[g +k��i�Q;�g)IM��~' �w�u ,w x�c��甌~4��u��*\v��+    �]��Ls�u�R�����'WR>U����z� X$�( ����4��nX\%%)���    ,�>�Ls�u��j����\kxz�d���̾�\�<�: ��; <�g��_ԥ��I��u��+��c����   �r��e�Zg K��k��1 ��ܗ��N�xO� XTV' p���,ɳZ� ,��������   ��jƹ�u�T�$���e���PK�����/��]� O�� �Ѝ9��A��$ol��<���    ,�I>���u��j��zp����w?��S��u , �B��}d���~3Ͻ7)�H�ٺ	`9����f�������   ,�>�1X��,5���z���p�J��8H^��ӿ޺ ��U	 \�g�_<���$yU��eT2x���?�    ,�iΧϸu�j���Yjf1h�z%�|��ߺ�;�Һ ��� pv����w[���$/O2j��\.�12��U�2��   @+5��S�����/�O�_<��Z�t���bN}�u ,#��:=3/��>ݏה״nXf�������    Go�G2�v����d~���\���`��ߺ���u ,3w 8�Dn�j�?M��1 ˯K���ލ�   �B��Ls�up$.�����Z� ��Z���0����?�: ���; �s��G�|k��UQ2H�_v�G   ���g/�<�:845I�_j���X%��I��vr�ݭ[ `UX� �!8��o*�C��k��J.�K��   ��U3�$�Zg �ҕ�Yjj��URK���������c `�X� �!yF^��]&�2)�޺`��'��  ��g�>c�<41�_Uw��(Rb��3�$��"��QI��]-��1g�������^'�����q^�g����8�޽�5ʉI�2��HCI�,QL]�T7���$R$��~�T�lꅠnV����W�LO�僪c �D#I#�����Z*R�,���O�?�: �"w ��z���,ɴ�� ��"E��޲{��8    #X��y���wV���~>�R;�uQ$=I�_�M�G��'U��V�� C`r�Lid�?N�?�:@k����$m��    ����V1F��R{O��T��)ި��?�"����, ���`M̆���M2��, ��H=E�R�-Qv   �,��,�}K�_��"�)R�W�r���_Yu �`�Mʶ�e���I����`H�����G/   ��;���ȹ�c _Q&),��U%�#I�wO��cU'��D� *2!�w���$K��0��݋��%   �`��I9Su��Fo��'�R;��)��I��2s���W�� �M��  0Z���7�f��>&=mI�%�U�	`t�;u�$=I�~   $IʜK.�V�{��{�UU�����y��L^�C *`� ���ٴ���_$�ƪ� �NE�{�   0Z���䋪c�(�H�H#=Qh��I��α�8m Tɂ; ���ɳY������L�Qu&�ѧѻ�t.e��Uw�	   F��i�l�!`�h$�I���	eѧ�F�ړejw�ɱ��: �� ���t/*S��2�Ug�6`���  �����ϧUǀV&�I���B; U*R|T��_�ʑ^u ���; OŤl�q��H2��0 $��   �h��ٜ��Uǀ��0�I�o�������V L� ����4���?M�P�Y H�   hMe��\>�:��2I����Su (R�&���_���[u ���`����W���In�: +R�]�   h	e9��VF(�v��Hz���婜����_V� �z� 0��;/�Ϭ��'W$�Ԫ��@=)s.e�%)S���   �HT$�ɩ�c��Wj?��aO�c /���~�e������U� ��w a&gCw#�?O�]u �^�Z��'�[v   F�syO=�Q�[doXj�����<�#�m�6 �Z 0�o~s6���؜�0ɭI:�������">�2��\m*RXv   ��F��j�X�����ɱ�' �[�ړe��{:��?�C F� 0�MΦ������T���UK���K-^�   �͹|`��4K��!�F�a �LE�n-�Ͼȉ���, �w�I -`b6<��,�쪳 p%�e����    $I��4r��P���v�v���Hz�ڿ����q^���< �wW�:  p���7��ˌ�Hm\�l��� ��Nkܬ��Q   T��3�e�ޣk�O�,��U��
L�<���3��=�c��t>>]u ��Ԫ  \��ǟgߟ$Ů$/V��+U�̹4�ez�E9�{@   `���=�A#ɹ4r��C��� #N{{{n�sS����Ǐ}�cW� �6ڪ  \[�e�I��I�T&�(���3p��ޥ�s)��iK����f   �z+�Ѳ�g'�IiZ`Ļe����sgn�iRʲ� Z��; ��}�>M��I��WI�Y�bOՉ �n��ƞ�]�J��S�-I���   �u������i�L#�ZÄ����vf��UG �w ha�f��$ߛ�)��L�V�	��S��we�Lo��o�]�   �V���HV�o��Yj7��*�ZV�]����]�9��8 �u�� ��g���3�������$��� �%4НM��Ij)��{�W   �
�8e���{��up�iy��2g����  C@� F�ws�$������k)����^u& ��FJew   ��Ppg$��ި: �Ig�캣;;vw�Vs� -�`��"�Or�l�q��$�Vu& ���e�"E�)��[vw�   �6�?`��[ho��hUEQd�ʅy��wg��Ϊ�  CL� F�����W���/{����?�# -�L��)s>Iz���u���	   p)�.f�(�Wfo�˪0n�iJ~�wwe��9UG *�� ��'9�Q�?�w��>��������>�: �Y��=IΤH-�-�7��   �烃�4�_joD�`���h����r�]S����L� ��-�_�ڴ(�=�Z���9}��H ��³)s6�C���d  ���}�Z_����=+ F��(�dټ<��m�|Ä��  À�; �$�Պlٹ,+����u0���^u$ �T�2�R�\����i���   0�x/���Hr>eJ�v�Ql��ɹ����tż��  È�; 0��I��᏶��{A������}Zu$ ����{��/�ݛ��   @kSp�z(3x���: joo˶[���{��^�U f��KZ�tf��ޛ�O��?9�3��}�Тzz<�MRPv��   Z�z;�N#�K� �vEQd���y��s�M��� S� �ת�kٲsYVv�����`�#eiQ`tk�L�º�಻�   h*�|W}+�� �4u��|��[�|����  Ü�; �&N���-�7/������������0Q���'g�\wo�ԫ�   |gE�4��������B��s ���=[w�ɝ�lI�n, �v
� �e��hz��O��sO���r8gN��: �J#eΦ��4��%iK-�X~  ��Fŝo�3��n��K+�"���˃��S&V A��+R�ٲsY�v/ȯ~z8�=q$e�  +S�\�s�I��S�޻�^��;   w
�T�9n�c���r�7���̒�� �@
� �w�9�#���;]�����޼��UG`X��= ڷ��,�'�'=   ���Xh����3�=�n]���ژz�Vu `�Rp �ʬ�S�w���rh����_ȩ/�T	�a�L��)s>ə^w�W   H��>5��e��J; W�(�,Y6/>t[&�0��8 ��� \��(ҵqA����_���9���7��\��  `�)R�7�
V��z�gL����;ͪ:
 �"��kf��1y��7g��%��?ߗ7O�_u$ F�����Җ\(�   CÇ�[S�B��J; Wkܸ��uGw��Z�Z�Vu ��(� ��ͳ���xO^{���͟���~^u$ F��4��{�ݽH[o�  ������4z�_j��S�ղj��<��9nL�q ��� \7KW���%3���/片_ʹs=��E �.^w��Hۅһ�   p-y�=2���F����p ��y�ܜ���ݙ9�ƪ�  -L� ������}��߲(���9�����7��)sv�!�fѽva�݁x   `4XhoD���a�䉹��[�ս��( �(�� �I�;��m��͋�؟��|Tu$ ZNO���'g����S(�  ��Jz�XhoT���ўm���woN�^�: 0J(� Cj�����?�;������ۃ����UG�%�)s>e�'9�"�$m������  ��x�<|���J; \_EQdɲyy��2��	U� Fw `�E����l��<������4N�
���<�{6=��.�����   '�e����,��иyִ<�2o�̪�  ���; P�������޺8?���9~�dՑ 5zz��&)R�6���   ܇Z�B{s�]��*L�0.�ߵ9[���:
 0�)� ��>sr~��n��#��'�/����H �*eoٽo߽�]w�'iO�>   p͕�O��� UikkK�敹��m��P' ��	 0l,\2#�����s��������: �R�2�S�|�3)RKz��/�  ��q��޼��@�������;��;S�N�: ��� �J�^K���Y�5/���<����\@u���8�\����\y��  @+�z�ꔽ�f�]���f֬i��n������ �
� ��4��#{�[�����=����H Ы����}�����  ��տή��p5i���sc��X]u ���� k7N���~�#�.����`N��QՑ �"}���)���'���"�X�  `d�z���ڛ�
� _�ٴuu�gS::ګ� ����aᒙ��?�;��������|���#�W4c�$����H�ڀu�z��   ಩�_J��퍪����jY�ra����|Ä��  \w `�(�"]d�ڹy�W���_����@ `8+{��{z�)��+�  0\��7�=���f� F��s������[fT ��(� #N{G[vߵ:]��u0/z+e�ԯ �eʜO����E��һ   T���k�F�ս���4u���u߶��ZTu ��D� �n�:>�xG�~���/���W	 �P�{��'e����{�   �>����H7~\g��Z�[o_�z�Vu ��L� �fϻ1��{��Ko�'��@>��gUG��hp�HR��w   ��%��µ�v ZC[[=]����sܘ��  \5w �e,]9;��ݜ����{8_|~��H pU��ٿ��^��"�xY   ߤ��^���@+�E��\�{ܑ)S'V ��q$ h)�z-�[g��[��#���_����V�V�\xo��7�%i�-�ג8�,   �Q�{Qh`t�={z�����e�̪�  \s
� @K�Ӟ�w���-����^��g��,� ��4؟�pȾ���\x�[z  �V�,�7?�Hy�� ��nȝ�nɚ��UG �n���6irg�hS��.������8�nՑ �*/�~�|�#��
�$Eu  �;�x�ݙ;]Ə�̶�]�u���j��	 �6w `T�y����?�#Ǐ������y�7W	 �H�����{������»�;   �M��i.�+�0:ut�g�U�s�tt�z ��g= ���pɌ��ޓ���#?=��?;]u$ be����p���{}�u��x   �R���I����/ ��V�ղj����;;2qҸ��  )w `ԩՊlܶ8]����G��/^̙�窎 �)/��5)���\zoK��   �J�*{�kR ��(�,X4;�=xkf�|c�q  *�� �Z�m�q��lز(O<�R�y�՜?�@
 �)���}����{qa�VU<   F����Ph�� �2k������,\<��(  �Rp F��q�sߺlޱ4����x�XX `����PA��H=Tz   �� p�n���q���]���(  Â�; @�I7���m��[��џ�����H 0�����ދޒ{��{RT  ���:; \���e��]�yǺ�jFD  �(���    IDAT \d���y��;�e�����[����H 0�)ӓXyoޛ�"mi��  �����?� \��c:�q���q��tt�W `�Qp �s�ߔ?��=y��[���ʇ����H 0�<}��I2`��  ��o��'��v�� p5����Z�,w߿-�Ə�: ���� ���Ȫ�yY�zN>w<���|��U����O�[ro��7��v�  �R�5Z�Y����F�L#g� -�^�e�ʅ����2eb�q  �=w ��P��ҽuq֬�%O=�j����9{�|ձ ��)s������楸���  p������ڭ���WE/��{g{�ϜZu �C� �
t�i�����K���/���_˹s=U���ҷ�޼ݧ��^KRORWy  �e�4K��� 0�fϙ�{ؑ�fU `�Qp �:�ud�}���ey�ᗲ��c9^� ��F�4U0���Eo��Y|  �������3}���wkV�^Pu �K� �*L�ܙ{Нm����_���K�� ��������u�ڀk  �����ƀuv�M@U�L����m���� 0�)� \7L���ڔͷ.ͣ?{!/z+e�` ��RG�b@ٽH齨(!  ���x�]� ��ɓ'd��y۪�j7  �w �kh���y��;�����|N}��H 0ʕ_SzXvWz  �ev Ə�-;�f���V�: @KQp �fϻ1����#���|�y냪# ����%��k)RO���;  p=5R^(�7zK��� 0��ӑ�-�r�ݛ2fL{�q  Z��; �u�pɌ,���r�Ȼ��_��w>�: pI���]xt��{_�]�  �r}���evev Y��۲v���}���?��8  -M� `,\2#��rw�=����|��UG .CsI�1�r�Wv�+���  h�� m�\� �D��mY�nI����L�8��8  ���; ��Պtm\���o���#?{!}�yձ �+�Wzo���Wx�ԣ�  ���C�}���� ���^�g������2eb�q  Fw �!V��.�>w<����|�ɩ�c W�齿�^�H�Xy��  #W��^^(��/� ��V�eي������U� �� *R��ҽuq�mZ����#?}!�}�eձ �k��-�4U^�%���{����  P�������Uvev he�Z-���ͽl���S�� 0�)� T���v����X��K����U� ��f9&i�e�5���+�}�w  ��({���������Ѣ(�,\4'w߿-��L�:  Qp 6�;ڲe粬߼0�=y4�����lձ �!�W�\z/R��"�޵����;  \��{�9w9�> 0ZE�g���g���U� ` w �a�cL{vܾ"��/�sO�c�x1gN��: P�2e�K�=)��|��Pr�[y�x  F��s�F�ϣ����EgO F��(2w���u���_8��8  \��; �0�1�-;n_�[���_�S���� $�[{O�N���{q���� @+*{���`h#�D�]� �3{������,X�� 0�)� s��:�����޶8O���<�䑜?�Su, `Xj\(���x�����"��  }�q/�V[ .OQ�{ˌ�{K.�Su  .��; �1a�������z��<���� �e*S�'IOａ..��{�+� 0��+�/�y  �ά��r���e�UG �
(� �0�Ə��Vgӎ%�� �U���{����  \c����n[d ��f�}k/�Wu  �w �J� �^�J����~�������~  ��A%�*� \?��  �A� `�St �J9�bE����w ���H�2�F6�� EQd��MY�ln�q  �� Z��; P�2�+��h�����,��3p ��YV�� ?EQdμ�s��,Z�� �J� Z��; 0��/y�����I�����ex  �R��^^�Xb�� /��  �O� �E,�?��+y���r����c ��K�\�6uq���� �������Aľ�  �[Q��`V�gK�/���8  \G
�  -n��1���]��������<��K���٪c |�K�ߛ��z�ڀ��z� ���+� F��(2���-Y�hV�q  
�  �Ę���q��lھ8�=�'~9�}�eձ  �H_�}���.^~�/�+� ��}��h�]� h%�Z-���ɝ�lɜ�ӫ� �Rp e:ƴg��eٰeQ�?s,O��|�ɩ�c \#�^~o*R��f齯�^�8 �p0����v `4�+��ޭ�5gZ�q  ���; �(��і-;�e��%y��y��/���~Vu, ���-�]���,�7���{�	�� pu�$�v ��hk�g�����͙6}J�q  ���; �(W��ҵqAV��%/x#����|�; 0ڔIo�,��H���b��{�m ���y��{�c�J� 7��mY�r~�ܳ%7M���8  
�  $�/��힟���G~�B����c ��Z��+�)R�^g�5 �*/��_��� .G{{[�t-ɞ{�d���U� `Qp `��(��k^V�����:���Ŝ|磪c s�r[�#\x�t! �����K�{*M �
Ǝ�u�Ks��6e��Ϊ�  0)� pIEQd�ڹY�vn�<�~��9~�dձ  F�f)�
��k�E��Z��R&)R�� К��6�\Y�/��i��Pb �z7~l6n^��wvg�؎��  0�)� ��-�����������/����,� ���W���H��[��~_��~��c��O  �ڛ0q\�7���=���h�:  #��;  �mނi��`Z����y�W/�o��p� `�4�y5��\�X~�/�+�02.�7R\����	 ��f��Iٴmu��\��6g� ��)� p�f�|C~��m���y��W���9��W�  �K�=\���5���{1�6 \{��z���]]We ަϘ���e����jU� `Rp �;�a�������sU�=u4O=�JΜ>Wu,  .���7�J�M����u�D`�+{�.)S\�;�a����  ���(2gތ�cC��ZPu  F8w  �ڄ�c����ٺkY�>u4O<�R�<u��X  \兺b�"|��K).���-�,�
�}�y F��K����$Š��o��  h%EQd���s�]��p��  �"� �fƌmώ�Wd�%��̱<��+���SU� `�.<�?�U�z�Ņ�Zｾ�}%���x �^yaY����rz_��o���o�� 0���,\<'{�ݒ�s�W ��� �5��і-;�e��%9���<��+y��O�� �02�\y�_��"E�e�b������ ���g��rz9��^xl�
;  |7�Y�nIn۳1S�N�:  -J� ��^�e��Y�iA���N�y��?�nձ  ���̞��~9�o�}`��}|`����Z��Zyтz��K�}�7ҿ�n; ����9&k�/�wm��	�U� ��)� p�E��+gg���9��Gy��W�7�h8 ��4� ڸ�W�ͥ����/^�/R^����s�Z��ǚ����}  0�L�2)�����[פ�]� ���'  Cj��)�᏶嶻����^́g��ܹ��c �ER��w|��%�⢲|ٻ _~e5����<��Rz���+���7��b@M  Z��S�cWW�oZ�Z���_   א�;  ��r������ڳ*{�<�g5_�:[u,  �F.]��x��r���J��-�7M��E�b�?��k���O�F���W�%��sQQ�Oc��$W�]x9�  �E���ff���l����  0�)� P���f�]��m��x�x�|�|��c �0Q~��;���ۗ��?pU~��������|�����)��i-��o\��IҸ�W��,�����#׮B��  _U�ײp��y��̙7��8  �� ���1�=[v.���K���Γ�z%��Aձ  �E}�P�u�ߋ����%��{}��f��6 ��5��)�݂�w+�_�W}�B�������e.�D1��������5�v��|۟��  �ט1Y�zav���M�n�:  \�� ��R�ײ�k^V���c���S����GNV  �J_�A��i%h  �+3q��to^�[w����1U� ��Pp `X*�"��ߜ��o��w>��'�����s��WOm     �7���ٸeU��\���z�q  �k)� 0�͜5%�?�)�ݽ&��:�g5_�:[u,     �a�(�̙7#��ؐ�T  .��;  #Ƅ�c����ٶ{Yx#O?�j~�ާU�     V���Y��������9kZ�q  ��(� 0�t�iO���ٰeQ���N�y��?�nձ      *��9&k����ug��	U� ��D� ��(�,]9;KW��ɷ?�S�����F��:     ���z�lܲ*[o]������  �UQp �%̜=%?�Ѷ�~���}�h�=},��<[u,     ��(��<��lپ&6�HQUG �kB� ��r��	�sߺ�sU�=}4�=y4�yձ      �����,]>/��ؐ9sgT  �9w  ZҘ���~ۊl۽<G^~'�<�j�y��X      ���	�Y�nIv޾!�&��:  \7
�  ���(�t��,]9;�y���{�h�;�s�z��     �n�ir6nY�m;צ��^u  ��� 5n�=%�?�)�ݽ&��=�g-�~r��X      ��j��2f�����UREՑ  `�(� 0�L�86;n_�����~��y%o��Aձ     �Qn�؎,_9?��ܘ�3�T  *�� ��U�ײ�k^Vu�˛'�ϳ������F��:     0�L�:1�7.϶�]��Su  ���;  $��`Z�-���>�<�<�Z>w<gN��:     Т����[fd���Y�nIj�ZՑ  `XPp ���8!�<�!wܳ6���g-����X     @�hoo���d�ݙ5gZ�q  `�Qp �K�Ӗӽuq�<�~�}���|��4e��     �h���Y�~iv޾>��wV  �-w  ��L˼����g��G���c���٪c     �\Q�3wz�ܺ6k�-N�V�:  {
�  p���8!{�[���^����}5'����X     �03vlG���������Y7U  Fw  �Bmm�tm\����_��{5/|3==���     �z�tmX�m;�2n�ت�  ����  W��9S��m˞���о������ONU     "�Z-�,�9���ʚu�SEՑ  `DSp �k`���}E��\����<������X     �u2nܘ��Z��rӴ��  -C�  ����z�6.H��9��G������zΝ=_u4     ��6}J6n]�M[W�����8  �r� �:�9{J�hS�w���p��<��ky��'U�     �P{{[-�����`���  @KSp ��l���to]��������~���F��     �o0��I�ڰ4�n]�q�;��  ���;  �y�eނi����y~�<��k���SU�     z��̽eF�ݺ6+�,JQUG �QE�  *0a���}E��^�����g{5'����,��     ��ĉ�j��ؽ.S�N�:  �Z
�  P�Z��ҕ��t��|��ϲ��c��̱|y�l��     ��E��gݘ��Vg�����UG �QO�  ���7M̞��e��V煃of��G���T     Z���c�lՂlݱ&�fO�:  0��;  3�mY�ya�o^����$��=a�     �RQ�y�Ԭ۸<���N{��  G�� �06m���o]n�{m^}������?�nձ     `�����+nɶ�k2g�̪�   �B�  F���ZVu�˪�yy��O����9���=s��h     0�\k߸eeƌ�:  p�� `��6cr��Aw+����O�ɷ?�:     TnlgG����m;�f��U�  �w  �:ƴ�{��to]������{�Xx#gϜ�:     k�  �Z� ��<gj�hj�w����z�?s̪;     -��sL����-����  -D�  ZȘ��ٴ}I6m_��N~�C�Nd�3��婳UG    ��f�  Z��;  ���3'g�}�r��k��og��Gs��{)˲�h     pEƏ���nɎ]]�5gz�q  ��H�  Z\[[=���eU׼|���rx�9��|�񩪣    �ת�k�{ˌto^�5���M�  F�� `�z���kuv�Y�׏���O�ˇ�J�a�    ��a���Y�za��\�o���8  �Sp �Q�V+�pɌ,\2#�}�e�{=��>��>���h     �B���̛?3뺗�k���j��#  Qp �Qn���}E�߶<'�����+/�:���T    �7m�Y�~I6m]�	�W  � �$IQY�tf.���_�͋Ͽ�����[����h     ����1Y�xv6n]��K�(��#  È�;  �c;;ҽuq��.���~������{O���NW    ��^����7eͺ�Z{GG{Ց  �aJ�  �F�fLΞ���{��������y�_���Qu4     ���7LȊU���5�iڔ��   #��;  pYj�"����%3�婳y�Л��䑜|�㪣    0�tt�e��9ٴue�,�%�Z��H  ���  \��q�޺8�[罓��о9�����L��     �@�(2����^���+��9��H  ���  \��3'g�}�r��k���r��9q�ݔeYu4     ��ɓ�g嚅ٴmu�ϘZu  �(�  �D[[-��ߒ��o�g�~���3�;���|\u4     �����,\<'뺗e嚅��jUG  Z��;  p�M�ԙ-;�e��ey��'9��D��{"�v��h     |�z-7Ͼ)���{�tv��:  Т� ��j����sߺ�qoW^?�^��{</z+���T    �o1��IY�zA�7���7V  � �!Q�Y�dF.��{НW_|;���ȉ��,˪�    �kܸ1Y�l^6m]��g�(��#  ���;  0��vv�k�tm\�O>�"/|3��>��>���h     �R[��9�����K��{Y::ګ�  �R
�  @�&O�����ۖ������'���r�����    ��ZQdƬ�Y�vq6nY���U	  @�  ����E�3����{�r����о����NOO��x     -c��bՂlڶ23f�Tu  �A� �a�����+gg���9��ټ���9��DN}/eYV    `�7~L/���-+�`���j��#  \��;  0����H���ڸ �||*�~+�;���|\u4    �a���-so���K�f�ⴷ�W	  �[)�  #���e��eٲsY�;�I^>�V�=��?���h     �B�^�ͳo����޼"��c��  pE� �i��ə>srv}oU�z��9����p���9}��h     C�(��4mrV�Y�M[W�)���  �)�  #ZQ��`Z���:����w�$��^��-��ƀز +��s�k���:&"��j�AO�C���З9���LN�TOgW�]I�$�l$�al�Y�,ˋ�o.� ͒,�����zE�s,��y���/�w�Ͽ�����ؙ������s���4=    �Y�Ȫ���X�zv6oY��  �{B�  ,���|�|��޸���>�����ཱི�tj��     ~����ٵw{�zf_۹9���'  �Sw  `QZ�| ��ٙ���̍�[?z*o��G9����*v    �+���Gs����pg��vӓ   ��;  ��-_1��ve�]��2������ۧr�䥦�    |�����s��<���88�����'  <w  `IZ�"��to����|za*�o�α7O��ך�    ,q}���ƌ<�+O������3cQ    IDAT�  Xz�  ���~�P~�ˡ��s��T�=z:o�(�����    ,}�V6=�Hޕ���g��eMO  h��   ɆMCٰi(�ߍ���K{�TƏ����٦�    �L_��-��g���<��ެ\��$  ��!p  �K)%�w������W���n�����{�t�]���<    `�j�[ټe]����S����ꇛ�  Г�   b���c�>����    �wk�[ٴe]��ߑ'G�d��MO  �yw  ������_�O���bw    ��Z�d��59p�qQ;  ��A�  ��Z����u*ק��    �ԴJɺ�CٻGF�ߟ��6=	  `��  �w�����щ�{�t�{�Lfo�jz    p��Z�lڲ6�����d�#k��  �(�  �v��]��d׾-��_=��e��Oe����    �еۭ�߸:�vo����ˆ�뚞  ���  /����<��'���{�����L��    �﩯�ʦ-�d�yrtO֬jz  ��&p  ��J�r�~���?��8��.]kz    ��v+���˞�;��3{E�   ��  �*�d�ֵټum~�˃�x~*�=�w��8�.^mz    ,Y}ٺ}C��ߑ'�ޓ��W6=	  `I�  4hæ�l�4������Or��gMO   �Eoࡾlݶ!牧�dŊ�MO  X��   =�����ūy�3y���;3�Zk��    `QX�rYvo����9pp8=4��$   �"p  �A�lX�����������l>x�\Ə�·���\��y    ��>�<�wlΡû�odG�����  �� p  �q+���3;s�����q+?����w����;M�   ��SJ�굃�9�h�xjWv>�5�v��Y   |w  �d��ޞ���s��\>:q>������3��6��<    hL���]�*{�n���=���ƔR��  �$p  X�����s���9�h����L�||)co�����ԕ���   �}��neӖuٳG?�;k׭�  ,pw  �E��*پs}��\�����s��d�=v:��?���SM�   �{fٲ�lݾ!�Fv����\��$   �!�;  �"SJɖmk�e����u8W>�·������|�����u��    ?���l۱)�G�3���y衁�'  p��  ��k3�®���+�7n��������޸��<    ��V)Y�~Uߵ-#O籝[�n���  � p  XB�-����9�=�N͙�/���'y�3��鵦�   ���ۭl޲.��ٖCO���M�RJiz   ��  `�j�J��\��;�����\<?����cgr��˩�6=   �EnŊ��u���ٿ=gժ���  @��   $I6lʆMCy��ϵ�7���'9>�IN~p!�o�5=   �E���5k���Gs����ڳ=}}�   ��_%  �5�Z�g~�+��dWnߞ�铗��ؙ��Ι\�2��<    �v��M[�eמ�9ph8[ݘRJӳ   �Qw   �U;û7fx�����f4���s|�{���O37�iz"    =f��lݶ!{�?��'���ʦ'  �@�  �A֬��?ݛ��77fne������lfo�jz    h����Wex���޳-��=��>I   ?���  �϶|�@Fo�����tj.�����y���;�Y��    ���˖-�d���9xx8�Y�RJӳ   X��   ��V��k�y����3yy:'����&.�ΝN�   �J)Y�fe��؜}vd�hz   ���  ��bͺ�<�Ҟ<�Ҟܾ=��'/e���?�O/L5=   ���M����=[s������W�  ���   �w����ޘ����d&/Og���|t�BN�w6�n�iz"    �V���ٵ���ّ�˗5=	  �%D�  ��f�`F������t�}�ą�;�Y��    ������y�#�1�9�Fvfˣ�n���  �%p  �Qw_wO�+�]χ�Ϲ�   p��R�z�`�mۘ]{�g�����  �3�   ���kWf��u�;w:95q1'�;����s��T��    �e���e��<�{[���Ȇ��RJiz   |��  �������M޳)I2}m6O\�G'.���'�v�F�   zS���]�*û�f��my|϶4=   ���  �c��e9�=#����gr���L��������ħ���4=   �1����趍��hF����U��  ���  X�J)ټum6o]����ܾu'�?�����2q�BΝ���    �U_;�6���{�f�yt�ƴ��g  ��"p  `Q�����޽1I2yy:'������q��    ?N)�k֮*�۔]{�e�Ȏ,_���Y   pO	�  X�֬��]}aW:��ON]·����ɩ˙��4=   �{�|RS�)�����~t���K)��Q   p��  X�Z��m;ɶ���<�;��r��L?��r����Z��	   ��:US�I�)���ȅ#In'ɮ�;�Wq;   ���  �%������3�{c����lN~x1�����ϕϦ^   ,!7K:�%�WK��~&�~��Fӣ   �)w   �����2rx{FoO�L^��ĉ�y�3�}�޹$Y��@   `1�K:'y=��ͥ�K��oz   �
�;   |Śu�]�+�/��������*'����������I�7�   X0j7h/�O:��d�����>�~   |��   ���sW�7�}�[��\=�I�EI�EMy)ɲ�G   =�^L�?��?����[9�~�Nӫ   `!�  ��ʝ��H��o��,8�F��8��e��f7   V���cI��\n��vο��vӫ   `!�  ���ڍk���}�1O���C?i��$/%y.I�  �{��^�ɱ��c��on����jz   ,w   ��.���$��Y�����xa>x�E����'   ?PI����$��$��9��In6�   #�;   �G�fl:w�ybC2�Ӥ��$?Kr0I�ɍ   ���t>���I�oI����3�E�   ��   �������y$/>|#������R���78   ���ze�B�?ƅv   h��   t)�^�]��gdp&+^h���t^�)�d�ё   ��ԋ�����9�F�[M�   �   �S>��t�
�7払3�*ɋ%�5�$˚�   O��ԣI^+�����7��nz   �uw   �ar�z��Ϳ�ݒ�WS_H��VZ?���'lt$   ��N�9Y����Z3��o�»I�   |7�;   , gsd&�?̿$�j�侒���TR~^�mN  ��fR?J�j�j2�n���t�   �pw   X�^��N��}�.I���pM}�&/&��$���&W  ��So���5�H������'3�^   �w   Xd���D��$�N��y~c+��KʋI^J�\��'  ��VR���XI�}��+39�J��w   ���   ��y�B��̿������_$�/�W��\��&7  ����s�&o�R^������sG��jz   �`�  `��,�_M���/ɯڃ9���:���KI�')ͭ  `i��%���r�&o$�{3�N$�4�   h��   ���禓�t߯�de����ܳ%�Ѥ�bMy)ɲFg  �ԋI}�$o��Wfr�$ך^   ��;   �5����$��I~�7���k�K5u����$ۛ�  @ϻ�t>�i�%�՚[�ﭜ=�d��a   @��   ��+w��#�$ɪ<�+i�$�/t�J�D��  �%�^H�xI��t�q&W^M�]nz   �����   ���j��A�����OF��R����{RF�hp"   ��lRO֔���Z�쿿���uv   �G�   �ȑ�_��"Omi����F�΋���(ɊG  �g��z���V���ɩ���jӫ   ��G�   �73y�l��I~���W�����J�ɋI})ɾ$��V  �S%�X��k�%��0�S%�M   ?�;   � �<7����~�$�����:)ϖ�g��l�M��  X:��򇤾QS�h���S��GM�   �.�;   Ш�y�$?��$+�Ԗv�hIk���&y!�#Mm  X$�$9��#%�HM�\��[M   ���   �93y�l��I~��g�G�Iy1�K5y�$+	  ��&���c��#�k7�   �m�   �������}+s�`+s�%��$�&9�����   ���$�TSߨi��,��W�5=
   ���   �+w�'o���]��������RG;��%M�-kn'  �=w.ɑ�e�Α�;�O��Ż�`��a    ?��   XD�ܞN��}��~&z  ������M��O�   p��  �E�����ޯD�O'Y��N  �/��Iy�Z�\jz   ��$p   ��W�|ӥ���P'y��<YS�Lr8�`s; �E�N�w��VI��N�fꛓ92��0   ��	�   �$GnO%H�}aE���N-i����t��ond"  �M'y?�����9�p�92��0   �^$p   �3y�l��I~��gC9�������G�e4ɾ$��v  =a2�xM��R�tR�L�w�t���k�l   X�    ?�T�M&���K�<�����%y��>���IF�,kj'  p��%��$o�ԷJZo�I}s&G�5=   `��   ����|%zO~����:�)i�&�@�F����f�  ?�T�w�2VR�krdEn�y!G�7=   `1�   �7/�M%��|���<��v�<���HIF�N2��R   sI>N2^R�tRǒ��t�OR���k��   X�    �gy�j�v�=�Uy��N��R��ɡ$O$��� �^�TRޮ�Mr���ʪ��٦�   ,uw   ��й��N$9������#�Y���:ZS$Ir �w  �>�&9���%u����Tޘhz    �L�   ���nM'c�/���P'uWMk��:�J=PS&���N  hԭ$�d,)�Ա�5>�7�M�iz    ߟ�   `�̑�$G�߯?�|e�ݔ�`;sk�H�C�^|���  po�N�~I뤾SR�Jr�j�(yy��q    �xw   �E�z�8��|�����P��d`$�K�#��G�lnd(  |�/.��d����tƦ�j,ye��_��>   ��C�   �L��d��Ϳ/�К���5RS$I����$��/ `����DI&�2�IKZ�����    K��   `	�ߏ̿/�Γ��R�'�Iݗԑ��K�X�V[ X�>MʻI���5��߽���|��`�   �3�    |͕�u%�k��.#CY������H�pIg��<�dCS ����.����:�I{"�;������   �0�   ��nM%����3C9�&��i���%��H��I�M� ྘L2����d"i�Og�{��sM�   `a�   pOL��d�#��.#�Y�;��[R�&ٓd��s� �7M��$'jʉ�����v���92����ƃ�   �"%p   �>�5��������s��s�$�I.�ה�$�z) �s+ə�:�I/�c��'�����q2I��}    ,Aw    ��쟊߇rhM�?<�2�y��ԑ$�=�  ��$�K�DMk���ϥ5&b   �W	�   �IS96�������<���]%sÝ��<���x�Mz+ @î��Ò:��Ú�DM��/�é<v*yy��    �}	�   Xp�s�b��I���v�CCY��d�����_��ݷ�$+�^ �{`2�DI&j2�ԉN���?JR���~� 7   ��&p   `����T2����_�W热wR/��K�Κ�#��$�T �?���dRN�ԉV���|�I��Ϊ��Wf�    ��   �%��+����������[�lN7�/t2 �X�L�II��iM$u�v/��k�u�ۯ�   ��!p   �/|���䑼�����h��();;);Kꎒ�Ɏ$��\ ���&��&'[�G59YSO�RNΥ����~��    ��   �{��W�%96���ϗ���;�p;uKM�ܽ��)�I�%�p��{h2ɹ�z�O\`?����F    X��    pϼ2�m��d(��$��s)ídKM6�d�&�I�$���� ����L�s%9[���N$9�J��g����    ���    � M��d�#��kɋ�ff[;����-5e{Iy4��&ٞn��N��&3%9��$gJ��N�ْzz.�3%������w    ]w    �!��a��ߟ��yx]��o����ǒ��h h�l�����zI�u���ԉ۩�f��$��    ��$p   �烛3ݘ�l��%�dd`yVl�˝�IkcIٚԍ5ٚԍIٚdc�n7 |o�I�$�BM9S�%�LR/t�9SҾ�"��\���M    �-�;    ,Jc�n$��}��{���_���X䦒�����0    x��    ��}�>ʡ5sY�����&�[ɖ�����nI�9ɖtc��}@�M2��Y�\R'�r�$�:�ْ��iM�u���~���`�u    X��    ��2�c������}+2�!io�K6���I6u/·�'y��n,��$�$Yv_��C�%�4ɥ$�JʅN:�&�Ӥ\(��d�b;�ܕ,���v��    �""p    �W��t���M��w�O����V���ds;uKR�|�:�������`��Lrn��_\X���>9����;�3�u!yy��    �%p    �ڍ��F�A��w}�����Lk]+Y��YWRIʺ$k�����.)k���뭽���g�&�%����V�gI�rR/w?���s��^n%�&sd��)�ǿ�    p��   ��l��$�Ir�|[k0O�+i�KZk��uI֕��$uM'uMIku�r|V�{)���.��`����%�+I&kr��2Yӹ�����L��rҾ��˝�}6�k��n6�    ��    KAg:o~������Z�5kJ�֔��%�5I]�I]��V�n?T��N��$������� =a6���7UR��ԫI��d��ԯ��X�f�JMk��֕��L~���f�    �.�;    �������|���Q�rhuI{�vZ�Z)�JʪN����*)kJ�Ý�U�q�ʒ����2�+�&J�"��Ïq'ɵt����\/��zM�����$Wjr��z��u��^k�^Mړ�t�^���d�֟;�ƽ��     ,Rw    ���N��d��{��j��Э,�K]�Jgp�{=~eMV�d()�5YY�����duMJ���p~ ���K����$���>�����g�m��%��|�~�$�kr=)��Ε�2[���N�d���Դ��S�v��v�L2;9�3�7���    �}�    ��=��fm�_u;wZi��˝e��si=\S�Z�֤�������Ǘ�$�t/�'���V������&�K겚����������W%i�����{ֽ���mM%�$I�^7�K��nH^�Z�=5e�{��$s5�)�͒z����j��RӚL��ܹr'�ݗ�k�ӹџ[�S9�ş    ���?,      I�Y^�:��KM�ؘ'V�v���VZ+2�P��%�ۙ�������|�{K�ꤖ���/JJ+ߡ�,�����}�����SM��Թ/oj]�޹��V굹���Y;s�%��$wҞ��Knwj榺?n�+y�ʏ��     ��$p    ��\���I�����&�      �w^�          �A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           @�	�    IDAT��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�          ��           ��;           =A�          @O�     ���k�    ������8    X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X�          X���;H� �^v��X��$"\!2_з��52         @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�          H�          � p           A�          @��          ��;           	w           �           $�   ��R�  �IDAT       H�          � p           A�          @��          ��;           	w           �           $�          H�          � p  �33o�        ��;   <�{�=     �W:8 ��v   x&p    ����z{ ���  �3�;     ��� p�;   <�   33o�  Qw ��� ��g��    ෽�Ϸg �(�; \D� �\ <��;   �������  �Y�"w `��~�=  ��  ����� \X w� X3c! g�   @�}> ����E� �Zk�|{  �rn   J|� �ޟo�  �;^� >i
 fƹ   (�z{  �r�; \ċz `-7� ����B   (qa ����E� �Z� �Ĺ   (q�; ̌� .�E= �����̼=   ��6  ��@� ��  ���
w   ��> ��F�E�� ky& �'w   ��> \X wq� ��L  O,�  ��| 8��| ���/ ��Z��  �,�  ���� �� wq� ��L  G.|   J�{ ��o$ \�kd�z�4�    IEND�B`�PK
     uK\���'  �'  /   images/16bd2965-d7b7-4d97-b402-ac1747e7568c.png�PNG

   IHDR   d   �   ��P�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ' IDATx��}	�gy�[���ܷ��h���˒lɖ�����l����`'\��@�	K6����s�,` �p6|�l�-!K�!ɲ.��h���������kzf���R�z����{�����J.jp�|�4��"YK��d�J�&�Z�J���e�"I�DI�I�I�H.��#9mJ��\'��n\\RB� ��ʊ���&�m�0)�N�2�'N��l��&I�y�#$H^�$*Q�Z/%9�NH%n'�VՓ��;In��7�Lp�)|�߇$���$O��%�v��I��BxfY/n�ɴ�2�H�Fr���� 7���|�d��Y���!�Q2}_�e5KNH%n$�(#�P2�gw���t���8�AS8�����nM�[�B+� .鉗��J� <�b�Pɍ�w�	@�~H�X4��;%�SI�^8�}��$�J�U��u��٫�f�'b^�R`ф0|�]�
/�[M����݀�.Z�.�غP|F�.�9��G��M�n.���J���T�Μԑ��Ht$�)j��
$E��h�|��^:��������:�n{Ƣ�Y!L��j�� �����[��/��w,�x��-I�Fj�����·�?j�}��񡜖��<�z5hn.�
�$DgBRDB"�X,�h8��ij�Q����D0�"L�5�UPTA���w�=�;��_�����5�
�,��"���?
$����d�D���G�ŧߣ�����*Ѳ��+*Q][�ʊ
���������0."�ԩ�vo�0�T��+�"�H"�!�"9Ә���P�A��12B$�4�)�v�ޮ���������i�K?!�dBd��D����ÚϪ(g��,�8l�J�Z�*�f}-:�ա��uu����FyY9�%�P>+��-�5r#��[������W�SDP��	arj��q��}&�s'�1�B�Ѕk,�jxK���w������=���X��MH�*,U������7�\J�`ե���ݬ����5�smV47����,���`�v��u�Y��@!W�#K󣾮+��a˶ ��}v'������s�`1� ):�O/:�G�Zr��Tk)��l2�y
j�T��[��R\�V]X���njA�5�hiiEuUY�;�|n���d[NeE�*���ڎ��ؼu g_���8s,�]����N��&��G��Gd9�0DǀR���KH������IW)�G�
�+;���-�ظ��m+QUU�v'��/,�c�X_�@VZ���+ѵ�"N����.���d	���8����Cd)7ҝ=@��}kE�2'!/P�;�^xf���J!v�?��n-��<n�pK+v�Z���5�%��D�2f��˃l�a���XM�ۂήs8��^�Ӈh<Y����h��tQwӒA^>)���B�Ue"����������z/nt�!���©劦r���.\�z������(�j�Z���FSS#�V�į?���HD�E,�rYʯ�����/������������,�w\{��R��������'^�?z
�_:�(�s�?W��;L�Zʚ����47����� m�+��X�j���*��O�����"I1)�7PL�%-���u^3)3y��_�2���������m���������^<&�y��=^�M�����ش��{6o�$2�7ِ�,E��b�M;PQ��c�|Ǐ�M
�`�O� ��������)3������.�*���"Ctr�M�93�ߵ�o݌����b���9OⵃǄո��M��;�ހ��6BsioX2����k�֭2#��q�Ѣݗ$%�E>�'��I�*�]!����E46�0P�Gd��߁]<&�ׯ����w�������©W�e\K�l���W�^TJ�7m��^�o�����"Ia���a���!����[I���c��������D���;E��l�u#Vol��u�[�)Ȱs�^(���7v�w��?|s?�&�E���p��#�w����A^�MJ������ ���U��^h$d��?�ʖ���J��|0)ܛp�έ���g���聘��'*��]gS��;�"94"]U"�м~�WQ�P*�t�:x �T�5+.[�w)���-���؁���UA��(�u��$iY� ��ػx|����R.����T���`U[�UA�����&���[q��n$z���~�s-t���C�Yk��#)Q���ԫ���R/�b.�8��r�0�+�U�A�{��ذ�8��/*��!]�VR�3�q@�/�4UX1�1Z�V��(�q�0�wM55W���
�|�}y��X"���3x��GI���h�:t����z1*olx ^%��~fU� E:�v[V��PX���U؉!����$_'	kbG�oC��L�ﰼ��� ��>\�TH�)���X���Cgf�Nʅ���\|s��O59��|���R�ɒZ��@%�&�=T"4�˸���h�V�y�t�{�����������j"+��DF�R��)!�`6p磒J�B�j����Ew�0�-+X4f���ȑ���f^��e���������)�S�`�ӕ �5�p��$�Ť�k�� ��d'�j�e�v!��S���:Z��(0% \��0!^�G�tLH�PĜ�4vq��vy@i���i8.�MQ��0�Js4��]VW�U.u��!��TW%Bd!suS��jh:&fL.]LH�8 rS^M)"�%�4_bSc����'G�&7�EV�!�z���ȸa��	���171ފ��zq����?=(fa�$Br|W��9Yއ	�+9��j꡸�"���b�N�-a���K�+=�V����6M��m�������jxHb�qj%Wg=�!Ο3K#��)7��e�KI�`T!#ѹ��_�X��	�jw����1�S1xKJ2�#��[D�yLvh>�F����S�Ԏ���HDCW]�ΏC��cϳ�J�ٱ�[��®)���'07�.���Y-�/7�W���뇮�����ˋK�k�y��r	!����M�k��hH�sX	��l^��h?"�!Q�\�x4=܃g~q��쐳�gfL3��qD��|"���<VY�4o܁���!�)GW���������q=I�,�]q��Ω���'�T��h��^)K���֒����^|�޴��[_��"�����q��`�������l�3	!���e�Z�Js.���=&�4�Lc�S/��>�C�9��T��o�}�!N|���dp���,��=� 2�gFtE��E��p��V"���#+I��_:�'~�y}�}b�|�?�Eq���㷓)bD�J�|������?zP�g.���|��
�#@Gyf�/��ݏ}��a=,H��=/�ѿG9��t����"�==Hs��$��o<�g�9,R܅DI}��mG�$K�gl��������ϾB�hΞ���V>񎗙�Sq��̳�140�O|���ـx,�7�H/[�Ë=���W�c��đDܘ-vX��1"H������e�4*�+�ʱa�j�!R�����v��G?Ŀ��m��͢���b-\cp&�������������`��yX�s�������_��ʚ�a��Cyd�]P׺v�;ӇH46')l)S!:��xq�i���]XݵB�a����SZ&���0������Nɇ��I����8�
�_���pK��itwwc���況�D��k�q���t(,f��z������C=x�;��λ����N�y!i�a����q<��+x��#F#�"��d��}濆B�7��^���9F�:F�b�˪�UiR<� ��gc��y�S�c7�����s�|�޺	�ݹ��4
E$�%���VϮXO�!����Q���q��"�Z<1sdU��5퍄#�׶X��������utt�g���5-(+�a�oI~�e����;7YU�=v�z�Ulڶ7߶�^�J<��Jb�aY��^|���(<9��ul4�c�/`��8v�Bɨ »�R+�F�g�{A�Ȑ����ٙ�)��u����b�0��!�Z�'&�L�������5�ڰuG'��؆����y��1'��"�-�/s��d�p1g=��1L����x���8u�����ג��n�42�5̊�bR�}%	S�^���]X��kVbtd��� ┚���(br���ɩ��3,~��+������Mh�CCS5�k��ۀ�c�%|~��a�(%&�G�1LM�124���1�z)}�D$7�.���Mg<��7f0a���}Yŀ�<��ɓ'�j�*��Ԥ[.������C��&ɍ�P�[�ԬL&IJ��Å���w\>�h"�++�W4y�wI�$=%ޓ�D4G8G$C$t��k.�?�%#��"H����/g�2��b�Wŷ��p��i477���U��Z����\A���Z�8�ǃ��伮,sيH'��Du*FC�(e}��Xt�_dY�:�;����C�E�ُ�B؜F:�j&����cjj
�����l?��{�ju3V��!0:�@`
1ʴ�Hjr�g���.�oF����J=)^'<{��$v��
���믣��^�#������,[���\� Ŋ�@��0ř�y�(����em��#��$4ү�-��t��
�fF�F011��FR~S��b�1��U��$�K�S�!4!�I��C��������q)�5��D")��~V+h�L"��}$A,�R_�Z8V���� ,�J=�17��*!<A9&�q�PQ���s_�Y��2򾉗_����Ʈ���G�>q>w�!�Rg����]�1?L^J����zjY^�l����C�/o!r*++��r�	9��is9�2���1�5��09��ߣh���[H�ctY/$����S~{��M���/�����[-���g�$Ā|�m��)�n��1�IY<��U�1lc�c����D���/��Lw���,�ݚn��ņ� �84�A��������Ec��f������;*�!�8��]��pia��XTX��Аx�hEE���P^^N-�c��������<��gY���]���3E�B󥊃tQlF�)>����w�uH$A8���04U��09������`g"��k������!����P8,^˯�M��YM���rCXUĴ
`!d0.����&�]�������[��@)[��=���	V+�zo/��D".^+��Rz*'Օo�^ȌK+늚����kn\VB�_�s���VTh��oFNne�^����+�Sݢyc�O�mEH>��X����S�Yu�Ra�ք�V�ke^������;��$�*sS��!C�@vJ��A=]�[�,_�C��񬊜	��$d�*'��k�N�������	Ɇ=�XBl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl���!�^0����2ERv@�	�C�]0���$�v�I�0������l!{IR$.8��H���t]?�r�Nӏpp9�ֈ�}y
!�O�D9���S�4\N<�4C7Pנ���}Kf��ϓ�/��*���$M���P��Q�`��e닖J�|R�a�x2N�ju��4����"����A�:��|�AI�B�����!����Q������V�;s��յP�(�Ε+����j������:>nmjA�5���w�k�pYrD�F�VA�?A"	k7�*���+{�T�|�C���^>t^��`��4�A%BL��RP�C�'��Vu]���>����~������ "��r�K ���&ʴv�M�"7KяY��-�����/:}+��*7��.+������N��b���Ā1J��:��{'~��Å�:�c%�!�u��E�:��d�Fq~WzIPF�N�g`5�>l����9��`���Z��(�w��l��~�G�f�������/G�W�é�7��B%���vn�]ܝU��,e�UC�G�3�R�C�s��r�
E4�.�\l��ח����(���1&F���|pP,Xq*�QOdT�H��ȝ��lJs+��?���F(�$�ų��>:�
Q8�k.X�T=iˏtU��.Ul>MJo�3 �$��at��&B\"]s��b���z̅!H`2��QR�u���U&��R�2,hT4�Q:���	�L��q"&/4�1X�VK�"�t���j��$/���;����8Q�kB�O�d/�b�a�������qQr�B8��������d2���Q���&�E�dckI��pW=s��1�-4T�p���b����X�Q��D\fX��z�}��Z׎s�/�%�b��}]���8����m�{Rӕ������l%#QY�XV��ׇ��QUU���t��;�$E^$�1� ���1Ƹ����Oy.Qu/(V̂��K����d��H$������.���`:z��B�uъ��o�0c��7�;S�%�Pna%8K����T&��NWM+�#B.v��g.�*�1)�5�B�I�}R��P9ç�Mr�o�@1R�K}〽�DHpOŭ��٫8��0p�d/"�(��L���
b���'+R�j��pg��^�dȱn�R[�a�R�aUU4"I��HZ."�+��0�8
��s�X���^:�������r�[߁DJ06k��O+��ٙ,�d�I�ݚ�s�KIT��XC^G�$^sxՊKED��1	���OR��2c���K�0:2��U͂�l��σ��W���(F���+�]`�ז!A���?�|�̦$%�b�|�t��THSf-��+?5��"B�Z!1@�{�����|��$w����±�1������uU3H�Y�<�h�&TV���w�h�4�R�}��$��U���,�9(y���u�5q��jx9ܒ"�DP$8)"%��d�	�vY{Dc�~ސG
�qL�O�=�X��5�H����T��܏�� Y��z�H76
)&Wѥ�O��2�I���[R����M�d�	Q��^-�Lq{ܯӏM�K����#C��s1x�l?V�n)h)���\����M"=`�MQ&�xb��M��S��82�G�\H˾@ar�;���$��9�DBQ*c���t�])�M5���'�E���EgW��5���4�J��@������V����=A����~�Ck�e!�x"�@��I�z�%��� �s�|��3@���.?"���"O��w�R��$-#���帒 +���EK���kr�80v��o�B�H&�y��GI�Q
��"�*���YLb�d1�+���S�!���&�S��q�z�h�su��r+��n������\ 2@��ŕ!$�OWHQ&�B���A[���$Fa���Y4�1�Ub�8YY0	rIq>��7A��
��Hֲ��)nNc���EO��J|G���W��d%��.�9��;怃=+��|?&)F����1d^���u��W���j�Ĕ�WLLHĮ8;!�Q0�-��rA�,l)L1��� �d~6�Q�vsg%�$qd4Ł���[{N��'QE-P8K�T�l*H��\'��i��1�j̋ ˩�Z���\,�S��a+���E�S�a���x=���|�*���+2�{.2s�('����;��e�1�L�n�����h$�-*�>);�pV�fa�������E�fb8=����,&}���X�z�!"�M~?[g���������� ���V�EH"�&�t�yۊ������t� ���8x1���������o�Bp�u.ddO��#bVJ��C�����5DL%(�N+�Xd,(w��4MOxUV�a*8}	ɮ�"F��:G�s ����3K��qZZ#]�����ර�Jŝk���G��W�5�B�5d���k���hz�D�^C�p ��y�ч�əq{f,b+Z>2��Jk`��"3Jf�/��z7�Q]�(�t�%f�g�&���߁����ZqϽ�����3�K�z*e�]�}�h�R�<1q
�CCc�@y�O�ã�^V�Y�,�ޅ���>c	��	�ZC�5�¯�#����<��$ A6ם^�3bx�um�}r�_�η��!"c��96Y���q��/�re�� etS$�kS��#b�PA��yE��|�T�.Ő�*���l+H�IȌpYە�k��kI��|UN����1����Vo��G��� �;�?�dq��a-s��lXV�c��j�*R�2�� ?}z}n��'��,�e�FY�aX�W�1�,�4���sM��{���Xc�glP�قw����2��Hf�����8B��Zq����Ԗ�����H�5�*�W
�vk�Xh϶�ae�W+m&svY�M�-[�sX�Ik�g��oW��0U��a�Dh�>@��Ǚ=��9�a!�P#�&��HF�G2s�-�3��+d=l2sZ�ِ|f�b��:	gm�ߤ���]�������p֧o8� R�.�?�\$���-ek��%9�dq�d�33�,plI��T�6g���
k��2�,P�@�%WV�7�1�榉�JlG�R�|��w�71B^ ���شE�R�[�X���L�Uks��Y��}Q��9�|��'�n>�����6� ^��#<B��wHn��%1j1v�bR��<V&��gw?1���x!�[��ZҤ�%���I��VY�QAi���)��HY��aqP�y�XZ�e�[z��"�"��D� ї�|V,���}):��T�������:X���d�~dK���d���n�X��8͞�]�F�̚6o�B[{���/�������ѣ�|�}�>&��oއ���O�~�s�:���~�(��L�"�aM��nB�#g~H�d� �ER��r����S�9ը0R"����܄��c'�l[�}k���0�𹯗d�Xp:��'?�O�Hē�-ׯº�8��y���I��'(��+�d�W��7%?�9T��a�������s�{qG�Q`�{6$M�Z�[o��߰A��&�Il7�P2�~�<�J"���o�e=�n�ıW/��ߜF�Qњ\b�q�����ȴ�l"�'�e�F���L�/4r~k�6-bV�l�M7o���֊��I$J�����k���5��ضc5���Ћ�p�D?���WN����2sU7�"�"�;�lrĲ�_�k6�7b��6�s ��/����`�oZKnl��VL�MR��ڋ��Q�bQ�R�(r
ay2��Y�Tx�bǵ[�pͦN9o@ԣ��aaYߓ�����Ĩ�)�Nrg7ܼ"���0Μ������?�r��١��r��-��o����jE]C��3K%ua��L	<쪛-��������.LM������7�D3�7�l%�$�[�K����&K;J�D�w������ky�s3[�nʥ�ei���ń���?���z����� }�
����t���4���qf�G��73�Ҕ���/8��0D2A2B�O���gHz(����Q�}�F���7Ռ�N^֪�r�	n��u7�b-b��r0os΃��)<J�Ff��dp1%�Y�:�┟���#��q�'!_vB,Xg6�z,�bæ,���.?lCH!Vܕ[r5�!�fp�Bl���!�fp�Bl���!�fp�Bl���!�fp�Bl�����g*���{��*m/��z"    IEND�B`�PK
     uK\�d)e�Y  �Y  /   images/ae99f124-1aaf-4a6e-8177-44087bd956ce.png�PNG

   IHDR  �  �   ��o   gAMA  ���a   	pHYs  2�  2�(dZ�  Y{IDATx���	�ŝ6�V�}��3:G:�%��Ë�� �4����۱�.G`X{���}?�טXs8>��&��s� �d��؆�C��I�	I��s�w����]]=�4Gu���{�U=3UL�SY���B If��[
{��b-%��t�D�T,4�HYB�k)�kQ ��IP�P���/_%���2���S��S��՗}�����Z�7��6.�E����hT�5I����&�����~���V�H""H,�֥�t/����tY��B�@���+�Z���')E�Կt�x��B�+b�_���"����g���m�{���*�ԯ�?Z}��P�R(C}����mBj�:��N}]��N��u���k�:QG{�@�@A\*[y�B��U%�Q�\)G�F��r�፴�Ĉ�ڮ��c,B\iiëj�\}Hz��RAV���,�	]�	�~� ��l�x�m�Z�X-��ZU�:*|�jՊ(
O3���.P;�@}y�h�T!��T6�5��F����k�AY�t��)؊kU�eRH�
�֫p�X-=�RD}&�D���k՗��VM)-UW���j5~B��R�
�VD 6� �Y��vSA�.�K)�T�����s��93�4Mj�F��KF�����k�H�C�i��;D��i��i#�C�+}Y�����7�K�UM��W�k]���{�����r��;�S���Z�k��ȿ�,ԧc���_W����|x���u�w�P�$ĮM�n۷�� f�fL�K�RRn��Z�s=хrt���?�Te���2�d�~��Zx�hxL�ϱ���0cBߋC��o�:{�\z�~��Η
�L�r�
��%w����~��vK]��cp���w6�@��r��^ARިB�u��a�"�+�4c)�I��l8�a3A3����U�����p���j����~c�t.�E�(|_OK��y�V�[*���T}@ �AS��ե��Tܨλo Ie�{O'/+U�Zr9tҌ��,YqP���enqfĺ�n%'L���\v�ԉ�ؠ�>��TԿ�R1���·B�W�0EDp��VݶJ��Һ����y�HsPi~:9ҍ�����^0м,tf�-�VRS{5��Q�u�������:��������p���Uk�5M������y@�9)^}���y���ĥ�|V?:T�^����3]8���T�=�֮jh�=Lm]�l5	Z�N<�K��?NO�����A�W5ռr� &	AV�\���Q���{�q�d��gNq&�O�j�����e��\��=��ԠB)��Kg�z&L*�.U/��H�O��D$�tL��0"S��e��)4�^=�����9��k2�۱3>!X��2���8��4w���'(b�:ay�����T%�R��P�R� b@��2��7�oQ!��ɾ�{���Z�2�nԃD0z�i��<���g�{F����7AW�m�?�����H��m� LDp�ߦkt��Ir�d����3�l��U"�	�7�C��{�N���D�۸�4��A���o��.O�a��5)�b\<����z��wI!��#J��$/ݸ��Е�KnI�O4����N�U0uSc�DBI,��
�u���R�֐��� �!��T�
o��A������ �z_Qn�p�Ǖ�n`���^�o,��dp�����?��U���J������!�ƃU�IA�dJ�޵��J�n��D.�eg�В�l�(�6F2 �b��[\@k�£<���h}u���>�7�N��;R��ܕ��$~���G�4DI���� �@މ^z[P�E���D<	0��KK�袥�F�ؙN:��=���[#�[R��W!_�[	A��T ����U�����j�~�����/>����;Z�i��:�vH�_�uy*ߗd��	j��\����"Z6�P�K��j��+�$���'6k˩�:�ZIu��q�%�R�W�@z�h!�T�� � ����_=$$�/��R5Z>/�X�>�L�^.�-�C�:��`�y��2�7�����W�d�W�A�@� ���{��ԗK�k��	+FH��)�>�xi!]�ZI��4��B�U�`��.w�*��l�W�� �!���S�)�*�V��ma�>�ʲ	�N��h�<c9�2)���B,ֈ�?���~A�ɠ�o	��(N��o�K#]��Ě�� �����Qy��f�M|��K}s�
�v��X��0��۫ZH����/�Q�q�+7J�	!׍whqy6y���>q�'��h�c���7�Z#�թI����w�Q�p���-5�Q���<�]���3���w|"u���V.�%]��=� >A{��|Y�ǂ��	lAds��6f��>J�?<^ �on��� �X]���V���D�1�],B�;ɡ���x�p�<^�w����ق �1�	��ѣ*���ڎ��� �e����O��Nc?]��LR,��ޗ�E}����#�%���7}M#M���gA���(�<yƼ? ɆO�x�9�|u�T�+�D�
�_���-:�7�w�A`+"1F�N�?S����.��P_R`���F'a���m�����
Z�N�^wy*_�`�o�@لsu�?	�8�
bm���8�x� ��'f��;�jR����]ݪ>s��j�M0�D���]�R�gBҭc���q���sD
06>Q�@�L�ggIP���y��{�&����Y�Zm�ܛ�BcmS�a|��0*���	�w��R�Q�go��nT��G��O�
�,pz*��G�!�6ic�esq�\?[F�Ow�'GZ���zC��̥ZG���!_�n�� �aN����Y؏�چ�gݲ"JO� ���9�����P�a�:Aܥ>�?��~L0cD3��s�%Rjϒ�+bm���J�.(4fF���'vW�*�y����j�19��#���+B8����!�v��tozP����:#��� �Y ����/n�O�[o$���U���u���BM��U�˄6�j��k���t�dY��) f��]rA�W���p5�����.�w�����P�R�`Z ��I�*�R�R�)�bms��Z���>��r���>=�k�;41��l���@M��SA4��S��X������T���I�OyȬ6QS{��\R�K��t�W� ��BM!K��.�6��ѥˋ �O7^>�>>�L�'�cm����ݠ��{�WБa� ��H٪�o�V�B�e���4]���:�#���D�Y�a��z,�;�9�$i���w�տ#8o�)�s���a��]�t��"#� �����Y��¨�NXN�'4���Ͼ;�z�� �΃�s����Ats�m.SgW+� �>q�nM)8�Nj��F}��tW�I}'�{5HpND�ȵ��w��B��V�y6�+V  ~�$_���@5�Gw�Vu�͒R>Pu�w��U!�4�9py����gD�'T���1���é ��O(o���v�6����G��4z[��}U�L
�h�\�J�ww���p*O� ��O,�r�P~v*�=�k�gT����!�0�-]zSz{F�K��[����d�#�[�i��G�h��.�e�:�Xw;=�9y�=��y�z��� � ��C|IĘ�����R�PN'@2��N8o������蹎T]qkGF�UݱC�5�8�gPP-!�Z�72/��	K�u���޾>���7^hH��CC�+shi�񚚚J�锞�f��dg��aJ�D�'�7�+3z��~ v���Vuȝ�vl�1���R����r���W��r	K�
���jko7^'bP�_����v�����(?7�X��Г2���hAv*�>��N����o������]�D1�ܕUqK(jXl�iy��1�$������=�������g��YYá��)+������")�kE�Co�:es�_�� 
��B�{�]*m�Z���ɵ�[�2Lې8�巙�A�˙`иlWVZj��7>1�Ku���=b��ZA���o�����"A�	?�^��Z�3�^����rqi%�q�p ��Rf��8�"$&�_|��5���3�jBnUuLa�W��Y�0NO���1�u<�����qq���B!jnm����ͥ��2���<�����Ç���Gl�v�iٲe�Η��ڌ�@ @��4z鮨��ʜN��@�;^��׹�0�1��ӥ�ME��P���9�(�Bs�3麵���@ϧxv��ijhj��(U�����Ӽy󨤤$j�U�.+**2�p���t��)��/�A�����Kiq1-�;� >e=�\�ξ:���^ڣNwea�_s޲d� "�J�}�պEe�t��R���]��T��	����***� ��ə���A�˅^H���F ���Q}}}��p`r�
��pp�?|��Ջ]�nMD߃Bܯ� �ڲ�I&ID#�%�Կ��/��k\
�{�q�ܦX�>֬YC�-��߇n�ʕ�r��qڿ?5�h�qp:z�*T����Ȧ�jt��K��.��[���sg2��AT��[ޑ"y����֯Y�O--$�_��F��̙��������i6p��r��!#���%q�Q���s���!ć+VSz�F���E�Su�Ǝ���U����`U�frK� *[u�*]#~Fh���K.($�B\�ƺģ�[��V�^Mv�A�KMM�ݻ�����/1�Q��۴T���jn#q��Bo����@�+��d�.�8����Y��X����7,�;u�`�q"V�삂��k,; �6F�O���R�E�>���ZZQA���g��7F�Su�JU7q]�la�TAė�%dB-!1|�ZB�Bh��F�y�ȍ7at��ɨ��o����2�[<_YZ�k�2]s�����2]�wL�{BV��0ZBb64P(��8��C�]v�ʯ~����G���Z���۸Jћ3^�=
�t��J�Y�'K��	"�g�1ASM!~��%ĵ��6:�;��W^I+V��x������=V&�+�Qa>�eƫ�Qv~XOzT�H\5ң�r��D�A4�PTmn	!��?oSgq��k��ݭ�9}�R�Ǹ��xy9��7`�2ڨꮭ��Q��Ȉ	Q�!�{Bk��8��/Wr�����x�Q�ܵ�{Յ�}�}_��(�� �O\q]��
#�{Fw�:�9�z�XB���q�Chp������n�f�|Υ�^J����Ge��`���1X8oA�⺈뤿�Y�~@�e-!_�㔠6�FF�~�j�U��K <�@cs�3<Nܵ�^K������<^���"c�#�_\'��#�j��v��T�֒��v'd�	Ř�������C�g����F���Ss�>���O���ȁ4�X������0�ў�[�V��-�	7�Q�Ϭʓ�Y��a{��2��a3���E�x\6�7��ݻwG���cR����xǣ����iB۪긖D��5����}Ǖ<���̪���b��h��<�h��}���M�%�� ��U܋�Щ�����T]w}��.J	De�ʕ*�^&��ׄ�r�A!1�=�)���,x_��D���3+1͇�G��ԣ���iǅ��T�w}�_}�@BQ��e�P-!5t���L�'�`��͝;טK(Y��>�>}:����(qp��-�3Q��r]ȗT��Նڗ��>���{�A��m^��{_�!�H::;���?�|�ڵ�lx��A�ǆ�Qn:�$
��ͽ��i�Չ�[��OՁ_�����>��32���sy^V*]��{'�
�/���2J6�ϼ�ǎ�(�c� J\�q]�a��=`^���@�zű�"���9����T���y�!��ZL�S{'+�ws�1�㭉��k�0�
�V����{(N�mM��x�S/w��1tO��1��,FQ����վ�1�c�1�K�XC	q���A_ճ��2�\���^,�0��=�����RSS)Y��1��/"��X!��8C=��F���/g�.���[]�d�V�
�_Y��{X[� JvVA��j��E�x���n��蹷�&_Pu��!߫A�#qD$/A����y���w�r�Y2_����<M+>f�����֮:p2��L�X(U�����H\���}B��n6��e�e���D"���*�^cY��8|,���I��!��y���T���B��ue�W�0ŉ�	��U�ߒD?4�g�9�k!�YuR(�g�0��1��r���^���z��"��	�U���V���@\Q��KT�`���C�d��n�y��s(�d�eu,zD	/'#Ũ��4�����Uw��W����E�K�sBPԓ��Ҽ�J��!��ׁ\�=l�:Bh\w�/.!��}�L���\�dNy*P%��������l�aV���Ab⺐;/=�Q�N��qj���mDe��wJ���K���*�J*C�U�m�6��O?��X���A��:��s�ۣZ�����@m��dS�"Q[��_Z���хՃD��t��O�Yr�:��Ɲ��Z'�Rթ��u�n��Ќ�z"��,�a��d�����1K>\7r�ѡ�II�K��g3ِ-������
�;��]�ƃ��|���u���A��:2��G'�Q���ukȿ�)���pWm��r~^��xn$Yi�h���Ar�2���|��~�����֥�vA$��,Y���|E�F�����<�w�1k]��:&\t�E�2��ڢ:o�E�������7��Q�:�h=و�������
�+��TSs�C�$3���}WW�%���́QR[��2��Z�xt�Yt׵!Տ�&lDNO�z�����o�]�q������Qƭ�9s�3�3\w[{���?�\���s_��w��&��'�����U�jU�&+��u�k�G��ԹW��"�\�M<J�s�EK�4& J��T���	�Y�t(\�r]��V�\��;,3iփ��]�R
�3sy�:xk �̈�u�G����N�� ��G�fV��ץ_4�Pc�i���L�����h�z�B<a5H�%�
	`_f⩯͓�<y�V�XAɌ��+\��p\���'��En�F�hV�ȹ�򟄤��r��<r�l"���EO���Ad�&���u*׭��Y]�V��C5տ��_m���d��\��3�3CyY��nz�A�U��#�]�Jx``�RSS)�[Q�,p�ʗ�ڻ#�������_m<XUO�`ւȑ"UsPD�ZwA!4K|��o��g�KSK�,�dduY.}�2&�׭\���3Ӄ��
��d�2�׬Q�{��Ԟ�e._67��&��g[An.MA�-�d"�֐:F �p�u��ӝ�5�R��o�oc��Y	"��G�ei\��q�`ccDٱcǌ�Deee�L�����xF/���Ƣ�Hrݜ�A��T�C�]����S16�-7'���Ҩ�?�I�}��%]�>���c0�k���UyRG��s�U?7��όQ���YzE���77&����NE��>}���ꨢ����+����:�h}'[z#��GU]��~��n�!3DC}��
���ֵ���*L\IQ567G�=��g�%M�ege�`���}soԳEe\W��Gf���� r���M�?l._2'�ʋ��LN�:�?�Z�x���ʕ+)��>Z�S��L׽\=�qA5Vu����m���=f,���?j�����!8��ߔok�|8�[
s�Υ��a߮�ת5������:��
"i*���c4CS��H�ܕU�D���%��9�A���!� ���w�y�n���lb8]׍}�1�.�po���\v4rPT!ĝ\w��;��w���$�ZC���h�y�'�h�L���`T�_��W(��>��1����wp�.��s=���~L����o�Ky����|�-/�ή.�5=�z��q��ɡK/����l�l�� �|q���/�;���������gO{i�?D��ʋ2iI9�k��Kq8hтt���e�U��͍�AQ<h싙�j	��L	S���g���9�үF��%~�����]�k��
�T����U�
�؉Q�v��e��kq���3Ɣ���u�9�T;b��S����������D��C�{C�J2iN1><0�
��i^y9���<�+r�mv�e�Q<�裏���Y��}�}�J\7s}�12��$n�_�0�D�i�����Rc�PSS�:��9����c;�}x��w-G�f��bc_���� B��Ρ�-�T=d.[�̢2Lx�h�ܹ�70խ�qžs�N#�JJJȎ�jmm�\���>L����>��d�N�� ry�����q����鷴��N�>M-#��9�֭[G�W�&;�	{��5��R�ZBB0��6�������ꙩ�y�D�(��P�+���0����_�9��+z��֬YC˗/��t��!ڿ?utt��f��9�i+��\g��"ʹnW/�"�j�����r7z���;=-��N�������\����giѢE3���sA@M-�Q)))T1>�c�;�a\g��H50�s����T��)"!����-.ϡ�<��`��=��K�P�_D��=�����H<z�|U��LӜ>���Ƭ�<�C�E�p<Z��� f�ً˳�X�)��:��DN����2s�g!ZC0{�"_�ti��F�8xٽ{7����4o޼����N�V��=Vp?���0?*�T-�>���T��)"Aѭ���,*̵wwYH\�s��9F��Q�|��'��<�+�蝟�o��g�e\��3p7�6㕧��ޏYQA�1�Cfz���㺛��As:�Ud� R	y�z��\�|ZC`\��8F �����m�A2�0����r.�b�j��dg��pn"EWq��ZEoM�Ϙ� 2���֐� �ށ-q��T-DH<p�l�@��Kl��pWaF�������DN�k�t��|�|��{��`�����6��թa�p'��?c�A<X>/7*�T��[���m�W�;��?%A$��}ӭ!��N�Ee�� ���r�˸�Ád,�t7��ïvb����ώ�R{�@D�6|������D��6����EV�Ck��C�~��O�А*ׇ��W��4��555����0�+_~K��b!�p��ѡ�I(U��n��5Ծ8��}�A������R4�)�8@�T+&�B��:�[E��CP�d�����;������r|oH� @b�:�è�x[D9g �f9=^����r��  �U���΂����\��y�����I���Θ�� `�q�n5��r�z�� *[y�B�$�4�/�3=ct ���:�D$D%gB�����=�9�t!����f��� @b�:�����ȮܺFw����\��9���]�q喔�! �D�u�gG#�kB��s3De��o�$�F�^R��r  ���zs�ܜ���&���)�tҷ��l/(͢�LtR  Ht\�s��!r8,��2�A�#)���|1:)  $���A�(_W��dGZ�t�������-tf  $������(##&5���H��Q��I  �pݿ������i:���]�D�\m.��(�  I��~s)8+��G'�}&D^i*+�M��k �l���h��(��h�|��gRA$��y� H^�� "�h����5��N���\�, ��8>5?S$h}��ۖ7ռrh"�c�A�У[C%y�T��J  ��88��"�S�ƭ�����p�e9��rpY  �q��h�V��Q٪�VI����D  Ɏ���#-eBegG������?� ҅�*�O��,\� Hv��	m��"��25A���fsz� �(�s�dǸ#r�D�5^�eo9'z� �0΄=�#/�q�9ΐ����X�7��.o4��]��J�Yi  �q&p6�vFN���^����;n����\6��� @$�s�d���r��  ��P{��\|�c� r��^A������9E"  ����1���J*�8KB5U�z��-"���"�q�	A   88#�0M�7�%tnA$HX\��    +�_D���Y��3��/�X�m��!�,  �bd�Δ��w6Z��DC))7����g�b4  ��3����+��g�z���{b��D�L�h �x8+�A4�)�"%j4��B� ��qV8Ս{=�`D�k7�]h./-H'  ���Ȋ9[���h5���L]���2�旙�   ��pVX�'�li#�o���A$������  0N�*2��Be�����ޔC�7  ����:|�3�PZ�'�n���<�vi:*  ��X�'�l��6*�\�*/#!"�ig�9� � ��pfpv���-*[8c����oDRX��p  &���<�g�z;����kx�?  ���5 �p�<^DB���2��  `����*c"��x�m��e�y��<  LN��X�Y�t蕎т� �R�j�;x �&  �����i�|�h$kv��.|�ZT样  ��s�d�u�$��A���4  8�!'B�[Uք1wV�j� � y���P} @]�����E�j�zta���_.YY��uyYefb
HN12$"k"�H���1�pi�M0��'N��:��ԩ	�����ZZ[c��?o-���E���$�da�!F�|�l���}�$Y�r�F@�;r��>�T����M���@����ޣ��|Z<JK�,!�D6��mp��9�"Μ���'��g�Hj�Ek�� �}��g��޽���N3����}��%?/�.]��.��BHT�%m}eÙC�A�2(����Ѿ��hϞ1/���?������O�K.���W@��
�����_��#Zi~s�A�������4���V�p�
���������xe�@������e��Y5*��Á�Ɵ�|6�<�V@���%g3��Ks�*���vF܆�=��|�m�#�x4M��n�������\p�����ͥe˖Y������7ޠ�_�Xt]��}8 _S�r �x��F�;�xg�%�9�_�]��s2����'5>��[o��ݖ-[���ᓑ1u�oq��r�}�Qoo�FUUU�u�֘���|���u����!�xf�%a�3�vݺT�G�ޜ� ����wޡ=�|2�6���7衇R�u���p�UVV����OO>�$����=h�j%�ݵ�@���A*sT��޽�ڒ��e�;ȡa�9�O����oR�ɓ1����ۍ Z�~=��?�V�h m߾�r;���F���)/7� �g	gJw�PD9gO#�=l���7�5�����FKbt������~�е6iepn۶��Q�������?j��Ku�-"�xÙb���"��?L�ģS�OӶ;HJi�����{�숃��ޣ{�������o�ܼ��͝K �3%�j�­7���ڗ�ξ)=� �p�W^{-f=��t����qPz<�s���#�QaA��L͞�fw�3�B��I�� ��*���ΨuK�,����7t�u�Q����0��w�Kǎ�X�����Fi�8a��`�)2<���n#� ����?Q �*��k��/%%%o88?��C��;��wߍX����|Ge%��Lɞ�5z����[t���r~v��F�c��ߝ���>|8b�3��M7�@ v#S*��F/�9͗渫����}��r逻F�0<���È[H�xߋ����S��2S8{���շ�DDUj��g����{z��>�\���_L������[n�Z����jea�=�1�Ζ���!��,P��6�����TS��RpT9wL���)��>�}�{ߋ(�c���_�
�gKD)=*�R���b2���r`o<�)�%d��=�������OG��p�\�AR��8�:{"�8�R�.���� v���\AA=�裔�x���Q�i.%>&�Ev�a������!)K̷�2D`c?�ܲ�WЅ����xy_��D��1�c�b�V ̆���l�%��F�$���ؗU��.��|�AJ��<�ħ�~Q��Aveuۇ3(E�4��-"�'K��bv�d�$g��\i��ǆ�Ƣ;��!eI
��#�Ԭ� vu�ȑ�����ݴi%�g���*x��1B�Yf_�����O����G���������O�Scf�p|��r-&����Π!E�yT�NӜ vp��jmk�*O��ШJ�^r|��X͝3� 줳7:[T�H�4s��4/� �ƪ5�qn�Z���A�cǎ�r>V"�����lQ���ZCQk0�ؑU%skh��U]w��`'�٢2(E���5�O{���U^�8-Ø��2�� ��*[8�,/�!��n�����6n�h�����W>;w�(�c� ;��� ��C ��^����v�caD vb�-c���V�*�+V�:�"��lnIJ3w�Fg��6�n�+W�$fu,����&�l��	��Yl�jޡ��R�aV���̦�������YT������ձ�C��Xe�Hg�N�ks�4vcuv���G0��X�EvcyiNeP
�)��;@BH�$���9+�pH������#--�zz"�noo�����ca���N8[�8��9"n�G�.yc�G:�hLQe�"���l��ė���6�H-��duv���@�/&>fh���Ȗ>������B����S�T�8p�.��r��ca�����X^�S4zi.����E�<x�`�ձ(�8f ��*[�Ks*���ZD-"��J����:"��l���"B��XU�<�gkkkҏ��S>�<e"��l��"B���t<݁yN���j����M��<)�c�) �nt=F�H����6:+�-[��>ڳ'��+aQt���l�Ý��o7����0� ��*��E���$�s��|�D`G���N_��U��D9���s�ݸ��p����)Y���������lQ���5�/����6�����'e������A��n��ؕU�p��j2��" ;Z�tiT�>}�hlڴ��	�3�# ;��!S��?!��E�4o�\*..������<邈�ٌ�# ;���C)R�&�h�h��]u��ʟ�Q�駟�SO=E>� %�W�g3>6 v���-�A)�ե�~����V\p�kk������B�ַ�e<C���Y*��ВE��c`WV��|i�4��< P/ZD`sW�3s�(\Ask!��>�]��؜�9M4���M��2�� vR^VF_x!}��g�O?�4�^������R"��ok�>& vfuۇ3(%ӡ7����!n�jk��?�!��}�{T^^N7�|3%��^{��73�w�!�V�ү2(�d͟Z\n� 	:�,ԍ�fi����4n����w��}�ߠ���ot��S"��O�}��ǀ���q�p�D�4���S�p�
���x��o�r3#/��ͥ��QSs3���"�y�o~�Fq�(����!d5���8 vǙe8{ζ���D�=�"�7�puuuEu^���ύ
|۶mTRRB񨱱�؇ÇG��^r�� �3�B��p�HYGB\9�7�ҭ��B|�%
����.]q���������:�'ܚ�Nǎ�Z�S<�>��L��� é4� l*-5�n��f��
���ΈuG���|�+���ҽ��K�����%�w�}��rrr�}�}���"�ZDR�:����;@ 񤰠�n	#i1%1W�>���{�9���ﾛ~��_[�B�X���B����~ni�.�MhA�q��ش�������Ff�?��F?��O��k�%;y�w��?�1�ڵ�r}vv6��n�Xr�,3e${� ҇D��!�@X�h���o��o�Iu'OF������E��~;=��C�~�z�M�w�'�|��o�s���o��$� �U�p��D�Y'�\}"6�vx��W������c�6bW��p�4�u3�z�޽F ��s�K.����f�7���,����ï×�����'U�D�'X~6n�B��
���ظT/[�l!��K7�teddL�����K���:UUU�֭[�ݞ/ŭ�x �Y��$�I�������pGQ/��W��ћo�M�P(�v�h�f�/_�����њ�g��y�7�W]-��I7^=Ə���Ye��6;Db��5�۵w��b�+�o��?c�}�g565�ܖ���u�� ��\r	������e#A��5|٣~VMM̈́��z�L�,ϪU�(8K�D�cC�C'0o�ډ.ܐX���e�
����8H&&炻cs �U��hbd���	�4G>2�Kh�� Qp��O#��޽���>+�G~^�1VO� ��,��3gė��t�F��p#� �q �r��Q:~�������i���������-\HK�,!�Dg�%�9�_�����'���fA�h�lpHR{� �e��$6��P�J�U(}q�Ԕ|����Ѣ��� ɂ3��$�$�<Pub�ߑ�kKQC�"Xh�DAr���K/����������S-�_�.�G=8�deQN���Q"�A�j��?�Y�<����VդZ��"�d��#5 ��i���3F	��]Li��}"  87�bʚ� �R��a�[Ѕ  ΑU�pք�;"��AY��n��hJq`�9  ���of�5�����C�t�<�#�˥��}�*����   1qvX8�Y^`�L��A�І  ����0�1�E�j4�&��>�$�j�j   1YggL�� R�2�c�j   c��#cL��(X[���]�#�8�^o��vP��  �	����'��	��1okqi��x�u}xY�jb!�  `"Z{��F�%�e���^d��Ҳ�9  0��C"���n	�K��E�   eyHL�Eԣ��C�A��5@=�C���   �X8+�,fe�l���2����h��x?S_F�����` T  C����8[�VX�#��D��^  ���ek��"�����~xٙ�  �UVp���>f9���"�k�5?��
  �pFX��L����AT���F�����rCx9'�  �ĸr�gJ���u���K�0Q/���G   f�f�%c�g� "!�T�����ã��U  pg�e���dcQ�����2��K�hِ.�Ls�-�$  �Q���d TS��X��E4��TwE��&  D�qh��rl� R����"  �p�ݶU����q�Hh�M�#�Z;��{�r�&Ҡ �DǙ��`fd�8�M��������M�և��u��"�   8�H��2�{'Ԥ�$_$"��D�A  �3Ύ��wBA�I}���^�C|c�  �,�����c"�Pj_�uz*?V��K��O�i�"��  �g��j}T�1��O��� �d���! @�;iqYn$3&d�A4��v�N?/kl�֮*���9 �d��Y`6(���~�	Q����-{���`q @���"iw��C��zHWM-�(��� @R��-��h­!6�'R������4w�SKg?�  $��9��I�b�
��Q��˳�]^^�¥" �d�u���ᬘ����=R�*�E���.�hi! @���L
��e96� ��?����A�:�Bg @��:��~39���~�IQC�K�������;Ӊ  H\�I���1��uN�gk�mU?0"�N6tSg� �dbDn �D�u=��f�����)5��<���Ĳ�����]� ����ုjB����s�EJm�2b T�q�  Hl��t��~�s"M���"���{�N5�мL# ������L��.˱s����'\��j�2���N @�:j�I�$Us&���<��R���("��]tIo!eg�� @"���uA�g�ι5��+-B��*��� � ��Щ�� $���$ɓ!_��bw��!����'�����	 �����2��8O�D�L��&#��@7~��  ���\��q���>� �h]���I����"�  �Uk�$=w.#)�MI��į4�� j���.ZT�M  ��.o��-�vޭ!6%A��ڧZEU�U�/�E �7�֐�
��퟊�?e}���DAl���^*/�   �?\�s]n�u�T��)����-���}"qUx��S�" �8�ux4�~�W��T��)}�T��*���nj���\��
 O���:܌����9SD�U�{�*z�<*��D]�)%  �����ê5����9S>�q�HR���껌��%y�  ���ާ�n����Զ�ؔQ���N���h~x�����]�V @<�:�L}�u�T��i�T�Г����2(oek9�* ��Pk���#u���� 
���qy���/����O�� r  ���Q�<�W?3?o��j�$���'C�h饲Bt� �#����6ӧ�5Ħ-�B������+���um"  ��:�LJy��_=�FM��uB����o��x��3M=4��� �	��\G�	���b�DA_�.�*R��&��W׎  ��EO9�T���-M�i��[WI����F������wҒ� ���u2��f:��O�Ϟ� j��x����/]^��h+� �&�N6���6���8�?{ڃ�	����5���g��k���  f��\'��������3DA�N�*zI��6�����r2g��   �NnX����!Uw���0c	 t�qr�A$��J�� ���u��(�㱙�f,�����������g�;-`�" ��œ�ql��鉐��g����kb������-*k�����dyQ ���7�8����cF��~��n���q�*�xB���=|����E/: ���u���D�s]=��ˌ��\n��>���#-���E� ���Ѝ:7���!�s3���Jw5���5�^/��������U�  0����:׌��Y�uf'��;�py*_$w��sSq^i-P  L���F]M��u3͂Y{�ghP<�pЭ$(�ֽ�����,0  ����ul�
j��,�� j<XU�\]�����������x�E  S��V�cͤ&i�W��,��!B5տvz�U����r��v�_�E.�[ 0%��׭f�����b�E�>��&�#R�[��{��-��  �?�S��:�a�e�D��{�#$����7����㭴fE 8\�r�E��;�,�� bA��'\/��6��z�G\Ȥ��t ��kP�u�����%�E1I�aAb���ÃM���9  ��u��s�&lD!_�n���S!�G��M����f�t9z� Lם\��II?��w�M�&�X�_�c���+$���'��Y�A�x� `"N���3����1و���iݫK�c.��@9�)3�A  [O�P�KrB8�#��]��T�u�+B<^>|`��5�  �q]�c1�������S�Ƨ����ĝ��'�]t�d:�\�G  ���v����-�z�lȖAĤ���W� Wx�G���Y�A�yi  _�	\GF��eʽdS�����e���JA/��}p��n��� ��M�n�"4���� ٔm��j�^vy�O�//ol��ki�s 0��n��t���e�1[��t��T�g]x��3�T��J��| Hf��6�N4S���!Ճds�"���{$i�0{�PAN�+�$ �dt��Ǩ�I]�=�"��W��������?��v�����)'#.v `�t�u���w��خ�������տsz�nA���r�+��!n\WF  �dWm���BD?�:��D���v�+�B�����{�.��a<: H\�q�g&�|-䯶̀�WAdCߑ��P�X^�qq��� @"��T�Q癩�Pבg�.�B�W��U��Fo���>�DiZ��Q A�uu���w���)��]�`m�_\����g����?d�/*+�  �Dh�5��纑�P\���u�+�$�����t����QQ.������o�m\�E������Y�SqDL�{��Atkxy߀N��oPa�lt��8��;�ZBF�f�r�Ր�)��}-��۳�##���������8�T�F  �h`H7�2��,��u`̋uq"��ȑ��JWm�,��?��u�m}�)�@7\�" �x�ø.3�$k�����@�sqD����@��r��m"Q��LS�[�@׬Ƅz _��:��h�^�tg�־#jOFB�����S���U�(����@��ht��b �l2�.3���qg��J	DL����R-#��yݡS����EK	 ��>=�B���\'$m���HB��w��7mф�ռn��6JSa�^��# ���'ڍ�ʊ.Ŗ�NJ0	D����E���M�����|�Bi)Z67�  ��șNUG5�Z�@�����2�X�W���SY(H<f^�#��e: v�C��cJ]ꏫ�g(A%l�������u
 �b��{��Ϩz�XB��]�eD$�����5F�
 fɘC��|1�~�\������x����r.c�����r� �8!��t�R%;C��-��"�X^oϝ���U������ ]�։�t 0c��q�%�[�b�~^o��>t�D%M�0%+�����j�
_�-�79��8с �wL�{BV���"!��	"�x���l�m�����<�A�U��\��]�`�>�i�ܵ&���:�J=%��
"�}�V��Wu��e���P'��< �J�mƳ�V�%�!�u%��"���KVx��H�/��1~��`����a{b������r\���F%e1�L�t�M׷gd�l�M���O���X��R��|p����
���	�tO�,i�����������9#ƃ��B �O�`5��0�"w�N��q�$u���\/_��zp����W�ukK1�+ L�1��cN��Vuσ�Q<��S�b56�!��7H׭)��2 [W�1���̪L�|�� #0�V326���F��?��0�( KsG?��B��{ �&��&a0="��Խ��j>#���( ��h	|9ߊ.�-<MA�c>#we���y�q��  V�-A��̪�nI�I��(��^�^���c�°~e1]0/�  �}~��vh��V�K�3Ѧ��J�14�?�2w�����2r���^k� ]���  9}t���l�\�ZB~�h	m;@�h���U��*����?7���`kg�1F]N&'@����]�F�o�{RO��})@0&ԜР���.����<>ݭ������G�t����d $�S�=F��Y��D����lN��&A4A#P��ܕϑw����۟iݲB�T� $&_]�=�{)����I��&A4IA���x��K�� ���]��D�@��NJ��6��3�cmv��#�%��9���u����F�UYSa^��m�t��b*��ï 񮩽����=�H	'�.������!����9=�^!��!��������3F���0�@��I�3.)�k$�T�$8'���x�8=�'T��V��p���._QD�i����}?<�L'�]1��D?��&8/�)�U=\���/ս@$����?�PK�
�bZ��h vw"�Mh��+NE�.tR�����7�	�?�2�m~]:��֙��4��jA]�`l��C�T�U&%�Մ~O���=SA4�>�����Y�m��<�:�:*�O' ����>��`��1aO��U�Ch�!���mT������$�e^��� �EKh͢�ٵ�x+}z�5���Bҽ�ڪ�	��h�j�^.]��=M�R���m�����dY!�0�����Ҟ�-1'�c���R��׀�z��h�����t{�~a� ^� ��<Z���� ~8u��f�hg;�!�����h��UO�y�xOʡgU�\a� �u��BZP��u ��dC7���e�T9�>B�/�G���� �!�6��^�ZG��Z=?�چ?�,D������T� `j��
:|z�!z���Ӑ���3A4�T���NO嫂�d1��
��.^Zh� ��L}r��zc>dxO�|X��n�� �!��~�˽�a�Ϭ���.`����..��"tf �,��e߱V�S��Hп�	�Y� �E��_�|U���h��� ��7@K��Ѕ*�0���:{�3@㌔m��I�H��3��"�j��g�U/�:WW�����H��E��:���K
� X�о��2�Ij��|$TS�k�Y� �	�@����H�?#wYm��ώ��q -)��#�Q|��C���&_�4���	lAd#������Խ��i����z�������'��"OE�)��䐼�4������{��P�n�����7lAdC��Ay�驼G=�ZHeV����y%��ȧ2�� I$��K��6:��3��!�s�� �������u���>�)�'�A�e�3����Y��T!q�Z����N����V=�Hx�~���7�Y� ����#��wl�����9ֶ����ZHyT��@������کn���FI)_��Ёm~�Cŉ����]�ʍ��cVs��*/��sȳ0�
s� ^�t��O����O$�h� �X�_�� n ��Lp����}�]���ձ�=V�i,<+��yyx(�
?�z�T;�Nચ������_$�;�85�{����]�BzH�"ֶ�A慧�X>/��e�]t� �42.��~�N�^ �[�8����z��p;��zI�m��~���Mü0�t]�sP-�]4G%�'�.1 ���S/Ϲ<��%�C*^��ڶM}�?:�l�2H��S����;h/���۫��/����A_�3	�O���>�\������DbY�m��_s��X���g��$L7~܀G�H�a��W���_$Q��������� #��k�ўv�Y���<�>��T�Hy���]��=��o�|_�
 _��	j��U���*�n0ZHBx�ڞ+ώ�)v�j%-tb�X8w'B�ƀ�<3�IYe��|�o$<Q�P���J�޵�t�x�ኃ�ĭ���l*��3I0���~�t��4aR>��P��zA�@%���)Y�}��{���$���H�o3���4�����M٩0��k�N��PsG���'I��~74$~�x#b'#Q���Q^��WHy�x��W0�|z��B�Ƿ�f�Jɨ�{�xF����!x&E�j)�֐��� �!��/�qEPU�����Fw	�o���(�xx��H����������i����9�i��1X��+I4."��E#��d/�� 1�7���^��ƿa�,�&NL�K0*F�2�I�d��ʐ���sn�"����I����y M9��<���8S�����O!�Ie�)>����c�����(
�)�HLJ`�.��=pł����r�$�����1�j$9;Wǉ('"���V]����RW�m�З̍Dlhe*Dʮ$b�0Fں��!�!��vo�r�*�ə%���T�Z}�w2�Gn�Ysm���]B�|�fj�(��)O� �;Im/]}�  `�^�cw"��Ԋ3�lC![�"~m�5P�@9~V�yH-��bs"<�����8��ǐLݻ�(J	�)%��O��2�|�<����z	pbS�K�/�$�KR̯��VW���M�'�Ys���p��~B�ڡtl�>(�>Q!R�"u�����.�F�J��R��0=x�����!m
��x:�T	�<Az�0��\,�k�Ug>,@#������$(J�)�("������zY:.s� ;�s-	���	2���t��C�׹�ݑ��7G�u��_Z)?��F��g�3�; ���o�@Q"�@I�\���7h���D�9[bQ�7˹�R�}��8I���D)�V�55��6����Nyi�w�}ۖ�r�d�,���$�9@�r�3
�w�ѡ@Q	"�P����ϼ�Nk>�E���N�R�u%���菉�s��6��ɱj*���|Al�����˱C�W�q����ˍ����yP�#@�H92��v�78��{�u{������K�Xq
	�b2���������Z�C���������-㛇������&�a�\�7�[��űT&����چ���<��f-��6r�_��R�=_�,u�il��x淯AQ�"�ؐ���
�8�u�uB&0=�_����J����)���/ v	ǒ��~E�T���b� �>�~�B���� A7E )�w��@��U>�(�Q�vbD6jsM�~�R��)U�@�|�D��#cY��8��w���؉ O�I��@ �@�1��)��5�9ݿM9��)'_<���:p�b�u��N�Q'X�D����ū�?�9����El؏�e�`��1>_?���Y��(�@u�C*�~� =��M������[By6�P-��D�,Xa$s�o%[8���8˪�%�����5	p��K�u>?+>_/���c�����iB�g�I���y�˦�<���}� �����Oy��E�    IEND�B`�PK
     uK\hyXe  e  /   images/f7e3f572-2cc7-414e-8b58-58f37a09912a.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs  2�  2�(dZ�  IDATx��kpUU���y�܄G�0!��	
��Q���֖��iUmiO���m��~p>�*[K�X]�Xe�tO�8U~�}�ZSPڥUJ)�-�@B��yAB�!��sά߾�����ܛ��U��s�=g���k��^W�@���'E�\�5�y2�"��(�4�G��빖%5�e�鑥�e���)� �z|��A �z��|���K�oѿV׵����D�����L�L
 5֊8"�4�B�G#��~D���R?Y�X֒���PR�L�Z���bW���Ru�pGuh����ةF<?�z��'�鱤W7��f )���y2�N%~k<�o��?�ӶXV�׉�	ίn�1��m��}�;9�MN���������/��_� �ѧ��h�n*���,�JUY�̘�)
DԵŶ�! �`���<���cI_N&�w�J,��\x�7v��o�X�߫ m֦ߵ�#IӁ�k�U����]�-��� Rռ� `t��T[�47���ԗ��Dݥ����)RSQ,�S#ѧe��^�9�Z���RY�k�I���?i�\��yzQWo��b��ӏ�P��Կ��\z��+CZV�^����h�H�zSzËU�F��Y��j�ʜ��R:%�=��s�Io��N�݊�bZ�T$f�J����_���鉾�����{
_՞���ҮB�ߖ�=oK�$k�T���� =�(�,��1}R�S5��I�pEe�D\kߓ�J�o�@,�W.��)�c'������'�I����Y_ԇe��̽uf��L8 ���j�Z�����WΚ]4�L�ˋ��c�{�x%���s��)�qr�h��{w��K{�oG^Я۸���}�X`&������Hem�N/��	5su�\1��@elA~�p�pY��U�߱����kϿ���C�gN�ճS�pu�Z��5q�؄ b�'1���?i�h�Q��V�u���O׶.�(O���[�R��b�ˑS5���|-�M��a�a��F�1ԁ�o�1�:#V�_~���yWL����R��Y��µ��)�z��-ݷh�ߪ��Q{_W3hz>�����%R��a���v����_�u�������|�a�'A��ߢe�e��UK�eOk_ŗ_����X�˱U��tҹ{�=e܀��w�R���:�[��y����Y��V� <u�<�4G?s��?��D�����,&�[vu=p�/�е��36�R��qb�)K��g�K��s���͒)Q'���6�J_�N���� QR����
�Q^n ��k�Ǫ�ܾ�V>�ٵ�Pg��:oY�W�Ƕ�q_cĀq%Hx(�:�����ҺV�ᶳj+�'{{�Б#�D"��� �g˞={��,��Ç���U���˜�z)/+�Zo�^K�Y��J>�}�I��l+X����R��1�0ezF
�[T�o5_YZqÂJ�d���N9��&.�ŋ�ԩS�u��As��W_-s�Ε��~ٱc��޽[�kk���*{C��3�͛͔"׮�}��CU���>�����X�*�cel�o&{�ƒ��+�SO*�5eK �xw�㦛n���F��d2���ԏ��RRR"+V����J���O�u]�9cF�@��˯�$W�}�ɷ��[�#�6VC?*@R6#�S��0�|eYN���b����-[&MMM�H$F<��Ǳ�m�6������(k�X"B'	ϯ�u��]���M13�Q_�I_��?�pl�� U3�	onn6�`�±���~���7Yu��Jb�'���#}������e]^l�xQ@RAs��3pm�0�g. ��R{Ԑ߰|�z������n�:�'ٔp�BG�q�I���j[n���b0" �w
gJ��>���n��L�­E������)�'���,�:����?��O��i:tY�v�GG�j�ɕ�{c/���3�����w`�M��Ϙ�3�c���0ʍ����ZZZ�Gu�2Qx��G�/���<�Mz΢-�9x�x`�:�`[�qe�N���  �
�BbS�C�f�9�)\�s��PN�:e�߷o߰��X���\t��>���Kz��b�u�s����8,2�6XO���T����oK4�3��o7�lf  z�G}dޯZ�*�2z =O���6m�wd
:CwǺ*��f}�1�������y����J]��`!t��gW�@����u����g*�יF����58�6hkRDu�;O�n�j���6p�������{k���Z�X� �>C
.RC=U�ׯ�6�w�p�3�si��r�C��]~���3z�+(m��\9�M���a<�J�K�$/��VW��ȱcǤ��n�� ��ѣr@ϝ?w�L��Ct��Vͱ�[��#ι�,@����$$�β�d���DO�6�Do?��Y�z���닁'O�4�p.mLF��_F�贫7v���c�s� U鬽T�N�		����J�^S��zɦM���o6=�\����3 ���\	&�>�%:�=kJt_�7����OΙ�b�&�&o�T�C.��V̊�*�a�U�y�f�{�Ur���RUU5tܠN�:;;�/j3��oz`ؓ�]]H�)�=r���j����qirm3�`�-x��)Ru�<Z7�A��+հWVT�����c��ŒP
9��&1e�p�c���hp>����n�*K����?h��: r�S=�I�q�cl ��$6k��ܑ$RQt���ʞ�9FhO��AT7uh��@Z�-:>�5p�z`�;i�?#ז�N2
}??o	��(?#�:��"t��+K��;z�T@~姟~�����L�-���Q8�i $��k��_U3U'����L��d���U��-#���,-�$C��ꩲ�@�ҁXr���[��gv.�A��-$���w9
:F���`G�^�,\�:�"l�!��l	�q�wU�5:o�<}�b�u.������%���U�]�stKxM�X;C/k%��عT�r'f�R����n�}�;Ù�
�"�Fv9xW�&A�辭{p��}�e�1�]�`Y��t���o	X��g�1�]/'<X)�|�E)bVa>/+����stQbq�@�����2�"a���#GdoK�mk3K�+���456J}]�P�C>����`0�5�TH`S>����N
�>���j����?��I�A>,[�l�w�_*���{�V����0ZA��zNI3F}�<�rF�p�Ν����;�z�d%'�v��{N��7���n�ŋMJ��h݃��<��!����e�c�=:<mR0^~�ey��G<�6n�(�o�Qy��\��X����� ,(�P;$_%��?�6ɳ�>{Q02�c�����_�Rjkj�t���e�_��X�TՉ�N�� �|�VY�d�<��c>�s�{�=����?/1v$b��2�MK����Ln�zP-_-�m�p��ŋ���C������|sV�$\�P�,\�MQ�(�����)����r�-�n�si���44�+`�i�����Mx����5kָ��\ڠ-+O��4���(W�3 	*�I
c}ii�twwKWW���׏�Υ�
��{I�.5
)�'y(xD�UU2����?���o\�p.mTgq7b��'����钇��L|�q�|y�W��{���Υ����a<i6�\�w�^]��:�D�X�\~�����?/O>����۷��?�y��tKzD�{]J�R�S�TP"��a�jy�駍�l}����5?��i#���,ŀ	b;���R�7�hI,�L�GyD>��Q�z�MY}�my�B�=�^�>���y^�
�.Y�Hf͜i���_�	��\����_|a����sOއ�t*�����0um)���=�$���?�#G������o�[�Z��-P�;�~$|S�,�b�P�"�Ե���)a�c��I��p�/��Ш�M�m� �V�oS�"×���e�|�g�s�έ�^� U�޵��N�m*>$���g���"�"�e}N-t�o��t�[+�\u����� K �驅N��B�bn�4��o�����\�_}�� 
�S��l�!�Zu�����Ď����a	�0}Ar#��sF�ͮc't���z�X
{D�/W�Zu����X������cY_��q������V����PG��s�d�,�Q�3�I/)o�o�_zmC�a	(����l"���~t�F�ꃤ�,�P/�,�	�����$�2���P]�D���w�y�'�k	��e 3�?� �F$�1k翏�V�vjo����������*�2���ݪ�K&V�.��U��u�����S�$HO��\��f�L
2��㭺e�1�X;���j4x[W+x��e��"з@�G���6�^�a~@GF�ҳ��2�oaKv¹��2!�QA�/�>���TЭ�X;)Xgk�,@�lfl�).)/����2�͠�&�c��C}؏v}�B�;��9?sѷ5ld`����2~a������'Du�����7������y�P%�p�'�dCP�X�4?��s�:�S�v�Y�g����s~1�as{;���z {,8���)]c���`��{Ԩ?\=;��/7~�dk3sR�62�apy��u�R�:zb��c�zT��+,�~�  ���LU*���a#� �%h~
����p��i���|Ͳ���*�텉(G܎й�=C�hx��Q�� ��s	��/�ߤ���+Q�m)�؏���+�E��if[x�����,8���(gK�#�:��^tf8%�ˋ�E13x�uY�Wڠ����ȵ�_;��L��XV*�j�W'�i=jh�`��KUR�DP!,�R0Ӳ�j�݇�>�8��*�r�m���>�ۣ#��)I�"�%���6�4��iJ��6��`#KxA|T���+��~u\���ѷw(8�Ȥ�}oL��c�c�
�((lMLxC��`��?D,�]��0���)�3+�H�H���ư>���3=j8�� �
�W�+�<M\[�)86�S�+9�^E�Mi^��^f�62��"'�3p&}�3pm�B~nɉ3qLz�/��`#� +���������C��3�c�1�ڎ��'��OC?�sA���� ��s)���r�eB'jK����f�����F�ڎ$�\8 5|��p+���X��F�K���,��y=��[����Љ�(cS��K��J!Iu�ZQ?PZ���m��up.A��d&<I�0&<�����J�K�gt��������ҩ�E&��qc��u�l��l� �%h~`�����4C�e\���ӑBBk�,������w� �^�X��G#^�$�@����f9��K���,�	�P6�@��d�_�O�ɓQHyS��BB���;S�q$k�t�c���1�\~�w7�qd'�K���,�	��c��@������~��grmI�$��$6�H�1NKz#�l�<�{p"%�ՀB�D�1I���K���,�	�;��.�%��U��(�M�gç(2!4�a��J�f��e��@:��&�ֶތ�v�Y$C�4uL��4��<��0fاŸ���f_~��P��Z�fu�����-�T3�tF���Ul=f�+,���62v.�Y��l	 =$V	B�!�켩lKN�e��X�oh�$��ުo�z��d,4Q��Z�ߦ�3E��kK)U�wR0�:��&�[X�:q <S��
	l�g8[����K=�s������Y&-��5 fۿy1)2)��%����ĉ:����W��N�m*>SdX?�G)U�wR0������#��8���\�B�
�|�����cv���������+�4�����|T�7    IEND�B`�PK
     uK\P��ޮ  ޮ  /   images/98bdfb38-4044-46ed-976e-d2b53bff2879.png�PNG

   IHDR   �   �   ��ۭ  �iCCPICC Profile  x���=H�@�_S��;Hq�P��"��
E�j�VL.��&I����Zp�c���⬫�� ~��N�.R���B�P���~����{�2Ӭ��鶙J��LvU�A�!�Q�YƜ$%�q|���׻(���F�����c�0m��M��ObEY%>'�0�ď\W<~�\pY��!3��'��6VژM�x�8�j:��U�[��r�5��_��+�\�9��	"TQB6���XH�~��?��%r)�*��ch�]?�����OMzI�8���8c@`h����q'����[�J��$���"G��6pq�Ҕ=�r~2dSv%?M!���蛲��-л����������7��!0^�����i���3��~ �r���_   	pHYs  �  ��+  �IDATx���w�$�u7Z�:�LO��Kr��DI��HY֣$�ِ���'?���1l�l˰`6 �%�Y�-�P��@Qf�$7�l��I=ӹ���s�n��.��@�z��n�p�9����Ҵ���ݵ�0�C?�4mmmmaa��W_�?u���˶�Z�Up� 
�$ҲK7]�������i�뚮'hP�b˰�>C��4��>ıfF�]��8Ɨ�m�tMS���?��MQ�'a�l����8��]��d�+ު}�	���&_�Ou3�EQ̗j<?�|���+��$�4z����H�O�������B���������z�T���|�N�<�5B�F�x@7��^]]}�@+G�=�|������|x��9�w�&�R篌��'N�0�0V�Z�4x�Q�ݠ�+�y���7ѐ\B�Z�̪)y]�eu��������Aޫ:&k �T��٥���!���\9W���K#�7�2�]Z��:u�2�h�$����~
�˲�E�����ŋ�������-[�x�������0
-�����./��J�y���{��ja0��H��0t�{�>����f��W����A�4��Pr�QLF)�	Ͳ���4_WR�[��X���JU�+	��+�$�M�T��{B)[�x�w���S���G��ƫ�~�l{CS��-���6JD��JqY����Ws0�X�GƒDq��GXZZ�������ln��-G�D��?/�B@Y/�|襗^:r��� �kxx���=��hpg���26�=�$&a0�_�x�>�#��ҾŨ��)F�m?��DRf��3hSz�ƶIe��KW�K�ks<��7�M��O>�)@]f֫Ͳr�~��
IF��I�mb�,ǖM�E���b�����s�$���� �,..~�;�y�����;@I 	���i���o��<�t�r���}�b$���8J���u:$W��>C^뚙�� ��Iٔ>��̋�5����U)&����=��⩹r+ަm�<ʹ����8&{{�:��J�~}�o����Q�Q�Dٜ�s�<C#A�B�A���힚[#�	Ki��c�O*���X����/}�w~�w����"��{h�ĉO��Y���BX�t:�݆ɭ6�zc�E0�P�[6�^�B,�s��� }�3�1\U�l�����n�V� ���TR`�
#��/�+�P�u�V`%�5�|�TS�n2\��¢j�F>(,���Y�����mX��6a[]��b�3���g|0�L��j6�[�n�_@�s���|��_~��<�_���M��o���.`>$�R���-<X���� ���Ń����"elG�BJך�S�U�W�W-Տ�k-��x#Y��ڴ�j6��Z�����M�C�t;m�� =�3�*��Mr*����(�O}%�a����q�7�}���,�cۦ�ga��gʥ�5͐/l$!�	���&�ɴ!��,h��9s+�垜�l4Є �w��|�B�4�=���N�P�Ֆ����A�,�P(�-4~��j�ۅzjn-�Qyd'D#φ��tFTBj��r��Y��i���j�>fl���7-X&�,mcgҕK�w9Ҿg�+�PR8�)���.�mi�[J%�mY#�me�<�3=9���H% �-�*��Z�u@�)F^�e|����%��
������WЃkc�1
���y�'|�AhO ����|�˲�d�n�{��aXZhP����e��V�tR>��A��)��<߰��BB�o�^,��؎@"�X"ZK2a�a�1D��&&�.W��޻�I8���0Y��8AӸ��6��u�O|@��툖H:\��Ke�Dxu�-�6ނ��{-($��AڔIĻ��-��������-����#��|}�w5B3ưT�n/[o�m�����"_�H۰!{�I�A�'mbM���f���õ��ݻv��LM����%�/�H�~�{��ɥ�p���Z?�Q�i4Q�}�Wp\�Ƚ^�����?O�3z#��E�D���,����㯌�f7d��R*�Q(s�)��Z�P���]����2u��(���r�
u#��ٚ�X`�����@�)�;A��$����\ӂΣ��X�4]�hYd���j���l�c��[P���Es����3	�R�H�2�8�c9a�����B��/t<�uBo5�Sy��7�A�,yŰ�|�711��(JX&�w���,D�Tb���H0X���ܵ����ڽ�v��#��KV8���"���f\�*ځ�Y_oᩅ���t/CKB7�Xx��e�+���讻�����&��o��d1r�����.�D����ւ�&�e��v �J|E�NȖ���`:�Ne�@�=�N� �$�C N7l�d/�f��J.q���G��p �,��b\#j.�,��=%z�1׶��6:�i
�Y�'im��6-��{>���=j� H���]Ƣ>&�ui?x��	��l�,����{-g�Dg�������`t�ecPE�ŜA(��V��A�X,@�T+%�?==y���Pjvn�:77v�X[�2'�q�a\$\�B���2��ƶ������:��\v���XJP6���/~�d���Įg�@5�����Sn϶�ʘ� @]̅L^L��u{�N�Z�̸q R��Y�Нd#�#-�i7�G���#l��"G0ZP6dm�Pĝ���n���V�l��ʀu%��0�`��Le�0:�0�*a�õ!4��=�e�c�8�u 	b�v�"��@^�ȏb±&�5�����zER,&)���/�I*zF�{���iK���:�%���w,�g�A�EN#�s�Q4�O�ݻ��޵�=SSS�~����A�C�U�׋�&�`f�Ifr||\�V�r�`l""�J�����^{�����U�.ʘ-��C�P����OH��o�[��a��'?�	�^���سw/�<}�4f����s 	���C.O(�2� �Ļ_d�ZN<Rb���y���_O?�4Z�4�;�@ox��;����9��$F��U��,�2kvv��;���`�@��ج�<��-�$� T��
, �wwH���z��S�!����I4�}733�.�e�m�@#DzA@�Qpy8}�LP���0qH��~����i�/�%��&��XD�k�^�^��Xn�u���0��ӧ�=�?33jsH����Q
���U�b0��i,%h��@�{��ű�	�q1!��Ep��a&�.�d�ln�D2���B?f���|�������}�����!��uｯ}�*(.���G�H��<�f��1�;f��,��k瀍�d�@���~���
���aO`lx�u�]a��B�N�0~݈H��B�  S���bˋK�`��":E�vz]˱�����Jz)��`4cC��u��2���b<����g?�կ~�?��Hda-�G��q�P��������!��1p�=$��`��<�}�}���+�K�೥B�[f�����������+���13 ��o�`�X/L 1Z/ȏŭV�0v��I����k`\�S��?�:��>�	�I��رc���
ָ^��c���?���}�B'�YY�-[�@�#D^��m��Tߵcg������}d�.;5��%V7cx�w��#�wm=��^i4�{�!��v���Tj5��l��9���K���g��7�A ���R��@�,x�^�till�`�x/��$ٵk�'&gۼꉠK,3�0�A#��v������ɡ���l4����3�?�37�q������bЦ0'4��{ ^~��e��� ���n�E��KX�V�a�V��bA�5ym� ڸ��c6����[n�EP��/�|�Ңpz���u���I�L�٤ó���dA2k�a��r�
=h����<�Fv������?����Ҵ�Xa����=�����OR�ml�;����ï����.0�n�v�8t�:�^�p�u�5�)�v����������?
6����g�}�g*Ւ�Z�����;b�D�������|DV}~~����RW��p0��e�1�y�[����'N�8u�4z��7�x#��֭[o��&����R��c�v��b����ϝ[���?�~����)l ���� Ow�܉F��x#��<��s"�I+���a7�)l�V��U|짏B���r�R�(f7� �b�P�����{�G�A���|�KH+�Ke/
�b+"0Xi��{X��q����8���aN0���/>���2s�O˄��� gcRq�w�gV|ң2�"g��5�>������	�v��յ�����ޝ��ܽ�ܹs�NoǮ=x�����ךm�u��O�_���O��o���G>
Qr��љ�Y�P��/�V�j�1�����j���?����b����V�xj|�w?��~��Y]Zݱu�?1:����ܱ���3X�������������FC���������"�/��S�J���۾� h����tt��F?-�XYY2�����'��;v��D�.\��?�S������W_��������S����O>��g�윻����@�x��7�n�� ������� |�ŗn���m�[t >��2Q��H�X}�;n۵s;n�`n�CF5K0>V̱�(�M,p�fw} 4�c"����K�j��C��n����K�1'l�%����4m��]}�ssv&N<���#��a���-�}C�TV��'�[���?���=fz@:XH������>2��:{f�XB`��o�����Zh����ܨ�������[n�p�<vg��C�z}| c�͵`E��r�c]����#X!�� (��h�N��a�� � ��|p��]�"�3뇏�����&;�"��g�o�� p@P~���;x����;�� ��o�>�+<����7��q��������mG�N� Ξ=�ņ(衇�F�o09dJ�7���U+����_�}O��J�g�2=h�h0��2�2�!�!A�$E��X��/�����Z��-�T�4�+~c�E5%Ks���`l`�Mv<���?�\��e1	gCo�& �)��-( w��r`�����2V�:�-�]qo���Z�vk�/9���_LU�?Qg�	�������6��A�hV��({{�����i�6�(Dk?��#P	N��#��2"l	�� +`������3�:l���GXx�HHX=� ��?���W�ς��,���Ѷ�}49�%�K�)��#��ĺ
�Q+�_ba7y؊)����K/��Dt4^h�[T��J�\bT���0��� ���	���1/�V�I�u�D�m�G?�>L����`�./�����YHe�R��\[�. ����?��36jc�����D�#�|m۶m�Z���iE�����1c�..�y�y��~�+<"ʩ'�����n���x�hs�?^��|��WŠ���ORt�MܹX0 �F�~E�����~`��HZ-�vK� l���ȴTV4�Aa�p3D!6�{�2�����@�3���ր�03�^��t�6�Z���d�	H@�X���
>�(��%Oሾ�v��U;�4��;�s.��If�1���v���Ξ;w�ȑ�?�8Z��e�)|�BbO`fo��V |�m��n�W`%�}�9��?�  �Ń�I�J,6V�6�{1'bO�Y�"(�wb-�!0��|�)��_��XB�����:v<��x���F����b=�#���n`$Ҏ'�n'1t���6������vƘh<�� �E'�.�/�-�>��A�(��8u��$�K��|'H��b"RL2��ZcD)�T��œ���	�K(3/�8"Oci��f�=��W)� (�	\� ��oN{kWj�5K��b/b�1|/[
���|�� ����o�)� �O���`?ظ@����y�u��)�;�x������ ��{�$/�0t7�\���>��o����{/ǝ�Ї����O��ghP
������X�h|�dy0_���=��o�q�����_~�������Eˮe��T3��b5`�����Єef�' A����n��z���"�A���S�Is�����oAáWx=�"�.����SO��JD�}�V���X�p���Ahg��522�|��LJ+3��6�:	Z�2a�y�-�s��y�Q &��!F*��cؘq=�'RϘcㆯ��_�򗉡E����ÿ�ۿ�X����ȘE���5|
��bn���iE�dB`�����M�x�X�����/|����;�@�>�������Ho�OP-VT������^��c��A����c���6�\7T�^��_�5������O_���p(���������`�29���g?�Yq���@���7��F'�_�8�d�FW��é�ɋ�%�_�[xdJ�C�!���Y��q~A7��&����ǚ�	8,�z���	Ճ$���7ؠJ<	T��~Z���)0�dg��5s�3����כ�J�-@�4[Xo���z3T�ǟ�4ph� ��@�\K^$ F�
�:�.�hH�^����n���8��� ���H�@����ꊀn�E��$G�j��I�@ �W�c�!�@�`  +h���{62YPL��b���,�*��z�� �����O͘2���������� o���G�e��}h�#��4�'���4rr��1#�4��Az�#ȗ�k"z��!6Cl16�hd�N��4wC\��p��=�QIYP�i@*�Hx�$���!����}̲͔H���zF#�!![(��=��"��E��˗�ϗ_����K��P�Y^]Y�hqY��HY��[��{�@e�C@��R�a9\,�h�r�X�q��l����S$�A�E�*/�|�����6�8؃�Ǻ�wI�¢@�&-�\�>O��Jx� F(<@��XfB��Y	��ɘ&�V��O���)��nuu�#w�e;���$8�'��&�M�l�P�H&��b$�@��dv��UE�=r�KX�P�*�ݭ"�T���/�/	�@�$�:���uO�Rd�ZqȔ�M< ۔&�u0����Pe!���;2�$+I��$�p�$K�P	#K<S<2�\�ys��t�+ W���OHԕH4A���z\����߸-Hf�˘@W��/M�f
3�r�<3���1�	B[h�îV�lS`�I�m<�Y��#Ӊt6��	�:fA�j��$�*�Hn4о�qB�_i���-v��ƋN�I�H,���s�)����"^�z��s��P\��Vy��A��1p����	$�<��RȒ��!C-g�P�S��z�nT�WLGBy��t)�S�B^XT2��~j��b�n��c
 �Jp�Гl�:sAܚ%
���s�J��R�A�D� q��+��Ʈ]�`B(���UۄkA�a�i��[���I�=�`:�N��������ů	���">̖�_|J2x���H �_������^�D���MI�<)�5:���av*щ��J�	=I���T��QLaB��S�'�S#jm�e���i�A��ī�"fI�b�~l��E.,@	��8<Gl6��*֘sT��
���3��0��i���yu��i��A��[�� D�%gdQ��WKd�ʞ�5>���[bj��I٬`6
]J`(���vD1�����wEF�?��=i�V��3ǤDr6)�����D��w��V�I� $?!��IjnM��1�81rY�
�����c�cJ�����;���}�1��r�ld3)?΀��g�k�F�EX�l�y�d��<����2ߊ`:[.�9oE�S�jS�HJx��(H��=�8L��{訂1% J��4ܴ<ZF��훿g h�)��E��2;�W�G~��OWsd��z��(����t�`�3�-#Y��M�+�q�?���N�\%�s��E�>ם�w�M]/N��f=ϡ�2z�uĂ��\�`8�I��!���4q2�����̒钬[�eP�զ��d����/Ņ�(^�oAv�ɹ��5��@*�MwL"#$V�q�W���N���,�Z�%�j?�xRbH��W�F��\'ʤ+Z���7��Γ�U?K�g�FB�7v8���6/ONNK({~�yףN b3�U��_q���GoW��^-�M�!T%�T
�_�bR����Z�&�*��6�_�t�V�b�Iw5t�H���#�7�$�'����l']���i����E�9+w�Ҳ`r5GF.S3Ͻd �h���?i9����o�S�N��Y��8KRIS�d;��s�ԩ��(?EIj�R�My�̿7���,N7��:h��4ǀ�J���	�t<�l�~P N�����)W�'�-|�ZS�7{=b-6�2E�XҌ���b��رp��a{��p���op�T��]�*f��=	���M���َ�Q���~SN�����7�Fw`����H�Cō^d
E�m��nZ�<9
�Q�^�zV=������羪Me�U�)	)�HL L�V�bd�y�]�v�ܹ��nwش1T"Ys�z��%%�̄t�v�er\�{^O@=&AB�d�^XX �y"�Ns	�M0s���9�GSZ��g%_����X0ma���C?t,�%P��-�����n5���Y\�F�8�ph��!=����eX4���<Ї$ʐ8��xh���[���?H4��9��4i�^�@��Ȕ�\�<1)�ؒ�?�6����!��\Ov�������+;v���B�����bI'z_X��A��kf�b�IO�� ,�ԉ��V�9sRI�#P�Nzk��
��_��`��h��N�f�� +�J��e�����)H�djAL�M<^,��B�Z d����c��{9���H=c5%�CIe�J�W�� �NDZ���SN����������ĢM�b���gr'%����44yS��Xn���g㊪%�,'q�l�+���{�#9a����/�|���sss�S��h8��/��	�p4��h�^�N��^G$���;7��k��={����D"�Z���IS���ĝ�J=��3�F�g�H��l�z���4�F_m�K�<�+  H�T,hN$=1��U*�3fD`���iJ�!c �8$d�.�M�Ѭ����a��I?�
��$#������/<5��"t�(���1���+,oEW�3�k�AS1i��N��Ǐ�;/ɲ}ɳFQ8��E�U	��rjc�D��X$�/��H.^���O�/%1���#�I%F��w�	N]1O[��!���!��m0�A+ⲢP�z=�!w�R��q��1mKl��~׵K~�n1Z��t�M��n�v��Z�u���sg/����uΏ1�7�PK��We�i�=5)ZZO�0A�A΢9�uI&j�V�:�����a�q�=C�5�Vnc,��ޙt��R�J}(���b�DEW%MSUSw��c�+����ȱcǾ���~�#�*�I�����P 
�Tk�JY�[2i���j�~Is��9r�ȋ/���ǚ@F�.p#�<��t��&Z՜����%��K�����7�71�a@�b[�_��w�^����u�AO���۶oI��[K���<p𺵵��;QZr���,`b�36���ے�P�>�m��'F���C��"Q�(��n,�[���DF&i�Gui���7�R�d#)D���leoM%W���+�A@CXkꔚO1�����?��wFd::�{ w ��fLSt�:����o��&h��Ã�¨Ҕ�I�D1sHn��ޢRv�$Kز��(��	J;-�HSa���h��o�SO=uz�T��
��!�P�  �%��[nEo��V�߮�p�{��F'�V�&6�hPk�����8bue}dd��F�7;&� �bai��$?�T�*�MH���Tw]�:���7!�L݌٫Ŕ
�o߾��C�^I��=(:�2�0��X-��9�R���f*٤m]���F%&k~z:�cI� ���j	�@���7;;{��w�98 v�>Z�T�d����  !�@`-P� �:�Z~�9O ���ڙ�0��d����0՘4Q�2��.H���4xx��G�{�WI���r�������/�����7��Q�I����P�-�	��p�/_���?{����hI�Qd��9
B���"�R�����)�1Wp����
͑�2�~G<��Џ��g(�����ZufntV.Uȸ������k��u*&	�Z�� �ĸ���O0ov�����h�օ6ґ`�m۶�S>�쳧O�����Z[�P��J:m�a��*t�r;?$�����qpb� �5&)��ZME�KU=u��h+*�bY�km
�u���eK�5?H�����E��B/�qꍥ��k���]o���ێ�>���82JT_�����w����Z��Lt���De�u96W@j�R���Ұ}˝7����\�4����e|t��FZ���zP�z�O.=);aM��4;�ࣈ�Zš
咭Y۶mk�;���o��W�V���:]_ӝd*���W�n	�t�ږQ�"&`�{�䂦U%bUOI�6F<�⛔�(2�eUR�,+� �֘� �vE�5�V#J㌆�k�$��<y�R�c���������OMM�|� hF+�ʞn�h4�T�����%��)	���(�k W�~*��r-������T��UJ�����XwWJ!O
+7�#ZD�� �r%#rr|jjbϾ��쿦X-�W� 3b�V{��jղ�Rs�:�r��i��ьn���Z6k|�T���;<I���^0��88�T�^�`�
ű�kS#�ORJ�?ր7�Z�ގ��ڛ�������� �l��ξ9?>=�pi�cl�Z�*�M#U��c�sI�K���*�P��4�Wk ��#�O�L�D��M\'���E1�(3e��Q �[HCB���2�.V
p����Z�R�L��tFB���Ei�0�sZ�����Yk41Eq�q�}׽���Ɩ"@�5����آ�����ه6Y���%p�S�@(�~WT���	����س�v��\ﮛe ���$
�D���1/A��v�Z�@�8��'?��E��G�U-������fǺÉ�Up��7��Ǹdt���W�c�l�8��;���Jc%"�|$�S��y�� ��<Eݡ��nOݓ_u E��(F�<���cR���cR�]t[�}�-��HH��NJ��\���/���n��S�BQɔbd�+��Ƌ���Ihn�d Y��R�w�y'���ҪqP���(0�/�ܘ�=ڽ60�:��riD�=����A;�&��hvS��|R��0��(WF{}��	E���F�鶩dh��>�J�\Ag{��Y��5���V�$���K�$%�y3 'A��;a��yQ�$�o.7W禃>o>0���f�(86��$q:�@Z��$���|�Wˡ]�,W������7Ej�V<FWn��j�@^;�'i��� �A�@��'#1H��� 2�`��Bd��9����j3�����@+��B����^?|�K_����Ō#��ֹ�$
[�k�*���vu���7}����a�C��b�'��������A[Tm1�<��l����j��]���Z^��^_�A�n*V��F�R���W�F
n�<M&�=�o&|�@�x�&�hZ��� �0�=��P��[��f�-Y
�1���[`#Q*R,Ɨt��X��J��(f�)�^}�ݯe�5����TR�%Z4Ϊ�(���g�@�F��H�$丰$Yo�$�Y�X�*uI�$VP�(����%5^�jb�ǻ%�T-Q�KY��a�ۥ$	��{rS����B��}�c���bCK$fG ��,��`�J��"㘡�ۅCE�f�E�bj��j� 1��z�R��*�� ڠ��~��ҥf��p��c�	�G�S��8)��F�A|*Z�%��B[�(&
A��n�b��i�.8� ���"��,�S`f�[BE��8�]+v��u�"�H��Z�$w]i��ż9���{)���c!���cS�:	疲�L7����@[ˢ	il��
�P7o�2YB\�^JN��R}���?��O$�|�ʴ,�Ѥ�/��M�~H%���U4GA�l]�l3��p=�]�l�˴� a21	�Py,�T.�T1i�[gOv:m�4ݪ5<;<[�:�Z����va��+++���SSk�㓕jdxt 2��RC�%[�(��\��#G���`>�P��;�J��b_ Y�1nB�j\0G���$�5�i$��PR'����n޸W�+����t��|��$u�$�.U�W%U׵0 I�V �z%��x^//}�B�D���x/��Y�N��7�S=���m;��	E��l�'~�.���&�㉡3��G�Gc�h�uM ��� �b��	��B ��-�����h�6�O�8~�8�1=9s���G���a��w� o��p���S�������j{��ȶ�¾�<
̏�����G^4� �@L�N���=�\�<��FN�A��lSmD=����ʳ�����-ƩAtS()���1��a�N�82$�P��*��@�ٻ���S<���l�Ңv�`�HD�8JED���c$)���T�S�WvC�E3��ZPU0�^��e�}��gA�����I��۲unu��裏;vߔ
N@��9�R+�qą�C(��x|�Z�G2э��!�,;��:� $_�S<��/a�c����ɣ�._�<7|�]׽k����<p�K�N�푻T�&c{��V�Nr�Ｖ�� ��\�5G:ã&1}��J-��MY�Ծ�ׇ'���d��x�,֎{�k�ֻ��W�ahEiM�����!�:N�`\�u�ArE%�Q�ώ�h�$X<��{����>(�Xb3iD�*v���.�]#�Ӥ�%��\)��Q�Xf	���+�C&�%Hκ��$]2H��2��q�e
��NJ�I��6�"*TiH8�p;|�����E���`l�&���R5�&�1Rt�RZ�C�Z��Mi�.�YZZ��(�k�+�v�i�vϜX�2=�����;➳x�R���V��1�ࢵ�j/��zݑ��=w������.�>qzy���'�i9�5b���n[�*ˎTm��Z=�0$/t��DVV��>;B�7��AU�ten|m��}R�bjr�6Ta��^Y\j��,�p�=�u�f���g��)ѐW��لX���T�nKX�3�� D}���P�R�?���".$�@ �P��8�g��KKR,�
|Zl����sss��w�;��N*��Ǐ�����$x*��N�I�Sc�Z[[��Ĺ��D�Q�w"�T� ����m�:���G�k��o{����2�ls�on�X�ڝ�׍ɃJu���<��B�+��r�ŵg��8rlzn�X.�
�R�	O$S"N���h�h�3Y6"1�sI��PL�B�E���;���DK�ԇ;22�|��k��`Mp�!Ym�t�E?��{��������&��9{Oֱ$K_��c�,��`g�@ńDB� Yn$� ��#mKB�d����_-F֒�t:<fc \���0&��_�*
��Ǥ���얿�˿�������^�Zl`[�\��ɓ'o��F�*=�k�*�ǎnx@`:lN����>�K�"�)]^�??��w^�|a	�9Z�v���:��`* �X Natj:���ߊ�a�*�ܶ��_ZYl��F��,�mJO�̙ͦ�w¡�F�
#>WRm9�s:A�>(Λ��.��ʖM&o�s||R���Y�e�:�
|.���v��Y��/�y���W%m�%_�`&�(4��ǒ�8�o�<d].~�4�{�T)�qZ4_J����`�x�R,�C�`��3Z,��EK|�k����믃a<����m���������~�ӟ�tfjJ(W���$K� �=z���H!}��B&#hI�9�,*�g�Q�o�WW�&�c����S�瓖>Z�"J�^]�Ds��[�l����Τ�q�-�{�fc�h�C����A���k������&��L\!@x�j�Aq��~ꥏ%�X�
ˣ�ܒu3��![M�I[*�~��|
�}Y �������+�v��Ra�4]F^ ��ȅ�(8�E9��#p��$i���["lFz.�U��C��m۸AL�t.F$V	��:��SOMNNb'\}�u,��Z�X�t�� eT,H2C�!qM��'?y�{���~�����q�&9T�A��g"�n�5(��P��>>%ti荕�n�����n�[�k+PD06r��%ec�>�q?�֛]�k��F�K�.��Z���=*SU��v�g�^E�QLHu�C:b�E�]�� jd�S̢I��D��������?8�,��
^Y[os�u��ܶm�K(�]1��\I+�b�\&y��F ]=	2{�"�&�ą��ѷ��j�ځ���瞭[�b�z*s!1��@�%��266&y�a�IU9� �1I���6��)쏻��[n�����˗/}��Jc=mO�1�M��L�̥ Jt>[K�l_E�Ι�,/�F����s��k��P�^�),hdT7p�N�-�P.ի�_XX8q���� [[�mАX,������$$����kF.�҇"�M���m�'�P-RYO�l�xR���O��L�t�\/�4���/^��Q�D,�G�m
��H��R�!�]�͹T�wR�aN��L��^�*�#����jK���. ��s�L*��{�(_���۷o����/�-ᩂk���һ��r삤b��������z:���@h�rx ��������O6��aAgb]�%���P-:XND@��,,{�z��RV[�N	�ڶm�0���k#�u=1�]��q?����c��~�V��A�F���9�(�!��|܁����I�z�|�����&Zو��� �9�Q9�V��<V�ҭ/l�D�yh&�R-at̞�	�s*���+kR�Jf�z��I*���HRΙ͛I�guPL�R�ſ�l�39m�%�3�$��X\�����IO$�+o'n}�5�$X>�$�tF r�cz��$�8*;�����U����X���˗}��K�L>���F�G0���D�Y�Zn���Q'�mw�H$g��̪����f����k8�i�`�T�����Qz��6V�� ���R�Ӫ�Tdj���B�ܥ����Z{lh�
��+&���N�[	 ��FPu:�-��%�������l1�	p-���s���V�9�6�X"Y%���zŢ�}�7܂===�o߾�2���>�Ҧ.\�hKʵ���6���%�R�Pť�D��YTFV�_x��0r�u����h�J>!�\�<<4�u�QH[T�JH¤���>���t�c��v�%��±��P�Xe'F+���^y��[�M��^�����Ӓ�-��OQ��r� ���_��7,C22��;��\�8��9M)}��O������~͖-����J`��<:6
�l���X@�a�C @gqe1JB�;�4[��q���B����R�)e�*&�y!�L�mf��%���4�V�x�§�At*2k��|S)S�J�7	�t�M���E0e�QSQ�Q�S��d	زxzz0IJX�ahP*�I�& ;\������I �N�����)�2d�"ƚb �yGT�L�h)^ʜPzV6��mIdxQ��X�x�"sT��������{���M�l�Fd�����Q�ҡ8F'Β��b�������� ���2�iaJ�����hx����Lq
�:s�a[�v�����R�S����7�:f�٨�*ԝv�������x~�#&�FY�r�(?���X:��Fj/�9E�Q�)#EŘ$�-e?t�S�'�S���=�ȑ#�//����+�R�
Uj��D�@֐Y �2$�E67�+ibr��������زe���(=>N��ضHC��6J%)��w�^Hç���8�q�@U9!Da`R�Vg�I�.��dJ>��D�[f�%�é�b.K\*P	�b�P.qρ,��#c s�� Jͦ�`H����Qd!�������Ȥ��A%1ĝ�2�&%۵����5^*S9w�<z���@�������K�/C]�n%V�4�+�to��ۭ"�������KW�D�dM���\��8uS2��\�.%�X*�1� p��cl������Ǉ�h�k뫔��E��i *g�j/��\y8�8�0p����-�-˲6��.�����ɟ���Ǐ=��ر�S��Ԟ={L.�5=5{�ĉ/~�gϞݹs� Yh-�zI��2]�b���9FA���
b�)r],�����jmc�P�<��־s�v�J��؞C� D��2X}c}-Q�QF���S��>x��է�ГLU>{��ʈ�Fil��MQY�;�^�Q����(��ر�F�
����ǈ�a�K1�m:n!�yݳ�_{˵3��у�
���ë�g��!N�F�ӆit�z�(̩|�[
w3Z��:W� �DN��.	lv{�پ}'��<��:u�СC�u\Y��+I���.�=)��4|��7���ǎ���ر��~������=��sss���'A ��������p����7���t�Mh�{�}��_�4���ϣ5�,��R���֒#^�u��.Lv�BE�-Ȝ�~@Ț�M�����!m	e�X;��t��K�Iv�t��!��f���W��K�bH�K8,�l�岳�^R|[�܄�� �1��7B��ǁ��5˶($�놽�d��:+^�K4��`�򗿐���c��U*떱�ri��2�ub����n)�1�ˍՕ�z�+�]p�}B�r�*=!�AKR�zp �@�\v�  �RLFb��D3`Ld�`������G!����'&phh$m��<c�N,G�f�hP��~�����u׮=�� �~���޽���f���?���A�e<���h��~���]|<�!a��#5�S�Ƈ����ӆ�y%S_�����v*�ZA�X�b�����>ZK�D�6��"�t&���ĄmI]:�GC���z�ϔB�t���H-=41e������+�6�N+)h=�a�&�n�	�7P��8��8��X}��i���`u̵�Z����+T�SKg�]85w��ܮ��LJ���LlY�)�E-
�,
I��A��zLA�\�2�^N��2�7���M!JRM>�0�1{����e:m����		A�<`T��aCp$��1%�7�9sFN�����[�����Ç�@o{���\��9įЄO�<)�dTュ��%: '3:�6�$���&�샵��J���C�#Lc��j��8�����Y���ǏK����y^?�����X/��46��&���V(�8�J�d30���@�_���p�Ǟ+W+=�k����Fci}t����.,�O\\�04\��&�q��l@��ay����?9������q�������sU���xK\[���rQ�[��Zش2�)'u��~���9n״�<
})Qߘ:*P�Ӄ� d|����B�L�$��Ƈ�u�PIQG�H Y��oݺ�^���]��������ӧE��5+�E<rC���$�*r*��Nik�6|����SE�Q�7Z;�x�&����%D1��T��3 y��ETd�СW��`��f�D�V3/��B�*��ف�L-��7�F j	�lL݀�A�T0�$� ij��K�����O�9w����r�4V�w��5�uv����/9q���v����Lm�k�N��n�r2�Dlӊ#`Z7
��%~d@$��Xkl��E&y0b=���Y��8=ۖ�A�T	<�!t4:����  H�7��l�b��b��\������-�i�"�����*a� W�`'������l롡���IRUS��"MG�\�
~\�P�,��?�8�$:Q�/��D���JE���ǡm�kLK
t��-'Vhl ��CV�X4tZB �<������L�\�I��ư-�t��3���j1�ba�!�#�7�Юʥj٘�ӑ�/�%cF�p�M��.�j�����'~|i������>�ޱ�q@�N�E��op��D��G��f�fd������GR�R��J첩�����(ˎ��m@�T���?�1U��ש�aw;��;vC��êc�Τ������zm���Dm��X����5~��C֔	��:)��y!�Hu���'��$F�A섮K�X�B�&|2#�Ex����:��Z�'���s��J>��˗A��B���OU����@~�#�&=�Ӌi� ǵ��h�-�4j���դ:����#o�8�j��-3;�gz����k%O�c�v�J��+2\k���?W!�$nHbY`Y�X� o��V���}/�R(�b�t� ��8�R�H� ݠ�z)�S��yi`��5��7�xh���w�Cl]�PJ��� ��G���hc�ʙ�R�^��hb>u\}ɺt �"��E�����+���B�V_���3J��o>N��RQ6!iP����W�X�ҳ�\BM�/����q����$���#��f�DEQ� ��ZP��:�nԭO�T땰@z�]t�7L�N�m��¾8�bN-���cG�����.�b� ���ɳ���VD�~cJ��ݢ�w��/h�V�s�҂T���M p�S�3*TnKW�����cǎ�p�����fg�Oa�>�̓BsX/�e����wllm=z�*��b{KJ�dȊ��S�S�3;�=�����	�Celg]l6 �j�$}j�����é6�����m�CN��lU��n��A=W�/H�ʋ��4�)�Q�%n�I 6�h�F%ujV�ӷ,�ܠ\��g7��A3c�J��gR��G��0)݈�:iI��Y#j���]�,���!����Qr�-Q��!Z~�?{�̉�Ǯٷ���_G'�O� ��<�߈M��NK�
�Ǘ��%9�V��|v\���}/�� �@�+_�
T	[����?��s�|$����dY��m�.���M���u֏��N��9U���Tr q�0r��4.��g�ǁ8�,=�՗ň�L;)')�WAU)�hz�Q�гHA=K����[!��l/'%�'�NǑ�&eG�aI�7)�+�~/a��=?�B#Ԭ���x��`�X�(9©�R�JI��2'A�UW�*X�ޚ�(�'���b��k����7@���I;t���,��7���!��xk�c��4J������T��U�#�������|��)T!�Kq�xP9j�^D�Y�x�9JN�b)=����4$��kٗ��c������.A�Ks�, T���>�(�r���7���|�V�8엡��iD� �X�ښj�(j9�Xq#S����]-��buuy�^5��6T�z�	�Pڮ���.X<��-È�oeG��y�)'�3joF�vvQS�]�m��oM.�FC5�"R�Y�&?D�><;;])�HI.�Y�n�fp��M�<��D2��fkE�4(+##P3c�H�qb*m�)#G��� �E�d=c�^z�%9�J�E�R�9:���\�K�++�#�K�,um[����~�rKB%��
���R�^j��KqZ~M,����uq��WTc3+ybOj[T7M&/�US��d}�(B��xw̑c�b���Cҧ�u �u3́`.xr���0~L���{���T����eӇ<ڄ|e�`d�Ν�o��&F�$��4����EV�JrJ}�<$4�,�5���t
6�Z�������	@��OkW,�r��8��jdǤ��M���U� �����yU(��i�i�0�z�$�l��J^��� c�܇ke
 NQƠi`sP����(E;�����d�X�vW(�����w��T�ע�a�"�ث$tM:=K7}��HB-�ɤK%5��	y�ѣE�HٖQXr�a�����$�d�6���c��Q�W��U�5�mM��� 5F�Llup�r��S� �hT����Q�f ��Ph�v���VD�[+ur���:ۑ"�D����^�R$��o�:sMd�+�/
\hu[��5�ʯ^���[���9J��R���Ji�/D$UH�[[��r`ǱK=e� `�M��	G�-�A"'1�!0�XBE�	?,�E T���H+��قe�9�\�Z����;�m�U'�c<�3�����/�nX]i@�~��W}�
!%����*&fb���l+���X��!̞}�1�d�!vG�l�G\=�1���Ͻr�ylۑ�����-{��ǆ(a-���^��|�.��8�]Uc!NqW*'S��6���*8���1r'"e`��pT�l�R��s�6	/Ǵt;�a�S�4ٔp��ɮ[S���EY]AQ���őtp��fsHh,js#[��OX8p�+��t3i���Ɠ�!��4z��'͡��_�!5��&�/�s��w�v�����u�]Bxdd�����N1eG�i�4GA��)a�a-co��L!�+Gي�AL��t)Dͮ�k&DKlBy��5ݲ34�cf}��������-�f���,.,�={�����-�c��m۶�\��"2#/�M״"	=6��Q���6�EM�/�phW�5��<��}T����� �@F�={���.�t�Q�2�
%G����:�I����up(�˧����;*�DY�(��4 C�c��Ix+�(ݬT�������aF�ʘ	�ǗC|������q��N��YY�T��90̗�e�t�f��-��nx�{����o���g�y�G$膎�Ԁ���<�D(�,
U Z�b�I�rW�=2�ӡ*ǃ�� Y��/W�^T0���k���}�}�q2
�n�uilh���~���ɳ���WO�)�Y_j�~���p����UZ=�C
�TP����q[Kr���p�$�T�+֒�3Cm�g%�t��xrgbbR���Zm�^�ћ�5	��=w�7)x���;��M �-�:��5x��u���|g�-����������n���9l*�H�Ԕ�T�07�%�ܔ�Q(bˊ:ĩ�B\��F�pLKd����k��Z"�������reyU�&/;x^٤)�YU#�������̤�u#b�=!�i�H�����6��珞7=gb۬A^s���F ���r��V��ڎቑ��K�y������L��x�n2��$*T�Pc�oH}]�f|����L�<M�2��D�lUI.�SWE�	�3Q.U1�܅BI*xg�-�F/��eU�%Teu츞Y7R��F�'�P	�5�� %<ϡ��]��*���MH����'�|<�ͪ���r�F�o�D
B�|�M����*�
̉�l�WA�^�X^j/�ԪC�,���M�0�W���]��z���ْ��B J�[�q��'E[O�"����� `)�V���s���c����h�X*�@�׷��7 ��~����]"̩͎h��߉z���^~s����;'0] ��PL�$K|���TS�YJZ�l1��e�bz�Ä��[�OA�1�o�F� 'g\
�&)�jvB�V���!D`/��e�Zy�Zϳ� غT�V���B�S8�@��0	m���LM���Y8S�^7��f�[QHy�,�i�vfae�k��ۥ
"Q�AK
�zyɞ�1쒿�����'>��O�_��_1[�la�킌�������{L<9D��/�q�N�n-g���o�dQ�G�N�ٳ4w��^7�H����?pͥ�ةK�f�ׇB���Eg�d�tb_?z�X��z�ɗ�)�Z�Nς�<�%rĐ�X,%bQ59�ra�'��j��pBf*o�8�-`*�/�<>>�I�Ck^�ҥK���:�%p�[h��'�K沿e�3%$	2==���1��`E��ߐ5sss�U�&ծ���Rb��d��
@	�SAq���*�+�Y�T�+l~�Z�^��q��]�,�Q"v-NB��XtӮ�ɳ�r�	}�;r������������@D#�t�G?���O?g�WZ�&0�k���S�H�f\��G�pD����F7^s��AϷ�Mt���*�r�<��� �hE�n��my��pud߮}zbx�ڑW߸����*�ғ9U�o��"e8ޟ�g��a�nJ�����T�c�1���K���z4�Y�� �����1��iQ.�-����V>��ȬV�g<�{�n ��K@�=����_x��^{��Ї>E,�^�<��E��C=�k�.���Ǐ?�䓇��P�w�q�u�}��; �� �cȦWp�<2�����S�N�ɢ��uyaP-���p��v�z,ׂ0������� �M&st��I
�\�����K�	B�~������xۍ��Z��!$���э��y��&�kAl�~�.���5?��f'N9�^n�NM{~g���//-I���1���:�w���l��L5�[s�k��˧�<3:52>7�ЍR�8�zp�1�YS�1#�h����-�.�N'��X����D!.J�oF4�>a:����>01���/� dU�$҄N^��#Ʉ�sD7�ʦX������ѣPg@����-0�O��oan���'�&���������߀!}�3������.� _x)�H��z"�^�"�djl������l����`!�R�RY�\*��E�3����K ���W �t뭷rqX"IlL�K�1��~�MB�YS���Hu�KHpF��Kt~$��d˒�.��:�*�҈9�t�r�q=ûx����8-r���?k�����۝>�`��>��p�թS���uO�[��nEdW��</;�[��X,�m/ʹ22`sQ�d�!J�����",��򢓹���@R��+/����ᲄ�)p p$��5�aBd�8�%�a�Ν��}��=��S ���;s��?�A0�=���~��>���޻w/~��E�)Á��@�!�V4	��ٷ�SA�
4	\�I��Y#�8�,�Q�'Pe����}�{VH�*�H��~�s����Bj���ٮ5���D����a�U���,�,C��i���4������(0����1;���T&�&��?1:~���.�N������a��;�p���P�"���K+����4�,Jίqvi�Zx��6Հ1R\6�9(������\
���ԙF$�f�P�L.6���Yj��[�Ɉ�-���HԁdwH�}�qvrr�C��8���/~�x�k��B��Da��@<�Y��ZV|�4�ʫ��%ZZ �$�H��АlcH	�b��!U2-S!��)��7� ���o}�'���)�����'?�ɯ��G�x��d3�o�X��Z{A�چJnm�G�,�h��P��(�~`����GǆG5?	��\�P��a�v�H��v7
�^4��\�LLL�ԜBۛE�t�.'��]
[����7��;!Sq���a��L��"���g��+(�����4"SccW��ӼW�c�LM�Ҵ�A��t�`%�2� ;
�yek�&�6p?�c��F�;v�����ԛo�	x�����GE���Sd=�b�X����j�[d=�&��@,�wR��R.K#�p*)��~�� ��֤2	�I�im����e�:q\q�y��?t &�h'ST� ��`R[�P(9����3t�Q�١0b�\��h��{��J�
���tM64Uu=16��V:��1�ء�y���|�*��8�L%9j�(-��R����R�#��y"�Y'"�Wd{�ph-=q�v��L6&��! �U!����z���Ρ)0����Ν��,�r>�2��[��I�X!_!i����V�NML���\��β�C�VWW )�Y�	�%��;�T�π`���n" *޿�Aq	,�l�c� 崖d�;/�c��f�SO��L{2e�����1'c�#+������to�i�1��N���_�x���������,ֲ�:����٧o�9պ\��m\n�a.y"~�劷Hy����)R��E�D~EQ"%����U���:u���v�Ws�1ƚk�}�r����U�g7��s�1�1����bEC��ґέsܤ��%o��F6b;(��(�9J�)���$�G��yA�^��u�O��+8�J|x�)%�#�L��A��t��ٝ�iM$;�i	�A�C ~��կ����_�� �*T�Yj0A���>>�l333��!�xX�k�^�O[��XX[���o&gx�#�\n�7' �*�Γ�YNa�iś��ׯ_�"ȂZy�����~�n��*5$K�t��n�u�Gd.ޝ�����n�o8�]��"�񑣇`�vv�8��T�hJ\0� �V֗�$�jx4l���[�D=��t� -�
u�r����t���V����xx�6ʘxr%#����8��uc��5D�K�����D�c��s�����9@�S�����pɟ�韾��/���t\���ocp0���ŋ!7�FG��j���P�f�4mJX���Z����J�U�l
7��\,��k�a�h�-M+p%8x���1R�����OC���D��;H�v
e�=��׀�Bt%ژ��%l
\�h��D��7�ps|ο$ꐸ�U�xem�R�\�Zm�+��R��!�U�mW����A�*�Li�'���,b�*3`v��F:{@��S�S�~܎#�ZGP�L�!�<����+1!U�&�kAJd}K)�JՕ�l.L�$��m�d�ixlD�T!j08��׿���S�`}�x�����h� ���:�^�x����sss׮��O����AC�Pu���Ki�_�J�A�np��e��E�ɞ,т.-�̐~������Tp� D�Sg.�f�J� 4�q�?��L	��������}O�}���%b~��
BC�ia�$hm�b�21�JC�����?hQ�d`ĺ�p��S�G��n��`a��t��C��Q�>���W�S��j#cn�m)���V�M�>~�Tud�)�q��O�.�"d��ӣԫ��8+S�����W�$&��NVFg�d\`�49? ���h���	��FQ��B����B����t�ޥ+D���G?��O�ӱ����z�X�T���{��Ϸ�x��ɓA�������(�����Ż�̦�ٓ�o"0p�Q�͠]��dY:��Bt���� ��X+k��f���ھ�x�*��c1H�/}�KiƂ`�Aυ�Ǐ?���>�1�0�!��3?�B{�1f+O*]���\�2�S�C�>e]�J�@���p�\ ��ً���C�Cp�:a�S�K��~���]�S߾u������d	��Z�x�@�~��6�?���&i���,�����ZD�o� ��C9���;De��,X���X�8%3%�^��J�㴦X���m���Ճ??!sg����=7/9V�n�h����E��{�R'%�����%ɎA�T����	ǋ�d�x�:RL�B%�M�ԓ5����ڲP,�\�O�љ���R����	�`4|��?�D;��O(�˂�H��.$&u)w5�\���Z�9��YA�-��Mw�P������!��k���6�:�����$�ǯ�ߍM�Wnߺ{�2\<z|�R�@[$&��w++�g����e?'a�:/a�n@f��y��p&P�?W�4<%���|�"������I|a��U�k�Ν�P���T�,ӵu�m�z-�ݻ+���D �ʐ��ش�>9��!4�ۆq����<���c1K������ma+$e��s@���-�"�
�%W�>`�Q(z-����O�<+�����28;.c	1�u���eG�NE��4�D0�én:���+�3K���_��V��;ր�
�v�[�iO��㪢�۱�k�������ǪC���������.m�l>v����`Κ�T�Gd��M,M�o�	���ӄ/	Wi^2R���;���ix�x1�A@����?��@V������ĐM�q���^5���H`2,d�vQ��|9>�� �z(��2��	�}V�3���d�IE>��.\�@I>�D���|*w���/紨+#6���}@��`���.Ҳq7-Ҧe�,�y�©��>ք�� 7�.]z�G��#�پ�@��ף��N�M2�m]�˯�i��*
h��~���(=�
±�Q�h�?12��ފ�0v��vͫ��훷/���=���g��I��	3ų��\��d>�5^0�$�qpB�H�9��������L���S��P��f�M��^�(��F�Ǎ�Ngk���e��-�^��]������&�ED�q�%�&F�m��m��,i`L� $� B�e��:H"�v�g��H`
j�z�P�&o�J��E���y#����q<n[g��d	��8�	\���ۍFS'���'axe�c*/���4�
es�Xe��3Yq�t�$�Ɯ���	�B���׮_��Q�FE��w��f����B�Ef{m���o�Z;g:s���ᩡn�n5������t��w�
6ث�M����Q�"V9��$�ɰp�~t�m�����e��M�G:r�0�h�Q��!�x�~��n�j��'$�L�Su���f$�5��i�?�Y&�\IH,�E=� ,�{�[�
oY�M�lI�Q��'�E
ǩ,�[?��b^��b��,�H��)�Hh�ټz��3g���/���O�=@�q�}��_��WBbK|ά_´ї$�R�$�+�TXji���O����.��)�5�ram�L����z�ٸ37w����ၱ�[�t��w K�G�:7>966=�N��fX���3V/`�G��Č�t�
UM�TӔ��ߑ�Y,�f��$F�U�:9#�195.i�pw)M�&�����$� ��!y��.��	�^�-'q��L�C�:o$Sr�����m)�1��U�,IJ1rU��~�n &�.�[����l-���A�H�DR���F�ou�D���[�4�ߗ_~����k)╺,�$�HB����*ժ'�1IgƇ̵ih	��j�5�"�j;.V;1����������������RhD�[k݀{��Q*=v�p	�V��6T:�K'
��J�\F/�g%m1i���VZqR������6�L�xi�UhSж��֎��?�wڪ� � +X��u��^O�lA��Ȃ��徱�nY+�#_��`�o��g{C�m�,�e:t ̐:��W�� �$�%e��sy�R�m��.fk0�(iSȲΘ�6U�<�FHf�@I��뿺p�^�I�↟�f�~����*,ZGr��e�Tք�R�e���'
��H���Q� ���(Wێ��6��b��>���[�nux�ܣ#��A���0w��t��s��ǳ��WA�+�,C�8eP2)<\�5f�M툉�ɩL X�0��Y7�v
��t�p_,�bXfRII��^i�	xE��_�
��KӇg��j
f�6N�h������v��c��p�6�,ӣ�j��2&�xv�kJ���Xٶ�T�Ί�-F��t�N�q�	b��DL�����m���*nRp��h�ԉ��:66F���oS��;P:���#�\��� R!xQ�z�v]'��)�PA�8�ݻw�K,j�AV��"1%���=ѭ��¤G#�kt���-ȩcb3�톅DI�����,�Su��U�Ď��(G��Kf51�8�urL��i��s�!�_��t��۷�{�y@��=N�R~-ޝ>���b��L�-@]3�(��ree�E���"n�i�0Uo�JY��#fr�v�i�i)�$?HTL��ڭv��0;���i����BOH+�z���jy����-nMphf�8���PzĒ?*UK�Yp�p��	��H�C�ܥcZ���s�I�)<x��mV(��aG�Z{�Y�ohS*��ٺ;����6��9'M���.�J�OZ7��Z{�umuiph`��MX*��Z�X�J�3K�p�o�X�Ԉ9����C[�y�ߓ��K�<�ג_=:<���OW*%�>���a���V������N#N��A�i8���ҢF���v�.F�E����E�=	�͛��+S7�;h!T�!��'�|��bι�JA���8�ҏS&of;�9��Q4Ӻ;|X�>��|ؒ�@��2q�p�
�c�v�(�[��R5�\���5/z��E�f�>�V�;�2�tb�+�7d��r|�N2Pkn�NP=��P���$*�K[�l{@�i;�`r���䱶$ej/$���-�����ۘ�v�S��{�g��R�����V�����4ba[�t�8�wG�}�رCS������7nH����k�޹<��f����&5+��r�
�����|���]��U�]b"�Dw-��X*��͘�3@8ғv�a��������1��)?��XA���ji�"^]�sſ����Ҁ%F/)?�$ f.7Őz%�+]�N��ٯ�#ՉQ�ܰ7��������r��n*�1v@�kq?P�f�������?@��KMY��9�F�E)t��|�f�|F&hul
lomx-G2�n��a�c��ZY��l*��o�Ddh�����B�贉I��կ~uzbruc��ɓ�����t|�+_����K/���������!(o���O}�S'N����B2t����~����f���OLLL�b����$�dS��t$ip�,/���L��v�"ZR�ew:Am�V*�b��cYt�hpdz��[GF�
�\�$S��?뺛��-ʵ��:ߐ
7�
W%��{�L�̪9��x��2�v\.�m�T�^_��	l��ѡq�me}�Zju۫s+�SaL.<����2(�_z���;�mF����,m�ٸq�:�)m��-����1��W�6�C]'qOŴ]�-�*d�S��f���o@�_�p���K���zBs�̙��������l�4�ls�愷� 	;r��3�<�����X5d����S$r[r�%N+>MĄƦn�I�l�5y�cpv�O튃F�ߒ2�SCky��& ���ť�E"�TiI2$�S;��̴�y��������fe������ l� �&�QNc�540�*���N(�<2K7�_����83{�U�4}{����[�AG9��6 2	v�O����M��$@d٤L(/��i[��)���*�͘��g]��xz�p�}������uBy;��}�����?}V�����^}�Ua�?��?�|�ݺ-N�lA����y�A�p��9�&I�@ ^�Ό�ױ�E%'0)���)��}��^sJ(��R� �X�t�PhT�K�toyu����`��ŋa�u�V�<��y��� �m_��r���� �,YUR������C��q���Z�f��?~�3��]�Xݸ�}�򜭤Uom�lߺq{hd�����g�t� *@�'Qh�f������(} Cڅw�4Vr7������n����n��qˮmw��#� &���������(���i�)��`������ɡC� 4����o���ې�q�W\�(R�U�����š|��"�D���8��� ����1H�«�
sE�W���sv�KD��.@��"0I<����?R�JW�X���W���/	��E_��ܦRB�MjiIY�����QI*�m�]Lb`��]j�CTf*H"�t�d���.�
I�8z���;+�E��Ju@E����V�ywa	�::6~��X��sc���ܪ](�>{��ܡ�kj�Dͪ���x��+-4�En�G�[M�FO����1T^��b"�� f�Z~7��E�B�;D�AԱ�b��?��ݻ��o�~B���]"E-��P8� 4�����w�`������Ŕ��O_�L��M�ء�'�X�c��!�=E�a����/�˦���i˅�lʆ�,B��s8�$�e+�V��������Hv����[�|>07�ǟ|&	Ʋ@��t@f1�����;艤�P�ҕZJ�ńD�G���U��!�/�ҎpD�=8�n�K����Wo]�9Z��9����H�X�ټy����V�둑i���wn�;Ok�v���,ӵ�@�*�f�s/�V�c���G^kf�����������m�����&���v���3����N���ϩ'Y��f��%��@5�q"Yl�`L�o�������|�W��V?��[o��ܳ�ś���^��I#Cw҂]v�K+�%�A���6�pD]�Ԩ	�0���& #$4Y�l8��#iV��ćD�~�iؠ�����7뒓������˿>�.��s����@�����P�.Ӗ����e���iZ�!�"a�CLq�u�V��/u}���9e2�(r٫��7/^����v�g�<�KW��k�yX=X�,�b�BĤ>��g�G8� L����6d��آ�J���w���t�X�r�0\׮�Cn�ϡZl⇥E�X�HhX�F�H��W��ld{��ߙ�_��o.�����.PfK"�|�8���' U�/_��y,o8(�DD�=M.j�MC�CgUQI���Q��*)���C����[�`Ӵ
NF�F�m���?�K`z �A|�[߂P��������0��oAK���%�X��@	��jb��L{�q�V�R/��tP#�d׷Z.��nT����lo��;X,Âډ��|�၁�v����9sh
�������[o��������'�è�p�=3Ʀ>�~ɀ�ᦏ{����L��m�޴�	��bπ�jb�v�7�璌kF�r���2tft�cըՇ��C"�.1O�/8����{�S�N���+///W�"fhZ�{]Y���ǏC��Q�u��%��KKK�>2ً���$�rq��"Z�Pt1���(fh߇ ��(Nh��|	��,Y%R8q$�X�h��s�!I3|�ɠq�-��U��1�
�QL�˝V��jW����n!	�����d[�`RЮ1荬�ע�vū]i ��V{���܃8 =��y+�k�NpΜ:���w�ַ;�Ы�f�-������=n�������n��$���W�� ~1@��*��Q��J�m�tl�o�pq�WCayN�_�Ŭ 01�0���o��o�w����K���o�U�
�mm�A� (1)Bǁ�{��a��s�V���D������v��!.O�.�ҏhuuޱ`���	�\9C�7q-(�7J!�4��/..B����/o׶�z�7�x�96{�u��U�N+��1|�1�.q�F����R,�,���)u������јQ��n+9:>��ŉb�p�vT���T��0�{�*T�*z���#���r��2��4760tޝ��Ö[ֻH�a��սO�.�q�-4J#n+
�D�� 3=��ѣ��j�.у��9,2�~x��� X��CI�:��ڨ �V!X��r:?{��E�bR����w���;���3 �# ���ۿ��̑��L�8%*��H���[���H�t#Μ�*Ǡ�X�1�����35��lA`TϜ9c��V�R�n-���� �P��<��ݻw%
����O~B�^�L9���aMYæ���z{����N�QbL����"���:1#m��%�X_o�Q��P����Q�s;�ȥ}P�����ܾ[�&�662�S��՚���Z^[Y;Ҝ�J���1�g��)L��
��@�����1PzÆ������EJ�m"�W�}�������:G��(�N�PAA3%jlx���iD �K�.R�VyH��"s_�t�Klml`.!F;�tl,{���,~)KS�'�Aȫ7��J�\�/ȏb3��p8J^���	?�-�ҥ�29Z�W^y�׿�u��;X�������&�&&y�i�Xq�$-\Uį��kk�,ӡ<�tki���TJ�������S�3�kKQ�}axh�u
�V�Tin7 �]'��(m��"��˙##�s�\��(����=2��d3�߭�.�����Y�ѣO���`c������o���{��������,~��ÀO<�8��rr�(g�+��Yz���p`��N�i)�P;K]0��Z���r�e���I�YC��f�B��f�����S��ԏK3�pQXن�^��Xb�T|��}�1��Iӑ��:D�?���e�b��0����n7)	=�JC�h5eK�w1|�P�S�)�t�p�[�a +�[.��f��,ߩ�6.�e�����Ġ2�R����������N���̯.�1<2�֬Gʁ��C�c:�bjr�p"6����m'q���N���v7�9�(P�f)�K�y7�T�qa_L۞�>\�����1 ����-�F�&��[��Rמ8�b B&੸%�*Lʶ�^^ٕ=���:�ڎ���0���D���4M)��J��;�D�B��r�d�ţ�rr%�
��
H��I��Ʃ\:��N��x�iC��^������2_ɶ�zJ�K�;w��t\nc��2�h
�LrפK��eh*Ma�S�Z�!�jS��w��zX߮V66W�G�*���ֲ�#�^����v�Z�R���f�B��Wk5�A��i�� �Y���mc���E{s�Y!̌�{e ��Ձ�^�����;~b�����vjx4ڕ�'����^whhd�2x��틿�D�q��z~'sS��V�k�D�����&����N::b/2}��W�M�I��s�;}���ض\,q�Le�0DX�5hxis�mM����䖣F���߀����k��;w���G?�I��1���a%)��	�����Sf��bL�U���h��28P��m�ݚ��hGCC�r���aJh-�ޞ%��7�6���G?��)H�[7v���3���P'1�0L�Yt�:��݀H��(ǡs�p(`�~���xL{��^�Q(	�#>��X���&����q���m����񅅥B�����:[&Qә(]5�&<W��)��3z��l"Q[k��D�&I�c^��:���R2
�+�����7M�,��~��.��H�8S�f���n*�zT�Gq�#m������^�)}��w�����(��Z;Yia[��s;���1J{�tpK�a)�./���&�E!G*��
����b�V���Y~�۬��b2V�6�����`{�}��\�o�>���7�;ۭ���N�g���["��.�ň(,⢼�y	x�{{$�̒����[�b�� ���#N��V	�\;��\+)-(щb�郹܄g(�_����A��3�u���4Q���(ר-�@�����L������<(���)܄oOlv�2�0���B�@{A�@�&�|pp�-� ��~�����׾)y����Ksr�����d�tx�^ms�(;V���$�NQ�O���m���z�T�)^چ��
f7gO��Y솾iAyR�-����a6�
.q��[swo=z���i�O�斯�7&����w�n$�A�}�>�.�N��e:�+_y��/12�DD�:P�w������R�����U�d�Y@B�7^��ܼ���ZP�k�t�:L7f��O26fN�rZG��������^I_˴4�<	%���Ԅ�wxv����t�\L�Iu�S�� 76�Ҁ>_ц���CnO?�����<��._&����4nn޼y�����'�Ԭ��ʆ6$Ƴ~BR˩m�nY�I�q��@��+�W*4w:���3#�9-������i|����o_��V���k�����c��՛�ܺlx����� �v�c�ۖ�&�I�$�7�l�'�����G���1=��9�Nc�TK�(���#X��&�,x���ﮮ�⋼�%���bp��*HtI/݌cǚ�T3��%�4�Qzi]�.���L7df�o�.�Ɂ�R�&��t9��tE�#�T鞆Y�SH}������26| q�:�p`~?��O���#(�_|O����n�$iA�.�I"�Ε��C�p��K��}n�C�ʶܝ&%N��,�53��ݵ�ÃC��N�j5�D׏�����q?l�y���<�q67����ã��O�-(�Ċ-҅\QEu�$EDD%� R��ň%�rՒ���%ï���F���8�+�c��&��V�ji�.�t]v�R7>I҆	Jvd#SGd�<�d��Ͽ�s�'��4Ģr&3+Rά��̜\�qZɎ#-o.�uc�L��gv~[~	���s]h�#\�܀��j�K��DeDo�i��T�%�G8��<iI4����b���ƨ^�s���3����n,l�sƵ�6�K�B���Gf�ܸY(�~��?��K?��+��������)�)��V�X��T}�źIⅢq�'L6�b����^�篇|�̤31�؟��U<.���cǦ����a�����V�V�����9�GB�%tL��z���I��VDu�H��n�Ss9{�[�I&C9��{�߮2Zͯ�Hǐ�a U,��H��WF��l��Qk�j��a�"ƈ�c�k�~j|bmyŰ����P���\+U�D+m���D�uR���aǱ<�&�<�{��t5�2V��)�z�CIŝ^���­�c#��ʃE3�C/���n�&��l��?yz���R���.��7�\l�Sg������Z�i���}�4��J�Ax���[]��R-q�%�8Z	�xɀs 1�M��(K������T��0���0�����-���4'f��ư�.�uikk�j��<�{w�0�MI��J�.c.Dv1�X.yn�͞�O���^,Y�� θ4'#�9�C����t1{�X؄�e�>&ո�*�1�O�K�e7��:T�TM���>���x��t.^�8N��1���ӧ/\� s��-�^���qv�N�J��r����u9̣�w��-�L���!v�ҠѦw�\H����Y�/�/�nO����2Z��x�'#����n�]������� P~�ܹ#�üV�&=��PӃm�����HZ$�~�t��u�:��W��^���`�!˖�|��kI�b˝�-`�}�ZE��H�[\\�%.kT8G�Z�|$������J������G1CS4�d%3^=3�HS����f��8S�P����T����K��~�;߹v�p:�`&���o���S&�$�B�MC~3$�3�<�h)����J�,��r����YnhS���Z���ëk�^70+��T�X(O�ɚ{���w��-8�vmnin��9<Y���NM���C�O����$E�N�+lno%��2�(�� .��́�(�n�i�c��M�B~>��Ț��������t��A�[s�Ԕ+m7�o��~fN�n��~�g����*�C��.����y�RqAh����SO�$I�N� �%b$8rD�F�.�6�s��ܝ;�1�;�>I*�26(�Pȷ!�מ�I]	�S�d �B�[�d+�vO������JI���ހ͆85Z�����=20>��U����KE2���������=��pttx��d©<��d�گq) �.=�:@,���kB\`D���G+�Q0`V����F�u��ە4�>�k��B�,��k�
�Ŕ �J�7��W����u���d�'o�x��Y�)r���n셥|���zƙX�>�z��J�h��:Bk%�>���Mc����s%71猍MNN����N=zT�/�}Hl��{Aq�.�� ��%ٍ,�Z}�'�DBH���,�X.X���k~�^�Y#�����ŊW�v[nѵc�Z(c�k;X�ވ5���a�AP�R���fc�:��(j���L7D;;�Xl������/�*	��؆�
^�,�'��P��ٿ%o�26�|��37
j+��?dƩ{o1d��	�J�u@��~
�2��� ��$<��"��Ǵ���?�gH���%��5�o���J�}#=�Z���_���~����u��<y�th��T#�j])!#w�K�˥R� ��R�d�T$�:Kl`.'�;p�V����-�܌O�o��v:�F��y���!
Ųi؎90H���J7��O+�2���H��S$��� �1�@��^�M^����p�֮�0J�lA5�xx�t�I����;ԛ0.���0�O��,�E��� ���a� �J��ɟу��}dS�w3��N�,��p8o�+x���Qi)u��t��rZƅi!�<������v�;awiu����ō��}�s���7��֤�����_�q�l���w�<f�� X���*U�@e
Eˈ!�;[��ҁR����2l����q@�^0u�y�l�iƲ<�\4����y@ĨvڒZ?�(�J�whT(\
YVPq]?괻���
9�%��đ�����'��Zupxi~�: 2���czt��N��@!�����BS��O�M�÷�PI�U		�z��^q1�Q���=.L+��)�=c�P�r��	�e\5i��dײ�uL��{��������?��?�m�N�6#�%:<�'J�[��hbl�T�ll �l��.ᖞx�������5X7h���XE����~�C"�%��±cǞ��'�ꚆϚ�N&�rRB~Ѱ;��v�x+��9�Tʕ�����3,#x�^�T*���NpA����)_�Ņ_��՛oߝ��X����6�k�!�A���g�bȖi/b�räؐKM#]��)f'�]V�)����{��^96��:�2Qa�$�ݓ��PBh��{YJM�Brۄc<�Z/P%�y���v���B��m��(y�'�7Azj	�҄��~:������~���^\[r���p������P��
)��儛��E�Ȟ[��P����je��$��m/�)f5,���R�MO�de��	�+���`Ȏ+�����I�����U2�҃3���[U��Z�<68>>��Y+S���_�.7D#(I�Z�����(�ڦ�V��"��li8��|=��u�b��Oޫ��-O��EI#1���L�DK��=0:33�K+�m6�R'�4��%*3�M���F?���ܔP5S$w�N�CF�?N{T�6�#�AE�I�,�潥��,jN!�h����ޝ_�iK��i�9thh`(
�����p8q߹�r���U��S������ͻ��L����$8��B�$z��]d�۝"B䔾�h���(�dr�49P�^�CO"(�Fŋ�k��v���P\��K.R�H�Jv�3����>��1ֲ���.Ug���H���;333�W��cG~�#���G?&uX]]%^��h	�a���vʢ��|�G���Ӥ�^yF;�p�ϔ��ڎr&�<PrAa���ZL"MZ�T�>H@uxrS�`*e��i�4j������`y���Y����x�wR⁑Q�[��M�8�S-\&�n�s1y��1Nw�x.�pP%�F�g���H0�ׅ��z��'��5N,/���ӷ�o�g+�V�(K��a:����cj)Q*m��'�}#��0zz���!���%5C�����j?���x�C��WVVvvv66֤������=E��CA\�r�����ץ"��BFYFos�Y���3b�}���-�����)��8�k�#��1w������R�joE��q��4�"����R!q�X��Z�@�R���%f�����X���ɹ�i���:�)E%��)��mJQ3=%�ޭ��<~nsc����#�U��2	wj�kW�����=�@9aV����^i�#�x4��SR�8Pk;އb�;,{f������C>��s����GF�����x����C���&aҋ��<���0����<��z��7K%"���l��ܛ����:�d�a':�rz�8�:t�\{�p�y��D6�T�iG�K/�ts�hM�����m�j��7AI:�Cd6{�&���6�� K��I�O�Cb36����Lt���匸���Xmڲ���ˍ�0.
r�"eKZ@��P�+)<��/)$mPqG&��̫�d�������}< 	���� e��O�X*H�b��'��3g�0d��b�c�e؄0�-hH�8�pe�����СC_��_|�E�c����f�1!ٸfp	��Y�����1�5�!�-�L���T�ƈZ(������r��"�*�(��%&�q��� ������o,���٠�.���K�B)i1�r��?��d�0m.�]�~\p�v\pJ�S�l}`�(�-e+I�&63��#7�N�� �&���(1F�d�L!�͟8q���@�K�fgg�M���),Z��H�b_�`�	�	Is9��=��?���u�1V�-i�4�:ł"���+i�f�n�x.CG�Iڹ��lea ����M:���.��������1|�� E���d����AW+}ο�f��dz"�ml�;J�"U��q��k�a{z�4[q1���7���A�,���<� �'�	�?e�$ڥ2��>4T�,i�o?��G\N�:q��E�EԦ�R9|�0�@U(b��N��V���䦝ɏ:�hQ���e�Gy��_�����K1�fd�'<02�i��w�q�?)�*� $�R�AUH�+��"�8oePԨ�yM�Ɩ��sκ=g��X$"��E��#�>�^��f�D䃌��]35Y|0�b��Ifk�/���J׳H�lʿ��. �F��q�
86Ղp�so��D(�ed$4�/4�S�p��ԕ��p.����͛'N�����T��r�?��eZ�2�P��ޣ�l��㓕J�������ϟ={V*g�k�Y����#XL��M�D<���R��9����$���,$����;�Mx�gg�`�pfZ��3ETe���,ڨ~W�6�bBwɣ�'s�,�%-���UI���{�J��9.CM�!ô�&��/������s� G 8M-ά{�|7~�q����}�����0�q͓��J�!:��O=���9�����������'ؓmt�͂K�ˉ�XTSa��PL��ehs��S�:䌲е�ɱѕŅ������[[;�J	��iSr�;���:�d��M�M�,SP����tǷG�H�s�%��+x�:d�A��~3��d+*�g�w����$V���0�Dr�*���(A{C�t��j����>\F����4
��.�±c��o��"!"���=�������.� �HC/��S���f#ȕ��&S6#�t�,�������g#Ii�ϯ!���P�=eS�����:{��f}t��%���q�p��%�B@[ܟd��\���Q<4����d��>̣ϻ�M���Q�)�����g�}vk��BN�:%>Q�3�-�R~m����Ĵ}b+֑UQ�i!�A\�?/��l�{��v��J��ؠt.t:.����؆t#�̝�#J?����ڕk�T������WJ7��.�m��O�'�q�pS�����z2������(}`t����a��#X%�\&�Y(�eK��a�(��DPʦH�FvW��`E`���V�빔���.��8?�Ԑd�hv�Q5D09*�g}�%��N������b2l�W����_��?�S��Tm$=R�<Hg���k�j������7��91��J�n$c�%XۥI����h�$[���?��w�`Rgff���v��D<SA�nj/���$2�iK���4>N������⢙���T�N;͊�oH3�k��$�������T����&ƁB��=���odwi���J�b�SJrݞ�إ�Km*�/E�}݌��#%��;�I��6��g<���8WID)$�Ǎ�T�	��K�Ɋ��t�̊K�IH� 1P0� j����iw��a�HL�뢩y䒴���#ѭ;9J,��g_>7If��Y��q�+����w��d���6�[��=$�bR���ߑ���w���MP����~zz�p���8�%���Z%�-e���ő�#T'���3�	N+��\����Τw���j�o�$�j�_�1��w��v-�+62Đf�+eZ��'Vy���h��رʩ�tb���O"�B4��<���@�J,azE���q&E(���/��d#�J��5������PZ�WVV
�RƟ�sL\� �X(�%�L��X�R�M�����%������dF�����T*�7���ڮy�Lw];"1�������zp�3��"T�^sÀH�n>{�� q�;n�Ο/�����+ZWb8d�E�K����8��Yv���BH9A�f��Fn�2�;q�K]�kS�A��7�����<�@q�D�
���:�1�l�����#�$'��\e��;�>�!.�~��󷺢a����cc�OLL vHM���a�e��LIY��&	U��QH��4R�(�I��$$�ϿH��>q����l��s��'�}������p(%��x�G��Db��"�(l˒v�／�MrY�R��Pv"I,��܋��^62����$w�a�8����ػ �^C���=VLG`���l���������]'�5V����w~���Sw�ԩX��p�M�N�x-��y�[Y�r�k�X��fR���3L�Fq_�r���:Ͽ�V�w�{P{%��/'��^W}�#�m0ў���eLF���(���Rvp�7�$i���6�A�Е�`�[���5���CW�a����s��HO��t����=D��(D^���q�Ӓ�}%R�Ѹ��t)8��ԥ(����>��th/��F	���j .��i=�#�������'>�jQ�r>tE�a�p��|�(P���zqqq}}�Z�23C ��ޞ2�
rnG�2�X#_�.�kH���r�^W:��t��9��;�>�,1:�߂� S-��0����Gɮ��=>���o�+�X��Ɔ}��%ى��{���}�}�IR��h�E�;��Ag[[��8���<��#��h��IlR3$�I)�,% ���}�9��<�$�}⢣��I��b�����ΙJv;DѮo������֦�?$'�#�;��b���� ��m�߁?LzN��=��@��V���7Ϟ���������Ԕ�I�	�#M���O�]?�Ӑ�U�Q���i���[#�jC"еk� +�˫Y~&���{��Ĳ���Eɧ�%�Mnѧ����(�;�{M�A�u�3��ȅau/w]�0:c��]t�	��`��p�-=ل�Pl&�	��V_y�!��2�3�9�03iR�L��ΖZ)9�;�N�#�$���V�<�`�1ٲQ��K�a�F&fRR6"&'êLV��{��=��^����>�� �>HP��g������Z`��~:�ZI0� �kP�w�9s����ǩ�WX�֍$7�F�4R�1��i�n#�܈b�������-��˗�����b�L�����Q��)�'���BCf,�}��z�������)���l�������R	`�Ʊ�-�v��{�vi�]�b�_%���$���"��n��T��l�l����󟟘����n0P*S���Y��ʩR� ��8{-��#��II��1x�Ν;���/�L�e&՗b?��CO>�$�6�f7��d���9tH1>�x�E0� K��$�)��ڳ�"�2M��)ٕ��K���AI���?$���>��>���%�Z�|'V�����T5<6���OHQ,H5�Y�ec�"��7sAZC�*�3�, ��7+++��K�櫯�*ݳ�M�@�'O�<}��0���@�R�m%��q�|f\o߀�&6��b�r��B֢#o���K}�����Ǩ�{�e/���`_���I���O��s�-4��P�#4�)��k���'��.M�DLr&�ٚ�[P�	DI��:mp�l�KKK���0s��έ�sҡ��cl�͑#GΟ?O�B�^I^I�NX�=�Lj�a�2��0��R"�����a�]�|�u��d_T��8�J@��zO�~�7�~�`3w����A�v���p�#)�ס.//_�pA��������kh�d����Ȱ���4JZ�X�v����lnn�l0O�^P*�g�y~�\�N
�ٖv�;�:9ZL������Ӑ��LVDc��\���#���ӖjAQi��A��S�0#�I�o��`��z�]w{���>�t���$uE%lOTI�2�i~���9� &>0`M�K��>ѣ�uvfWL�ބ"�� ����ד���O�:�=�ݯ|�+��{�'�e��ĵ935-�.�&�� �<U��T�p����1F,ٸ�TV���p\ݞ4���0%.�fq�Ky�7�}�&KO�P����Q��Gswu��6��i �bғ9��&_!�.��s�mk��r�]"�U��W�ܛ9��s5��A��=�i����i��\��S�ڋw�v�Uom�o;vΰ�w���ζTP��O��(
.��h��faa�7���^)S���g?��?��?���V�Ȟ�N:;;�S@AA�HDԍ�����T�!ӆp�/���g�q��]J�x�X�]������yn#O7l2�<�.A��P$ҦϚhn��:o�9��{v��/+���}_���,�#z�1��m�mc~	�1A�ffR�M����%!�v�$fffpdph@��)�BAMi��7��߹u�@�p�IŎ	ACz~�ah8�Ye�\�"xgϞ�g?��ψE���"�n��h��,ʼ�R���^3� �Ľ��y��Q&(yG��iֿZ�����^�!��|ڛ�d>O~nz?�IL�,��{���Gή�?�Iއ���Z�Xb8�k;n6RO���Px���۷1�P3�q�v(;�����$�6k{gS���ea������{��Ξ��4]�?)&�����y�.Z�n�ˋ��XqG+�m��Iʏ�ɤ4�Qș��Q�l$�b	�WTή��C�V��EX^�)���o5�'��8&��������o�����@���+�i���s$f�.L'���㐙�*��۳�&H)�Dk @�� ��T���~�;��ZZI@	Ab��k_�ڹs�SMt떓m�����O��o��o���LbKh���h#��0ݳ�)8zDr�N	n��*.��x�������c�S`���~�0��YfkzW: R��~m����p_������Ԫ�ޟ��j��$�Zbr�5�q7�J�e��1̬�3���p`�L��-����,��248�	���j�-�j���-�I�Zrr;�C�˛���������뿾r�
�t7�A��i;t
;�l=�|m���d�8)� ��qg`�T�/����۱i�O��I3e�:&N�����\���Os%8���g��q�$.�����<��i5s"K��z���1G_#b��5�7�$V��T�zn��Ϧ��	���566��/=���(p��:�.�����C椠)�J@����N���/�077���rs�ƍ�+#V2�ɩwH��/
��y�P�� �=ƞ���������D��{�y�)ߏ�U�J�J��C϶�ɫ3�Y����������O�W������o�'�L�6tQ)Lc��u1��^�B�Y�j���?�裏�ʯ$T����q������@�$�!�����cG���z��K/�$��!�آSI.�9ÈřV��=�z��W����{��յ�@ QV��W�k��.�&7zeys��h_�1����%7{�Ȉ��J���SN2Ӧ�S�uy��&.���9u�Z`��fsL�a�"doV�T����������%-bX.�(G,4�&����Y���qۦmB,��$�(�:4u���| �iii��ݻ@� Ŗi'��-[cc�$�d,T�&����;�}f���6$�Co��#��=��w�|mUj�T"V��O�H�_�/(���u�ya�GJr+�w�{�0�M�}�oG�DN/{��z���;�Z�����*���f��e�[1W~L�?���ò�l*������*���    IEND�B`�PK
     uK\_����<  �<  /   images/1a257b89-3953-41e9-990a-6c271080df8c.png�PNG

   IHDR   d   Z   ��d�  �iCCPICC Profile  x���=H�@�_S��;Hq�P��"��
E�j�VL.��&I����Zp�c���⬫�� ~��N�.R���B�P���~����{�2Ӭ��鶙J��LvU�A�!�Q�YƜ$%�q|���׻(���F�����c�0m��M��ObEY%>'�0�ď\W<~�\pY��!3��'��6VژM�x�8�j:��U�[��r�5��_��+�\�9��	"TQB6���XH�~��?��%r)�*��ch�]?�����OMzI�8���8c@`h����q'����[�J��$���"G��6pq�Ҕ=�r~2dSv%?M!���蛲��-л����������7��!0^�����i���3��~ �r���_   	pHYs  �  ��+  ;IDATx��}�]�u����yoz��`PI A �.��1�eJ��bǎ��ɟ�CV�%"[+J�8K"Eɖ,S	�A �2 ��2�ϼ~k~{�s�� ��r��{��g����}�(�k�o�����ɓ'�=z{薦醮�ZǑ���D�i~�MW��=�9��"|X���/{�?���ht��5��.�֗V����0MӲ,�@a� _�߫���W���k4Hנi��1CS��M�hllܼy�O<��ߏ����~p�ӿ���?{�\�Z�LK�u��0y���3XX�%����<p����?����<�ɻ�g��j+&�$�岕����OX���5`ɬ���-	��"��pq��H�N7��Y��y��9��������r#׻r����G�n޲L;��R�R��� \�7��fL�9��*����٫_�QW)��K���h��}Q�D<%]ð~5�"x�=�����4�^��24�T�2q� ���|E\��J3<<���W~饗��5;7�����9�Y\(z^���$CͰ�4��͍�M(�ʸ�D^F"�)ub�K��2E�|o�)��2����h",%�,���A�c��1�c�_BǵbSw���1��c�^���~�T.J�nZ��L�V���'?���طo���3��tJ��ĚaA7i :Fh�r@1V�����Vh�~b@d�����bb�q���.�����İ:��:���sQU���������2c�dH+��e�"T_>6L]�����8+q�Qss�۷m۲q��Mن\��Ju~~~hp�ܹ�[7�@d!T+�lۙ���կ~��CYs�XZ���4� 2xJ�8j��1J�c��4��k��p��fV���P�m[�;� =�lۖ7L��4�gcM"r�&9o,�M��rCw鹡̝5��A5���c�����t6�9.�?�-:�v��^x���{2)W�{����m޺g���>;���'GG�� �b^�|�ĉ����{$�[�/�oӰ������X������_ӳnt|3�������k����Y�4�2�������1�e��t:}��y���!��۷o��F�ȝ�.|��|����@��i��?i���橩)?H5Y#�@X�(
HO-����(�0%�=��m����_���h�ihh� Y�H�+nʶ�o|��t�㏏�X,-�����=V�$�]�yQ�M�x��X\\��n�r��٧�{�o~�c��!��yƘN�a���ǲ1t(mSSS.�/
ܷ^�ֻ��~rz��ߺm۵��R�TW[{�P�LJ�J*�moo�~m7n���!ײ� ��u]�!�r<��Q��6l���+��������q��!#	
�|����k��O��g?�����tډ�����{�ukza׭--�r��.�9ʤ��H��g��������E\ڏ�X�^"A=lX�(ſ@������?�R�k��6�����mY�o��ʯ��L6��3O���7�� 
{��Oڵj��/��U��^�n��_��b���w~766���ݸ0����u�V8Է���g�B:33�/^��^�����Rwn�9u���ݻ�Z�.]�������׿��f�|���������ؚ����_�j^6�=����ۻw��mW�^���On�6$I �!���olٴ1�--��eC��-��a��-�-$�(:��CC7�8���y0y�΂TI�$x�2�B�g���Zn�y�gS���k�&&'��2����C*��44�x𡎎��Μ9���0��X�951տn�����'���u�?��s�w�q�Z�tuz�Э�7;��ڱc��Y,Q�M�;رf͚��7�<�{txx߾�����?�,���rНt.���7�|��ҙtgg��Ǐv>��c�>z�֖֭�t*��㏟8�������D�����||?t�)�l[��a�M��lX�`����gϣ�/^����8�rQ>(�`�@.\�|��41Ё�����υ��Ν�=Wks��=�~�kom{�������.��mmmE&�nĔ�Y�U��]�z��i� ۴j�*ֳR���~��_-��_�t��c� #���ffg*�i٘OGg<`�R.����ɉI��"�5�M�G��<Ũ8vk�·[�]�100��
�N ��63�l�P������ݪ�&h����2bxhP:r���� � �a!&k����}��1���x��������׿ޱcdppֱk�.��7���ڵk1��}_�:��[o=��#�Dp���@�333���������Y�>5}��1�h:.��ٳ��h�1�1��uuu�=s����p��ɉsg������Ĭ3g�f2H���u��T��S ̊<�n$���h�	��X�E���hoߺ��2��
�H�����_|��0�ڭ[�~�����������d��[o��������l�ΧG?9z
��d�X~g��ǟ|"�S8�ώ��c���ؘ �R���o`����
���/���
���	�'2Y�h�G}�'�c�pdXz`n�Y^�tٱM�KbW�Z��\�$�P~JAY��鳖����.�}��X��Ҍ	���o�)��9DQ$�9���L����'�F��G�v깎��Pe�3�r,1�� �:~,	�˟�l�QC��������\�����<'��(�#�A��e0I�e;�LI-4����I)��r9ܢ����0r��-,�h�$��<=K$N&Eo�4lJ��) 7i�f�s1*�L�\A<0ܕ'�'��I��!�J�aA�u�(l�����Z�E0$���Iy[d[F�W�kC<�$�k��⸞jՇ�8^3v��5���&a!�I���$��u�Kd'�r��|�ҥK?�REZo]�V�MOM���׈�W6�Q:#̄�Y.)-ɇEI�b�Y��]c���룅uݸ�أ�U˕\�Q��8ɫ�vPW�	.�G����L�RZ�lbj��`/�U����S�a1�>�]%���ز9���O��:)�R���e$��Aj��B�K*O�`4N�^�19>o����k�^���:"�r�222���Dv"���.�|S�Ԑ�/'��d��hEP)�z#�$.
4M}�x)�.��YZf���!=9+���@���K�KF^�e�+���e�W|�S���AD��׮���+$@�j�V|�aHn�)�G���Ct����,� +Y�%�&��Z(�vHI6����k���Srh�$����2m�]`�������K��;Fo�z�����~=�,�����c���0U^
	(l�Q�R���lܸ��&�l�?!�G��#NBv���3gNW+�z~n%q�M�K66��.��vm�5��FS14�s*mo۱�e�7�F�� US�P,��	%(� ��X��QF]��+h�������Щ�5��R�t�N$2��,��o�������hk�5�u�\���UAR��λ���[0	��l7��8Z,�1�"/I"�D�����z�/�~�;Z-�)c���+�.�v�k�C����g}/�N���;��"$d]%�B��eD����������5m޼�7�Dbhk���ً��F����R�%G���<�&�9H��J�B?���~��{t��{�(���$<Wu��5H��/����z��f���B�����Ka��LtߗJ�>��ã�}���^���A�������5��S-ŌV�X��}m���L�uR�s�Tj>�4����B7�v3錛Ѳ�b4337S)zސ�v��&dŶa�����יɂ��2.紡�kbb��M�����B���XΞ��<~�أ��޲y��8�ME��ԅ&9��@��N���EA�Z����ؖ�\oܸ��G��#~.�V�u=��!7���� #�Z��`v�2�5M7<�ʠ$�ߵ��{<X�hnì�5&S) �~X������گ�т�O�A0�Ԉ��O���?9�!6)��I��!	N��m���� �Q� .��xjr�\.�??��5�R�	3Cr�H6a���C�&e���&ͲȱF���7n<|�=|�����;��������T,`K ߐL#��BP*�E?��}�R ^ӨV��ٙI������+Ր� ����C��0�j%Р$��,�n�-�+�rհ��� � L�h4�8��%�K<t���?#�KYL�&���EhN���/,Ug`Dѷ�*�DP��\�E��+W����������������0��U�i*�� @�{�x�vy�08xZ�Ӄ�jvqn�ڕ��/lڸ������Ч�2K^e��h���eGNʁ�u�dt�ڤ�,I�W!Z�T�1��bc��ƅ�z|LP�Vg�q|���������:�R�T��dD��"� �z�l �����T������B!�J�;w����5�F�	פ *O4C��F hkZ���O���v��C�M͡�Z��'�;��[.mz`s�a�B�tB+�"H?����9eщ�u,�.V���}�0=|S��_����R�uS��$dQQ�8VI�KQ��m"� w��3!#%�S�R1j�5�Pq�D� C/�>����������pd`��+�/���*6%;�XK��P�jt�����^y����.�Z���v�nGzˡ=mUm�Թ���Ɏ�6U{�z]L�	aѵ�CnT|��9�fX�o�H�\��]{�lْ�6`+�������&'g�g�BKf"5D�e�^f��T:09bJ)�ч��4�@��ٚ�ҚX�E�f�"����]��p0|���c!k~~~rb��}c���R.���c�L�7Ym��}a���W��Z�5͖�\S{.rW�zI���7�Wu��B�����\>�=$��H>56��TQ� >l;棏�پ}��X(�:�E�'��
إ\bML/T��ɔ3��㤡X�j����f�|��>���L^�T�!���?�~�zgg'��/��7��6q����%/.���nٱ�9
e�l�����7o�-֊�E�v[���k�h��r9�ՠ͍/VK^�I����_�#�'#���S4Y�u�m0��Jq<44��ohh�y,��삁�K�4M��r���beaǘ��ӯ �T�p8p�ˎ�� 𽈩]�8;;{��1�&�����"�Z�r���?���K�1x㭷~i(&��'ѐ�rfkIy��c���ڊ�rSs���)�ŀR�R�ɘ7;V����j���Ԝ�j�1� U�f�@Kj������qJLLMpc�z[{����QT,�����&����J��?��%:�J�S�j9�RSS��իWc&� AX<��a�@�J��0?_*�H��Ru&����-x�fg�M�Fԡ��B��b`|�1Y�c,E�ZZ�jmG��U#��(���3>37GqۦhG&��43cHݑ~W�L[�+�Z.%�)׮Y����),��(uU+�T���!�@��lq����&O
�_C���3)CU�CY*�f�w��(���~�駼�!��'�<y�d),�4<�f��DhH	�4R�"�޶�=kg�Z�F�մ��!�ٙ+�/�i�X\ܰ����c�Hs8d���@'~��MN�|��C%-gfz��_�juO��`)a�Un-��R�t��G<��ÎN�>�������lvv敗_Y�fM�\;~�����ƍ�s�;�v]X%��-x��(Ѐ �|1-�k�����;��6R
x�L6��}z�9W�X����������V�Ѹ&��ZPmliJ�ٱF��R���9<<ԼL�-U�q�gC���-Ⴞd�@@�0S%)���\?�*=D�Ӫ���n����$oݺ53=��&9� ,|Ӧ��sCC7��y��3�<C[۷�7�8w�������L���SF�S  �0�k�A�
�'ֱ�O@KpS�ςf��e-7�T�r�{��<��(�WG@��1��ry^�5�����i�v�\�M��ת�lCn�i�q�\��������GÔ�r�z�A��08Lu(�OO"6��4�02��7qd���Y(��-?�٩S_�^ݷ{��|)��M��o���'�LO�ܹs�]8��Jцr��C����Z7m���іI��mM��>���Z���_��Ad}k�8_M8O��1+�X��~���V1��Y�xAWW�J�w�z���ۺ6<�!0�����S25;�j�w�UH�B)`$�2�f���T���{{��a��t:����K
��#�,��_���|N�\xz�ӣ�2�2˪�u$aHE�]hS6��88�,�|*UQ�������@1H���(�I#ɀ��;-�t���|�pR尒io@�E�o�[۔B�W�ʂ�p;�/1��4i�Y�r��Sk �� F��+x�B�R(aU)
c�
ȁ�uwwe�����������!+1�V�)�+鑐�p�Xq;<L�\�\�v}fv�����)�$M>��j*~�hM�*�P���M��3���^.Z!dD�V���Ժ��9�gcH�DE��DF�&��m�`1E[c%;\(�<"�����3H##[[[1E�tt�������ө�)�Ϸ�z�.>�̙3��J=z��j�A�Sh�fJ����mOX���yn��zz�H��L�s*�fK}�� (��I*N���a�S8�@���L�>�I�B��b8U�$��|=�U[jB]� 8�Ď4?���m-��ժw�����q�9*����;�G�ñ�o�m������	�>��{���kk �vPMn%��v'�������-MQ��%H���M�4I?��q,�n�+h�~�VҔE��ߦ�Z@3Д511}g�v�3����a��I#a�p�jz��P��I��w5ɺ`�.���K��V�!y����	+N�������R�\��F�92+AOp�Ҩ��ը��qq&����eT��������/��"�<~�~��?D��F2d�&qfL��*S���IfD�m�M�nδ���|�r%����Y���{��H��T��Y�Y-j?�l$�1D�T6�VNmQ���Ȩ����V��Zkk۵k78�S��>�'�t�<��uN{���[���0�yj��mYUf�I�Ї�hq�
�j���4 ��^{��~�K̠Z�A�1G�X��F�����~%�4fj=��×G[R]ٮ�r�������_������sG>�o��}���[�F�;-n����=�� /�0(�kOw_wO��t*�U}�J?~��:w-謹�Lj����+&���U[��R����f�P�&�a�rs���E.�0�>;3��d���~ծ���L*
z ��m[��ۛ���Ɗ�������tƁ���״���h��ؑ��l�jJ�;T��Mv��iKݺTE!��X'��xf[����M�[�o����óӳ�b�����Au^� 3&�J��tؐ�A6�rY��jn����3�^� 0h���a\G��b,e��j��%�U�_�����7^|�e\���;|�A����Žp�
�I�+� ��>�13��F��v�l�a~n��XnL5?���~�������uS�"���@EI�,���nTK����=%�9�	�s�![,���[���E�Ɓ���᷿�Y�z��mss�v�u��KW�\{���p)��;Ｓ~�z88��m���t��K3$����_r��RGQyǃ;�Tj��{7nݜ���}R�+J�`�n\�XBJ�G9�_�UJeF
Vۣ͌ё�޾�6��0<2ֈl��o�������rbh�?R����(����r����7�֙�w�t�9?p����D���z`z‚��7oْ~������z�M��}���ᑾի�y������< �#m�B��)ff��j�J�)�1�F֝�j�ֶV�������C�>|�T*A3���7:�3�Xx�j��͛�ǘ�Փ(o0l�|�3˕ڢ�Kw�R�Iobvb�s�Ss� 4�����d9Lz]�h9]��!�@��@<��6�,�:�!}�L4`5J��N1ma���%?k�?x����ĥK�&'�?��c\I5�Q����е�G�u�!�y�枞���6$�)ׅ�Z�ei�t}pppqq�f߾}�l&fBN�:�Fκc��RĈk[i��u {���-��J)��L�����Ld��RwM\����&��}`�L��'��:qM��0�J XD.r��i! ���D��z��{��]�ߏ�yuߚ��XW6��^@<�ia�D'{Z�C�f�iH�--[�lA�PI30����ٱ�1\ƌ�hmlt��J�����;w6��iġ��B3"0WEN�Q����Z� iom�)��ygG�MQ�Tep=Q�)��eS��69
�Ҳ!�����F��"(l "D����$�j9�`"?���<}���{�Сo}�[)Ӻt��+W_z�~�X,�GS���^�o��	iT�G�NON��5C�|������m��ZZZ0��Ǐ^��$CӠ���<����aF�nA!���
;��r�҄���B�����2S��ѿoS*�cΐ�`�F&���; ����)�Fj,L�S�@O�� ����{1eWY��_�������Tz�����mgrrZ?33�Jky�+hD&6	s0xƊ�Ł��CJ�)y����k�Pk7��Է�������g�֛�X���P0v!��I:7\�ˇ^X�]��}zqR/MvvuVSǚ�6m�ޣ��wLI59b�5C�r�l$;���lV$,`�7>��#��=�Z��������O\���%����r!V����k�t�����_Г���������P�3;�b�F=���F�_��������P���UpR���O��
@��C����<�C�`����NX��F%(f���V�˺��ۖ�צ+38�����9�ŬE���H '+d� E���j����TNY"�#{vَյ�#�Zݺz�n)���.N��4|B7Q�σ��`�gg��9�u(�͛��ķ��<$}ۤ>T�M�Z�P�Ϻ9tb����o����&f$�?'�\��
�s4�3"�ٲ�C�#��8�X��3�7���^��4ڡY�U� ���Jdl�����siN\`qݥ�_�q�z��Z��sc�A�)�nr�K��̕��vK&[�b�2�j����iv]�y]X|�c�"���^jnv���4�ff��śӳ3�VD�Im2IrcCr�M1'eK&�k��b�h��F����ʘ�ִ
��1H)�L��ԓ�q+��^�|�6�L.=?=�!�blt��m�Z�1����=�qg���{%6��3]b1�"Q*��K���]�W5���%��M�(0V�p�(5Y'����j���W-Uʲ�z�t�h	��w5�<U�l�$j=�P��q����ZL����H�Dhƃ�UYV@[^&U�R�2g�g�l�з�׫UlW�T��;Sa8���ű-����8��@D���!�	��w��M�L�s�t:�[4ds��Hnm4D=��>}�P\�l'�6o�g6�q�ͣ������$i:�BX��Py��Wa�8��n�$�0�3d�%�׏����W�.y�k1r��,ҽ�mŵ� �"�·��~���];w:��	H5==}���'�x�c�; ;���^�v������;����E��'��\��%�$j5ߢ�HH�h��6�MNMpa=@�1-cr�N���'���X"r�, 	�����P����Ξ�����;z:��_�B�?� R���'�n5����𭛡W6�Ȍ���ry��XNM�$��IF1p�Ν;?x�7��\�v-������۷/�- �~��G�=�ܦM�\*�V�n*��P����h>�I����rY�2�	WnE��Gl}�����C��|������Y��R�O��z���O�fTfkY������b�T�������Ե�3ЊB�Kg�j���b��'��"s�2'��c�S967c�B^/$ �{�iCf�����n���ٙ���|߀�
�o��H9�2H�/��&�&����{˖M��EZ[�C��0/����<���gΞ�	�8�>����o���q�$a1�I�/0,.�GR��.f��3��>t�Q6w=�7����je,�d�֦�'�d��.;6cr������C"��*%�6���↰$.�&��)W����"ٷN�ab@F�n���Ȟ���#��=6l�x
j����[��T
ŗ�ݩ������ׇ0M�E^:K��|�Q�������غ��c��a�H=SL�RuUg2�G����ΞY���"��654C��T�2Ҁ]}�)mt�ą'_}�3�[D�qw�t/K�^��S���-:�g�W��3/�XX��H�k��g6�6Gx���\�t9�ϗ
��n���׷n��� I�Ν�� ��KE-Ty��J�48xi&�?��%�u||���_����xߚ5��PW����x����ౝ��l��H���KG��Ɋ�#�@���窆_��ܾ���3p����|cO���fE���u���Ϣ�SN�\��[����U���/\�1;[��}>�"���%�ï.|��5T*�(~����$���	�8i��ٚ�}��A�j���+���|�X�U����������.���_1�s�����*U�{��b ���i-��Q�K�	1�9@(�X+�^U[ӷʴlD��\S:=��ݵ�՚����ܙ�����뺄4CW}���J_�
u����bajv��&'�f3�,e`Î�Dgn(�����i#�n���1;��UA���!����t:��6�c8A*�j��ICLaHg�@p�b	�	$N�Q��ٹ����|��ѣ7�ݨK���Ƹ���Q}P��Pnß"U
��QGg{���f.ʶ��Lz���s�b�*�g��XGj�SB��-J%Ȟ��|ֲ�/"��mln���Uʜ�ػv�z�f�T14��pj��E̺�-Y1�!��4\p��_o�/B���ԈH
�CG����C�,r�X��ȑ;v������~~��I:�&�C".p��c��O����&�/[��m}k�u3��yay~�|��P���V���K�k�W��I�F��TZ1�;;ܱ�S��l��u QH
�a�T�d�8�/V�4]����JVj�F�舞�b��1���tt�a s��+.t�x�%�ʫ��z�Сcǎ�47�����/�$�b��R3�t�Q�f��9��_D#*������|�r+�R�L���ic�֎O~���5�������
��Z���L}����%b���C7o���7C� ��H��<\X,j	��˫�*��e�ݵۄ��h���*�������d>߀tU��q�Z%�<M �=3��₈��m#{$�JHdSKg3�w�)EeU�� �t֪6UF�{�}f�M�M�ՠf��C/=z������3�<k�6�І�C�/m�WNF��'rgr05=}������������r�O��6WQ��:�����Rx�
K������aA��Z�L����dG��O�$MCX}`۶ ����a�֭�2�ei�l
�H+�l�����k*>�6� ��v��̍�LOn��`��O��l��rg?�|�����n�__�P�%�Q�!�q�!��k8���N��:0���؏~��L�i̧kU�R���;N��)%�ԡ7��W���JUk�~�&5�1R�U
L%5��X��O�j�M�|�q����_rlÿ�w��um]V�&q�R����{�����t7�9U����s���NCs6�����P�/��ǟ|���[����C�q�J�� ԓN��P�g��Y։)�(���4=�!�7��Jc�׹�d۪���pچh�O�_��K�J,u?�5�l��AB�ɖ������!FhǕg�J��B��K�b�\E�7����O�}ǵ[[ښr9d�%oZ�{��N��H�����*�
w�"�\�2�����4 ̲���	Z/�]�L�[�y�	E�f��2��&E=^����]S%�5�3��7D���=S��8�WT�<��Ry��}��?ܵ{7�V�����34��'�rټ������A*�jp'��Li��(������I�n�E�����a@�Q�m�0ݼi�-=�Rs�s3�sݩ^e�[�Ff(4-�9�G3�׌]��-hR�&Bi~��P��E�B�T���3��0��r��Tb��!�T�k�_ᇟ��)�
b��Q]�����g���������LPˤMON�~��ڱ�{��F�p�x���ySU���T+�v�zi{ժ�æ����ӯ���j�~#M8a>zk9թ������I!̎��}$Ky[:>�4.b�s�-Mk��mܸ/...NOOMNN�˥��B��M�uU��̎�I��I"H��Yߏx�9j� ̾i��W� ��lc6��V�u�r�USw�}�Lm�FiW���f��$Ir�w������r�ܘjٹ��൬���1�q�!U�"ً~��g�}�}p��G���7��p%��ؾ=/��Boo700z@�Yonn�u�Ν/��rllp!V�T	�(�J�y��J��TB�}z�ض��wuPE�7�z�����E�5n<��$���"�lpd� ��W����«�)���7�ܾs�NȊ�Ós��ۧ�D����\�_KJ���?���i[�ɟ|{��}�A5�����p5�r܀��nݼc��w�}���.R�`�v�Q��l�SE	�{/�3���kׯ]�t�pL�Q߽I!{�t�:��6M&*^�*"�E�u~��V����`��>z��;����$��3���-��W�dS�0�3�L�?�ޞ={J�bcc���\��f����ɩI`�?��?��x�b�
b�0��t"���zzM�
wK6K�I�H������1��n�KV�X�	�iO�)bfy��iڒq����~�v��i�~2������G�i�������]��Wuu57�\�BD�8��{Զ��������'�'&&���sKYR�P����FUc.��pϟЛ�xI��Sgh(6]���BB;=���p!3�N�ɺ��Û$%I�U�O���n�_"�e��4�i;������O"ά�[�o��2!1�\�Lv�A�{{zrbݻw�����
�"o�����Jx�x$�*Vǥ�4Z[J�5�9,s

+�\��$eeM陪���#l����[�B�V���']����?�ǚȎ2m�]���l��3��|E����Q��i[[����_�v�D]p|<�R��GZ��*YLCD)�<А_U�'�u����������F��&�-��^G������?#/�{p�t&�zu�qss���})�Z��P��&�|>���;��nݾ���Hғ�jK�R�2B�&p/T�u�R�"K7�R�"Z~�$�P g��nߋ�:�,�R�k�)����T�70b��\O%\���X�ͫt�(u56��Z���Ը�F��M>=Qv�p�G�h�d.�v�#J�,��:�*�����eۄ��%�JR���S���ꂸKRwI���L�
w�	
�KAG�%�k�c�ߨ��dԢJ֖e7��Ӗ����~4F���T��7�e*^)���^���+���
�v���}�.�5is�uEKI!�0���w��8��S.��M�+$j��5�+K�b�T���D
��H��=����No���h�����b�d���m�ۣn� pl7N&�<$)^������姦��9���o�	/�WN[�����ݟ�%M�a��9�s��rμ�*K��=0U9dЩ\�����VH�<HG͖Jccc�t�_:��~�	BQr7�mu�1.���[e���r�V\w���)�NF�t�Kż{���+=Կ7$Rf�C��]��⥆�{󴙂6��	[I �'jy����őё�ׯ���⎫V��RX��!]d*�*�dl/#O���&
�w�JJ��������KW���	_Y��9ᗔkvv�������,���U�r��i����09912<��Z��ݻw/u�V�%�|�-��c�#-���Hr��	F_[����J+�{�=����c����=H�$�t�
!���_]���߾���|�����f&?-����&�Щ�W�\�pfaGG�SO=E{V��'�X5K�C�!�J,�#��izr�[qݥ�m�qw��ǻq]�#�U��^�n"�$���zrެ-	w�JՍ�С�t���٧ǠSO?�t����mY�|�G>ѓQ46>v�칳g�^�:�oA����ʆL����Ul�1hk�O\��.wq�t�g� J�d8�N��*�յC�c�k	�n�F�T�:H,�+0?
ܩ7�q��(щb*!Ɔ� �k&;�'�h�o��G><27=��}|RKf~q&U�VXR��.]�422\*U Ξ|�W_}U�em޼y��-�??a�9�����VD>�N���$� -ӑ�7��Qtu`��>�&��93���Iw�n���X�)=Y����?ر�k�ƧQ����e��_=a˄~��~��jd@==Ȅ�-�ren~vzzzx�6�B�$�ɾ�������@�1w�C	s��?��������]7M�a���CUz+����ҕ."��q&뫮��eN<V��C�$�ֽrbz|�z��n���d���Wr��ęPٕ�$���K5��a#:��ƍ�B7GA�{y;�m۶�׾{`��T*Sg������������߽���o��d�N2��=�H<I\7M3�ɯ ��4��t).�M�K��%�$�b=�:� ���\�V�������[��iݍN����r�+���gh|��rt�N�����[�������0���<5�����������?�^����I��iZ���jIJ�2�՗��j���B��]�"l2C]"93.9�]W~>ɏ��K�p]��{ÀZM9�[�o�)&�n�A+k���Ԙ_��r���lkk�Z���"���+^��Lk��    IEND�B`�PK
     uK\G�BN��  ��  /   images/d6a4f4f6-fe0f-43ac-893b-20774d3ea628.png�PNG

   IHDR  �  �   ��V   	pHYs  �  ��+  �kIDATx��y�$�u'�""���>��{fx��b-Y�����a�`i���\@�DYkѠ z�����V^HkJ� H�]`h�0�W�6 ��C���Q]U]]���gD���}/���̬��:�*���de��E������"�(��":$�@%��"�(�C�T"�(��":4�@%��"�(�C�T"�(��":4�@%��"�(�C�T"�(��":4�@%��"�(�C�T"�(��":4�@%��"�(�C�T"�(��":4�@������o����O��I\Ҏ��qU_,���i˲�m�����xH>~������=��O�O�ж�ե�N(�wܦN������s�q��}��񼼞�s]�ZW�V�q$	�I^s��帵Z�q�:�o:.�F��s���%��4}/���=�JхY��~���\���z8F�R�x�������>^ﻳ���$�I�����~�K_��Ʋ����?���v|VH����#��y(�.�o�۱�����#�F�s��~��f�����s� &iAF8��k O##���S!��[��c��od����u����<�;��[����>�.�Ԉ����j���6�NL� ����է���^<�c�b[�����4F:�Mc��e_9�ո�&������1��}����ƍ��>+x/�u�F�[������A��������>�'�������K��V����/��F���1�{z[�����>�g��Ó�m��apoD�	�i�����M
r�����K�1��L�-�J.��࠻��L�����	t	h�=0XF�zx�J�[o��|�k_�×f_�׿�կ~<��_�k�����G���b  �o��	"&��=La�0�ݶ�]A�-Ҡ�d�08u�����i�}���g��;�p�A�։�c�@R%P�@�̙���ϒ�@oτ�A�yԘ(i�8�z������t<�S�<0܎��E+�?��b �h�n�$�h�.�g��2�{�����p?��_���K����_����iP���6t�s���|�3�5}K�{�O�Eǣ���.��l�E�����r��O�����i7�E�rB��o�&��\��7��w��{��O���#Р��>MF$��iG���a�e�Pj�M����V�����o�䘝��s�Ob�)xz�{�`�;�~׸�������Ӹ[�A��K2{��� �E�������6��旾��%Ԧ}��x��������)�2�D�r�t����ſ����Y�x�s�N~
��DP
"����^
�'k��+tԒ���on�j?�7S���w:N�<�Ƣ�����|�h��e�/J��r'�ogރ��I�uaS�~��c��A�o�i�q����!�GZd���H�^ZP0�����6.�}����'?��!�<�e��?�BQ*�D�'��_��k�����q�M�lll��$�5�h���N晈�^3:jM�5;�Nb,�x��|����?zw��p�����ߧwA��������P��k��&��.� E�r�D�����~�7~��'��L����Ĥ�H@"�MF�V�m;3A'G|/�~��Q���a��^����7��tþ��"�M��������>�D*��	u{{�[.�B�y����6�a�@���W_��������
N��kkk�$<(�U��Z���d�
z�����$��q��ڝ�����;ij4�i�����}kk�B�GL~�WVV��ŋ���ۻw�V�R*G@d�����w�ϯ�&��Ģ	F B����s��9ġ�ktԚ�I���:����z~���k�اwY���B�z�\�b�H����7x�����W���۷o���T�^����?����������7A�W2q��8��g"��If��i%�A�e�o��P�"��ä�B���� B�0��b��w]�����Ƨ^y�������gƎ��!N(����7J�җp���(�τ�C�9
���N��h'������IK�'M�=��D��"1y���wz�i!�	��O%�����/��g�����w\��[�n���T�(L��ŋ���Cu����M�Lr�K(a�|'��$�(߉"p�^�O�&�n��5�!P����Wj��廄O �R����򗫫���ڵk��͛7�)�T^�._�ܷ����P;����g��v"H���mE�	%v�N�w���i<����4V-�{�'�%mJ^�|����Z_*�`{{
��� ����������>��ϹpJ)�� ���	�CCC_\__��BD��%N��I|;.0	[+i,|�/k�;L���c	_�0��M�4��A���Q+D8��]���n���V�t��v~Ӵmj4Rs���N�d`A��t:�_�����������2�B�@���'.\�J�5���&��HC�O�(�yڵ�V��&��y��Q3���$�J���jx�vRl����ک�c�H����	x�c��aM�y�i����z'>���ς@tyll���t���{���S����s�OMM��|>�8�.���p�	�OL�%!�4����P��:���'M��.�tP-�/ʀ;��	�0��� ����Κy��uH�;�&*�2�[�  �<��&���l� ��677���������]�z��O[����x'D���_���rrr�_��>�(,����
(�� �@�Njl�}�:f�x'��e��i������h-�V1��P�J�1��mu�vc��Q�����c���nLOOuii)���/N��-�w���hrkk�fgg�%�4IX��JȰ�j0�^��o��Z1�v/�i�1��#�:�����t���^�'�tV4�!�v��g;���Y��]@�������w;�����H���R��q��z����/O�D�r ���J#���������ؠ&��3�LмH&�Ld�tҵ�^�ZI���~��K��~�����yMI�M�L}����� �i.��B�yL�)�@s��v�֛۵닐��ȹ� ��Hcy�W�r���*
���4�X"Pه��旗���ŋ������4��R�D�Z^D�U5��N!�l���\�<�Uϳ�A���ǉ����ޯ_MXh�d�=���v�5�;��ZP��D8%�B��:�?_C`Y��7����_�AS*hvvv`}}���
J%�%q�@El�&S�I!aħEC�O��PX���:Q����l��E��<tڅ�n�NQ]a��=k%@��t���6�>��d	��^������t-f^	f�%���ꪕ���������CS*mU�����J�MRI���M[2���n�V��Ln[�A���d�'�-�u�V]��+[���1����yjޠ(��[�@���=��L-��z�q9��b�z5�gJ�g]c���^d~�����qĤf�F�� �p�@X��=��"���G�#����
�������0??�]J������ɵ����ʕ+��
���%��4z4�f:B[�7B���&��|���pH��}����$|/]O���ǑN��%W�W���àN�P@\������;6��:~+a,lb6I@��Z��ׯ��;w��?o��ֿ�֬�TB�R�����/^�ǔ�(*�����ItҒb+iȔ�Z�0��ޛ�M���uwY�w�1��eN����k~�-K}wA�L��@C�N���p+`� ��𘸽 ��ы�A@�]�� =w	�i,a��y�N | Qatlr��_��_����f��)�(lxaa�]�p������B�Ib��c�����vS�
k"as��=<��IȊ�H!���w��l���Qp������l4��TE�L:�G��&C��*CD�A�4	�����>�V���|��Tf�WFFF>=??�����~��U�2�@Eӛo�i�����ߛ���
}���M��0������"`!O��E��Y%W�B\@T�&W��J��/>�S	�N�?�M���򼶴�uH~�j�u�u��<_��) �4�����<�~7�M�,��9��O��(M��<�/�����
�IS-	룇+�}Xj<I2'z�H.	M4���ZK�}�ǎ�5�=L������VEsX��=*R+08k��03;;㣃�����uҜ�!�΍*Dt�t�(�p�~��D�lM�iu�����̏��G�����{W����2{���}�ʕ+?I��b:j�8i
�B8z��VZ���KQգy�#�$ax�\�|�A� Ǫ#ʠ_��������A>zV�
T�i�O�]}�QB��r���`y$�h_N������:Y	��2�knWf����{L�L����LOO�߸Y	��"PAZYYy�?�V3K���0dq�đ}\���p7��&�����؝���$�O����8�C�`�Ǫ*g)d�
�
�*\ٍ���l����t�Vf�H 8Z
�&�m��
GK��g~��%�"�*�������@�k6��I\7��AQσ
i)w���/���fɇB6m�2wu[R��(�.�m���y���E2����A�{,��LNN"����R*P���b�%��@���#�<p�)g;���X|�h=�W�P�݆zM�2w��x�M���*�+��+���&3�[̿GE�����������;�i������],��{cyyy"P�.3����R'IK	��%�~�VQ\������Z�2����G�lZ�}%F�٦�;z���:W�E��0�Vs��^���V���i
��V��|0A�G�������W�yP��
J��St�@f������^���":|�z����C����@b�Z�����z?����*�
.՚��b91�x���t^eI��M 2��V@a�f�;1���#z9jMf���!M�L`��+7n� {}ׄ�4����[��?���Ȉ-))��i�Y�)��.��ђ��7��� �jɒ��J+&�i���y,�vJl���9t�:n��
r�N$��i�oe�'j%���K��,"z>je>kU�!^Es#��\ĹA���t����N
�U�۴%�m��L����0�B���DP��*����J���y�����嬊����bqZ,{T����X�؆b�uO]x�M����>!�&��s\�Yfu�V"�Y9��.�����*�>/S ��r�(�dq���iP����#])� �F��F�P��Lf�����
��<~���RP��%�a�@%�갾�+O�̡ցnU��BP�i��|�~1$�gHҮl6�	#�w#n&v��x"z~:(X�S䙠P<�ϰW-A�PO�
>�������b�/�^w*�sXC�"-�ةe����5�y�&/;;�֗������N_�ӈ�|ۉ���,WY587�|.v�d*9���"�̤9�ANZ�w�s�$���"�2�^J@��D��������	���2\,����A%���L�Ӌ�U�L�S��&BV0GNR�Y����a��"�csS��l�0	TXC��'�W�%�0_��m���k��RY(
pnj��Y(c���� @�@���5X\\ds����\��Q�t.�ݘ��t}4~�O��HhkT%��頡�fJ�h����l����gA���f�+_��z���qZe������N��oD�PE��S�R�$Ι�gAيA=��*Iy�Xu�k�gUa/�j}� �	�Kk�<�&5$W�Tt�gY���x��H�!�� ���+��}C}���^I=���xI�?��%����9�Y[�����eT�*����9a3�5�*2�;e�,�j	�ݻ���/쀅��B�F�<-��=9����iօ#�c�}�څ�tE�Cς�����a|\�B���L��<^����i�搱�,����N������k�?ӷ�Cñ.D�-tLJ��c��b���U�����mO>���A E�H(����ļ�2�y�����{��Jx�Քu�h�=��I�����wI6�@Pς����8Jx���"NH"����p$�	����ɋ-�x6���?
-Җ�����EJ�I�k��0��Ǣ�q��=AK<f���`uy	�Mg`hbr�A��m|�)j�֙�x�rvJ۰�dޛ���˰�S�s#pxq(n�����!�?�|�G� A%�� �*�w���Çp���_Z��*��e���Lc�3��.���0�U?�?y��#P9IB)l����'ge7�K*�0�<N�L�V����8�]݌��n��Lil� �H����q�t�a2�����D�t�:��ѩ='���y��� /dꭹ���!5�+/.£G����	�y��{���0�ܺu���qD�u"�i�6q��]����B�j����&t�$������.V�ՄD�H�K��I��#�"P9Qb�i�k<.	V<�� q]+L���%�t��D-�*��'M�L��I7��)NA�>TJE�X���-H�`,���`��p�U�{�"�v��W��A̩r�~���j��0�t����N�Ⱦ���{���?��k�Pr� �P����X�+��%
�T$�K�%gQ8����֓�����dؾ��uc�Jؖ�
P¾�n7�2sT��J��*^`�����^ZSq]���$H��X]��=�NBN2�it�$���& �h,+��Z�����bbE��Ь)A�\��|aR`��&Z���G|yN:�r3�6x�4;r
W0�g@�lR�Թ���	����IP��(�/�%����D�������}?JD;�vm�N1Z��)N������}&�/B�o�ͬ�\�P����+ˋ�����B�z�:8IԆ��6��� :�kU�\�@�eֶ�0��L��@2�^L 1:9����@���+�uUY��l���?�	R�jX�s?|p��,@�N��(����߱)"��qxO4�z���{��Z����q]��S����N��Փ3��<��E�;,�w���TZ��z�'��'��2�aP}/ⷤ��e�,�'�GU^
j䶐Oj���l����a{}���۷o�/�v�k�x��i��r��_�T��V]��t�/��@L�Q����FԔvn[:ynp�������#�\�|IZ^^�qW*V�_(����ADGL�԰��|l������ߥ��=8a�IPA�q_�)]a�~wcH�9�Lm����ˊ �P)|�����H�Z�;�k�da�rYH%}��>�T V�:`���"�8�,ȤS�{���u�0F�;���g`jz����qO���y(�V�����,$�bq��-���*<y�`���L�ٿú
n�����$�RO�~�,��}�4<��#Cpq���C�Y}��ݻÎy���iԌb�l��1t�I���1#��Q�-Df�6�U$4�P���.���IP�ZG08�Ɂ~$v�Nf,������k~�%T$X�Td@�x�����P{��N���C��m�c�2��k0��f"OV�u��L5a�(�>}�����8��*�R|%���y�a���qnܦ����9��HH0�UA��\=7��v�R�ppp�*
#�5�zT�X���\a��� ����(:��۫�F��>�6�ޭ��N(	sc}�AE��*s�ع)�t��}
�s�_A̷	���0�.^�Үr�K6sQ��M�*#����*P�]�����LO�!ˠ��Y?	�2q!����]�Rd���A�4Y@����p��<x� �;%�$2���q|]eBG�y��yR�Y/~�t:=���6���'L=*_��W|3Rޤ���- �����((��b�5�dL�T�6�Y3&PU9���`A�;���y��2�t��-$���|�2k ���Sد�5$U�ǿI� ?i+��� ��)
�4����#-����'��"(V�|2}ј��dx�5�������Z�RL�Bϓ"qL��l�pȞ�?��?I$��ӑ���}�d:GͶ�uY�뫬ۦ�_j�=�m�!K�c�9���*�R�Taaa��M����L"����>;�T��wZ��#3��/���P/�a}�)��=���W�N�fE	�:^����G �G�eI�pG`|�<�JC�*���2<]|�k�P,נ�S�F;�n�Á��q���xGz����W#�K�Z�ַ�E�D#�zTr�\_�i��?Eb�	(�0��')O��+XNS�xIt=Us+WY���#�����u��%d�H���"���w���P��� ?F�s*�%�&CK�T�>�{�H+���GZ� j(SSSV)�_�$A
��@ޓh�u��{�8��/�xz*�I����%��/,�� ǌ���;v�G��#��Sm,U�E�穢�@`����;z��?.I_uas�Ž2TQ�H�;��L�	��ТL���� ��-������`fj
�Gy��Y��� ��2Ps`��%��>y�ZVW��ޝ�0�����Ŋ��H�g��j��[�Ta͑R���,�﫾<h:�h���jl���S ��	(uI~
wc�j�>�ê���|]�ԕQ�Q���BUa�8no7�7�t&mU<�������+Sã*�we!�Q.
�V�&gf8�bk�C����8�* �'�y}��0�d�AH:�pPa��I��A��/U�N
^�oA7�4қZ��E�r<d����F��|*�L�.	�{U5�Q��T.�ܦ�1�
5 ����P<�`X�@M�r=�X$���\j�1�1��	Y;۰�p�1(^�<�]���jȩ�~>wFq|��2p.S��n��0�9�F��P+���TsL4��`�IyQ'�c�vI�be�E��e��j5��W���@%�>|H�Ӓmnj)f}2?���L��hqXz�Cu��&9�*�T�#�V��W���Tg<+Ϲ�@��dF�*�6'FQ`6��M(,P���z�'B%č��s{�)Mv��5�~tx��E~��~RO�K�!�~���wZ�|x���)P�p����zI�^��L�,̿#::j���f�L�N���E���c�A1WM�����w��[܆ŝN"d-Sg�W=ꎋ/�I����et�=g��$��Eɍ{��gjڗB�ᅾS���J�S.��6�v��ʊF�Zr�>�|��z	�@�y@y)��nn�?�v����4��{������*�'=��
�CF0 �D��ʾ�,�[���z������A�N�Y(�����-%��e�S���#ߩUZ����b16_P�}&� RR��Jm�P((���y*y��ft�B#`!3���٩����c��CР�0�!����M����(��B�!��V����Eqq�s'���S���o��X8MɄ�$B��R��$注�I���5d�5ē��4��L�����R*^�����N5���,�����!�gq_Z�q�<1�*ʓ�K��d�v�Ps}�"X�����.(w��Km~=�v/,¹�'p~v���-���~�x�
j5+K0��V6��\�3�yRP�Nþ����7}[��~}�<����D"1���o_��Ԙz
Tb�Xo�0�mj)�̨;E}���i�V��V@�r�O������}��d�Y3�sS��8���Kp���[b�#���[�ӄz���D�����ZeL��Hv��XA%���ji4�'M�|)��o^�ͭSA&��;���/��/S��T���%M��	g҇� uK������P�y�Oį�9ʋ:+BL�;�X
&�_��OC��!���bU��F&T!�O�c�ʕ0�KsVP�)m���x�DKq��C������taI_�ۖn�E&w`	�Z��]ʳ� ��WJe�{p�߹��{�Z�	[��h���{�F��h��4OEJ��R��L&C�N'V�S��!����N��vқ�":z2�sؗE/�D]Q�G>�G\���=�J��k�8#~ph��oU��=G'T�\8}}����7<9�����w���,�p�ؗ�����6����K����!�
-��� �� $�i*�KQy3:�����݈�QNrUPS)�3O��z
T���K��8:	��~MM*Jx<y2�x͞;�`�ʛP�^���w!��A�t��� �Ii6���9x�x%I�^��%Ae\<�˸0-�=�;w��G~���ty�X��-�u�-�Hr5��[��5�:I�*0���O�,"@Q��s@��u�]�P�£�ǰ�tvK>k@Ab�gq��g%
.>	ꤥ� aC���ṣВ�������f��@Sh�IS�1Df���v��H�Y�����P=���>��꧆]��N%�|"ږ�$�;{�Yl�l�f��@0�Z�¼��ŭ|0FKg��銫��D�#m������6�w���s��b9َ�/�T��DБ�/�;�K�$��S��j�V���o����R�9.Zd̩�j*��C,�c�1���P�B?�Gȩ�-1[%�����N�AI�,���V�����AM�-��:t�y�hA�	��k+���ن�7?"�J�תp ���:x�5��2`,��Dy�]M��K��N㲿$r��3�B�۹\n%8�	�L�H�,����LӤZ|�ˢ��`P�T��X"��r9U2���cՔ@S����XQ}�ŷafٳ�k���ͅ��/���G�����r�8��V����j��y�Q��fr�(�SAJ!��4�㠯~��V�^����ʰ�eZQ��I�Y��(l���`9A�a�kb���b6lvHC�>�M���j��B��*)5G�%[6��?W�"<S��6K�j�##�uq��=H����ډ�u	��ZC���p��4�V'ߗ�{uz�̲:�O����T��&&&D��*��p��TZQ��t��JRԙ�N���Ʀ,� T�F�\}����K��v$B���L�_��a�<��.�rU�K���#u7�����8΅�I��g@�k_�Zo�0�p]�h���'G�	����H1-��VM���))�/:E]�8ރ:i�C�WV�5�<�+�9"A��>�Jq�$Lg�[��1K�5��P0�Ey.V,��I�6]��2w�k��$��iAg� �?�R-=*�T*N��b��V`����"�2CJqI���|b�<e�wPT�r�o"څY^��Y�&HH��� !�<��ɱ�|�e�;�e$Ĝ��(�vh>�2p�m�{T�%I���!a���Ԋa�i�۟FzYYʷ^6��s��~栘8�-��N^�ﮥ�hcz�����}��F�I���S����5'���WtEa�Sf4����1҂�� rV�e`W���{D�O���̅����=Qb-E��:��%�� ��n)�"����Mc�(����:E���P[�!�s���p�K��CP0�V�|P�L/o��2�#:���jj*by�.�*:�D���P��l6�w��6�|�=E��S�\"1�����h�R���k'1Ξ|�d2��]D�U�43�#�(���BfS#5h8�ux�$�^����P���_y�����M@����"�m2�o;���l:�>W.�����'@�b��B�$�u��"�P�~�IDE�b�	PZE��r������7�|���؝�=*DT�^\�n�0h��D�QD�I������4���3o����c� �	P��_�zg��"�'M�b�ۭ;�Ԫ��~!�f���В�Ǚ��"�����"X�	��ɴb�7�qݹX,���g�OJZ�@�(����*Ya<�SFt��M�F�Uze;�$�����H�:��y$I�VsP��E�$&�_�z�Z�Ve��w�	|7(�x��zT(����^�n�V�z��Y��H@��؉Zi&f�C���Z����g��� �P""
J�w"���L&�XN�ZqO���ޞ�7�/� �f�z\�`@$چ��U�1�p�0�.��.�\'�"��"
S�Ln�Ms&�Hj�Z*GE�R�����ߦ9�[_Z����T����s�h�qHF���K;��q�	l�Lq���"����mxn�b�l�R9�f]=*�
&��f�n{y�f�^"��R�H�<I좌aZ�o@����.?�d�!��1�b���i��2L�T�{�AM�}:H��v�rRͺzT����ƨ����n�I��K�ZR����"�88�rT��d2��=��Q��1O=�h��J�|wvv��.�b�a'̨�֑o:�M���У�뺏|�h��z�:娈�1��#���� �� �������,���)�	���z��tow���>(
���� H��k(*&��}ccVWW��;}%�'�:��9v����	+++A���?�ޥVyl�-.����� ���7w��1yaŴrҒ��Cd:k��3.��~��7�*;��0��N]�s���T!���Пe��Xs){}JJ�Ԕ��[gI�Ra�e����������uX�S�8i���{��tܗ�����F)u�	�T5�~/��H"�M��O�$\�|��-I�+
DK;��G�������ŧP�����>����M��}m.�*��ׯ���)R��xШ&�Hrt�C���1��\�m�����Si:o���o���������&�7k�83�;b]P�_�'�ϡ�Ƕ\o����ݧ���٩6l�uf~��M�	m��� � ��Poz��	�nuW铰o��H��d�����+�arrf&/����e �GFm������Y�w�5���~ �If���*��`o���(3 w�܁���[����;�ږz�u>>���(���kp��5�ʨ6�A�,W���s���{�{���#���/5>�y�7>��o�3s �:Ugv���C�����>>�3�O�#�!yI�13S��z\��R�8p&�U��<Gj�~�Z�<��͵���K���t;Y���j���e 3
�.^���ge(�ϝ첄��!�%p��`�\�1���`zz��@<��O`ap����l*�c���;��Z�SL��T�ݗ%�$�X�nҘjPw�܁��>�AȍM��� *5��A�K��� �����0�`��`xж�����oء�z�`.�MA!�6��Ԛ8��3V��I����Z{Np����q�x��������R;Y|}��I�d��׫q���7�O�O[�s��"l�w	�'�"~'?2ݰT��W3����O�V`YgP��FL 211/^�ё$�z�R�����-����p��<�J,3�L������|r�.@&��]HSqȔ64�D��*�����e{{K1�C�~������|)���I�Q;��zK�\ �z�׶y�r샜��������O��>����jg��}�C���+-��}�������X�a�Ԍף��]�OX[;-�Y�g�}��T���������Sw���<�|��_�kk*�J�@pD=��,�Z�p���@¬��7�V�����o��<z����7�K����j�����y������iPGNe�l
&�&����/�Vqj�:�PcqP��^��������4J�d�=֬�6E��C~�d�' kׁu���Y=�����!�����5rրCv�L��
�	V(�-�?�]$y�ƌw|�ٴ� �x<H�.V ¶����+�Tp�`:*���]c>7��
 Ҭĕd�p,
:�-N��	H�I�3�g�,}:�5����f o�<#eRN��J%�v����L&C�v�tx	u�_�(��v�^ �e G7���E������l�"���L�3�05���c�����TV)V� �;�i<x ��bN�aV9��sK� G{��E�<
�6v��0Uk|�4F2���H��n��(h�`L�&����z�o"��n]�O��f���iH�M>���Nݭh�A�C������l������O�H�����k���+�c�+& �Iyn�w)��{X�sSs������'�q��&��q��̃��ޞ���;>J�\�9�Ze��}p��% ~�:�&d���]WQ\��K����2j�>1X[-~	H��
�m����.��s�\AIݾgkp���0��!�$0I �CI�|*+H/E���69�I?���x�z~ 2�30::yH[U=�x`�r���)@�h` �I'����  ��h>HTW�G!~!���������[ݕ�(�xwD�U�U ��
�D����<
|�z�jJ�����jJ�ʹ�y�����L���Xӱy�|��.k���e �����%RB��m瓭w�$B��D�r9j+L�D��8�<� ��8�R$љ�B�ML;,�
���r4�F2� �ξ���n�ӧOY"�P\+��lc�zqb�8� (��b�P��z�9\�G��H&Y�� ���$T+[l������� hX�%U2��FC�Y*Y��H�������mt�<���o��Ғ�y3����*<�R�T6�ck��+$�L���J�f3��r�j��/�p��O��c5��0�����%���ΛIg8�<�*蛯�T+j��r-��D�<k�U+�شt��;��ı��yP�����1�f��I�i:�UȲz\��栲W�����,2���-���K��H`��J�������Z��^��߁)s	�������O��a�i����8$SyH�����L:�w4W�UB�=�N����D��q�� ��a|x� ��k{��ւDO��z�0���@`B��Ū�*��:_�,~I�6PR)��0�ŵ͑@��GW�sB�^I����lK1���(�놆�l�K'lF�t�OYӬT�<�:��2&�Ӌs�B<��
 $�yH;S�@��Nǩ�|+�H�}0<:����K��)	�ο�������&�g�� O�{:~����s�H �L���D���v��=�3*xc�x���|�n�^,�w4!1�XZZ�E�ܷ��I�3�D�ß~���1\�ʫ���B��>%�5H|}�[n�+�T4���(;�I�L��'O`~~vcU(�Q���`�} -�skPc�ܩ�xMME�A�7��|��X]֟С�ڼ�)�܇��,..2X���d��s3<�ѱ�B2�4�j��Z�Sw�e=x4� QC��kpd��?>1͠4>���=�p���������G��Z^^�먹��0ޞ�I�Q�D�dL�PC]'�:i$P�mn������,�O���
��^/͡Uܖ�gO�0��5ӳ�������.�sS8�NL`��Q�7�UX�ulWz�A'Z_��p��n����������$J������b��$�S@|{H�@��dR9��1�ӐOŴ#X�U�\dLk�����̊�Ȝmmy���t�D�^�Z75��)�����sc0�������9fһ�D~�Pr�����a|t������.��>�����D��}��yn^y��8s�%v[3c˯�dEu��?�� ����)Ϝ��ɦ�|V�봹�V.�}�ݾ��1�Ǽ��{uf��^}��7>u�5p�
�}���x_�������?dp�յ?c�m��@�ʫ�Å�s
�]=n���A�077KNt��W�ʕ+�aM0ȑO�%s�(w6x|+O���G}���`�DI����p�ްp����t�u��c��3*xó(�u{�W��=-�H4KTvm۷-**�0BR*Iy^��M�$��IrHKmd#�JZg�~`N:��K4]��/edd��&K��F�6U��������.} <�_���P�YjjVָ,˔B�$D��H�R:��Ւ92{:���"�����{5b���i�j�j��344��qؕ+>k6�3�X� �!�b�T�S��,�+4ԟ�f�=�\�[{�'��Is`�~�=���P(�������F���:?��s� �H岐J: O�/��412�c��l��,��y#Ǘy����1=Oq���Y�|{�c:�/�MDԕdq�#�ePAJ:O�U�/'F5��(R�ln�XP����4�M��D�*������(�X_��(��-n�Ǝ��!~�t���K�o�k��R�X�䆦��h&i�ն`g�1<z��K��;8��JhuL���'`�����	d��g��r����nmÇ��C�%�q�^��s�@착G9�����Y*�Ѹ���	s������q�scÐLP䐮���N���7���������o�p�·2*pb��U�4�qm���%���,jO�s�a��(W�P,Vtތ���:,,�P�P�}�������U�����g�0�f���M���C�-���.��渁�Ә�I�9�r�j.k���%��ȔV��PA%^�9�g7PsՀ��9�_�T��P�K�)��M;0#�z�$:ȶ�3�UDR���`�F��fS#ɞ�@HzN���������r��M6;Q�I��o��/i|4���lV��" T���!���e`����F��e���O�}�j�-ʴ�憷���]�c��љ��}��sA0
��Rt�#���8�,�?X`M!;:���~�U6o���*E�IRf�\em�LYtO��Aǜ]�`�uyf
5�l��k!�����jI@DϘ�M�gy[i�3��㣐Nk�1Ki�1�6HS*�*�۹u��a�Te�e��|�c���f�|u~�L��>`�������/�kڧ�lB�i�pu ��E<���W��PɁ��f��n�^"���	(|6� ���e�<��_�
�C&Q`�Ʌd��D�!�ҾGz￵��n}�|�mx��k��8Y�C�m��U;����T �\�Ƨ`��y�"(VJ0��k+Oak��:2�JJ�밲Y��*�@L[�4�OfR�,���? }(�o��|�[j�j���2@����2��o ���{S��n&>��,��l���~��w���tiU�k�.�Bap���L��U���U�./���� ��6���l�*�}��0Z�~*n�iƚM
y��s���X=gz��z*�~X�܆�������V�P;-w���;���~�ܝcsZǴ��߮�Q���JC��:5��7vlt.�Ns����<l��T䟕P�s�_�p��E������L�
E=���5�L�t�E�ԍəGA�$KL�,W"���<J�Dbh333�%i�LB�˦�"<Fi�?�ܾ}���o�+_��|ޗ%�8TWG}�)�@J(���$l���r1E#�����{a(�@E걠�B�FR>i<ŵ]��5|I|^[U��d�U��M�^ѕ�ݻ~����TT�m���H�H�$��y����u��-x�w��Ǭ��y�q_獫��P;��#�<ָ��%�y����G��u�~����iW?��aumGe�#�Ҹ��Z��'F�<��1奴Д��F�VB���@�=�3A��mF�O�W~�W�U[9Ӡ��yAmSK�&�-҅H�x�I.j ��$�ڭ����Mě��*�����m�����O�'_���>�F{��oooÃ�7�own>���md�i��K�	�N�mA�F��D�v��t�UH 	?r�S ?����\����4$�1Xx��,����*��U�&Q2�*�7`e�k���K0��;��G��l� ���p߂��1(U� �'(��P<�5�')o�>wJBѣn��z����E�����6��Aqg�#��T븭�PY��R�������@��x����]y��j\u7�������+�`50z�~P{,�9<�v�.�Ri<&��c�����@���.UǅŻ�Zu�1w񼫏`ms��>���);IͫAmw��>������� �����4�M��l��lcy|�Ⱥf�zX�9廀����G(We{{��"S@�玾 ݸq#�7��tmn�I��[���������Q#�#��j�׮�իWu�+1��ww��ݻ��P(+� ��yo_$����r�SI����
�b�EZ�d{��)��$�ʴ>�>E-�dM���'An
�X�������J<}����>%P�U�����7j�)-P)�Q�$��D�i52�EӤ}}�r�۶�gw���[��_���ju^O�k�}9EE�(�@�7Zb�J�@y�߸p��&�x�
�I�؊J�iP��܌�$��å�.6-��غ�S��6��*���m.�b�$^sl��Y��>�f�5� 'ݑY�G�?x�]Xx�Ur�;��|^��t�}k��v+KW�8&���IfX�cC����K�te	��`uc7π������~O�<���)���!�<K
0(
����M���d-Ú_e���,��H$���j6�2Mg*��i
u��T$�Si���WSC�g�/x�9-ɬ�w�^����MT6Cmŭ�aw��Ke��d�8j�e�gyI&vU�317���ϐ<�0X��}(G/�N'�slgT���ͤF5=Ũ������h�K�.qE�R��/EAQ�0����BJ��^:�F�Xe�6���O����B1Y��<�B�h4F�3��L�3m�5��9��ɱM��R:%LI��BQ`������1�K��=,�J��0�4�*��唦�֨Z����ER[���0 �& uO� g���������$>~��p�yB8{>�N�� n��c�3*8�2�>s�p�n6��Y�bo�V�$�9�OF����`�`��5��'>�޸FU��j�
�ކw��>��G?���a�z��Y6�ٺz��S\;<�c�UP�-Q�1H�A��'all�)�K������682��	pc}*;�@���!i���YWs������� �7��Q��Qs�=�ⱨr����!kD��?P�*�d.�q��`Z��6��{#���!���j~����@i�j<WH@0�Y��6Ƞc���s����5��cq,r��ʺB�頰?E���3I��J��q��L�
%>�9�Һ�I߉N�8���T��������������9�>��~����|��QC�5V���;�1r�*��"gf�"�E�QR`?j\���"Y��`�*-:�VsYG�б9����B���Lt ��`��j~[F�j���#��G0w7��I�ۏ�]�YPQ4-1щ�I���sv�����f
�p0	}�<K㽉@�of���v����i����K	t��HAD�W�X2����o����������ܝ�����臰�����"�(2�Si/�vZR�Q|6��t���:��#T�F�`���L�(������aH�Jò��p��e(O_R�?��q�2���>�cligb�^#��F��s�#��T����x���Wa�ʾ5�CL'Xt�f��?0(,!<�3��2���\(l�3���\4�Eu�V�T�0 ����+q�t�Ww���p�W���}s'E�?�slgT���Q�맗�ט�Y zQ(��ڵk�5M�?)�(���P���w9���(�po�Dޜy|X��f2�G�(�|>���ʁ�nՕɎ/>�-��(�4ddb�J�M3�~���[%�v�8�A"a�r��v�g%|����coh	�o��̿[F��(�Q���f-8>vpe͝.�M�|j�k2�kЉ�9��,�P����T'R�k%A�4?��z��Sw�������Wɍn��M?S���?	��2i|����������)MB�F����⎊ҩ��S��THo2�BQ)�ua�f/mC�w���p.�#� �jV�ON�p��%�`�p�.���@ v��玏����$u6k�G.���,�������{^2�<L��r�ǋ+�C�)Պ2���=��s��m\3��7~���L���]ô���0n]���\���Ą	Z�����lS`�w���(@�)��:QR",9M,݂�ka�&\�U!i%O���	�35yY����f[�u�|�̂
�{�=�Rb��R��c�����1a8D"�f��l)ҋ}�9�۫�[�����{�R.W٠�L�dT��@�#�1U;jsuME\y:S��R��`�kJ�%���S�i���'kk�����|�k[սL�P�F�� ��>3���>3p5����3Z"�
�ʌHS�Ga���74��N�~�bТ�u����%ܸ!?[D�1��6[I#� �a��!�_�e�[�$t��0�����LϜ��T�Mu��t����ZGµ��QF�a�O��O��GT�t@}'��&�N�Q�~@�-O���>����k�O~��055
�_���{��߆~�{p��<jETO�P�I��\�Ȱ�&oܸ
�/_�t���.�`w���#��q��%�1*�5��tB��`zf&&G!s�^ڄ��Xy<KO�9��Jtk[7�R�s���؏����y(��V�T�.�A2���IG K�Y��
.>�	l��MmtK�Mk��@�SR����b�ڸ��M9CJ���a��ɏМ��*Z�B���}PEZ�˱���7�o(��&q�W�TB7&Sc����!j1\��^)#Ȣ@Q�%���o�x�^�Fk��3*T���ANt�f��i�;�$�dʡgOfX�' x��WP�P� �[��UTq��N��E��S��߫��4���)n���O��e����|��GJ�}�1�R��}�Ae���CP�z�B��,��h
 ^e���E���r�K�$hm�������fM��`��_@���lj�~�QOɥ��>�P����;M@A��φ/�9�1�����>q�c^�A4�[4�`�M`|�H��\U��X��|yvg��	���Fw8�c��3*8�bx#���G�O�V��^ �*B��1�*��}#p�7�ƍ�0;{rz�nVK��3�0{����Td��c.J����`0�vi�������-iCu^\[9������O��{�c[u��%20��87^��B�kd�7�PK����U��*�ג������^��(������^F���2��\�Ie �_���A��{��~�P�*���*N�.�h�������<����lxS�Q�m�4��Y&'�=���u�؛a{��߇���֔�xb�<dr��J@*n��l�k���-�X����5������9��m�u�dʰIP�������xfA��8�Ԃ��J7�WzI�jDl��g��E��	
�T�H&�EX���O�=�i�����J�.����J�WI�y4���jV�+!��KH��%NS���z/�Q蓢��sN�ʁ�$�:J�$E+[��N���JgK���YVU��d�5�5_���&_�D��I#'�Z~��oT@��}0$�l6#������ϭ��4'̓�5Ʉ�HNGkJ0�,��$>)#"z�RgM�T
Y,��{&����ˑ; �x\HgT��I�2*��n�0��q9^�M,V~�} S�~���!��؞
�Hf301=��	��eS���̜4��u�c&�b�����B�R�z���e��R�'G��NL��GQCl��%Q�)���Y�8�c��ָG}5������2�%j�mb���d�s�Z�r�(�8�� ��U��b���s@ ��V�W�\,C%�U`�)�.1])/�E!�!�0rb�ڞ�#�7����.�H��@Bw�q��$3s:F8�N@U�@��a5PV= 7����̌���mՂ��,�x���061#�܋F]��!,=y��~O���vH������T��~jnm�
.��,fA%�$N�v��{E�v[;�(ڋ4���	� �O�M5>'	fqIK]']X1�e/ז�E\�Q��$y�%���㓰c�c�
<��ׯ�XS����h-��iIi*�a�r�Fb���F�Ձ�,�A�"�H�^_]gf\qU�I��p��=���2)>����1�<!m�P�`���T��|&��sбb�#���_��M��V+A�0P��y��tޘ�����^�s)����s������XtmT}��I+����}�i��ϟ�\F;��ک��=zw���jb
��@q�5#m"������̂
�����A[Uh�9��Q8y�5���r\�p,��.�¿��4L�ӷ�*�B�-�M���)����v�zI(���L-H���Aܢr.N�p�|�}���d^3��o|�u����T	����g`��Oò�df�zY���*Lx�x��L�bt������)�i?�Rgg���㩣������JɅ��
T)B�$3��,O_�7.O�+�#�F����-��[�Ne`t�:���a��l�oAus�)�Ff`��u���r��gȮ���҇`0u�p~�E�6L�k6����8ܸ~΍��[��䏩(Gy~RSUx�J	v�v����(���їm�o�!����Z\�;��~p�3p��{��>��`�=��ׯ�����p�@]v(n=�w��{����w`y����z���Rug6Q�_���)b-�f�4
���7�J�tb�~���8���L($��'=�
5��pc�i�C~��i��P�ݒ�Y���,ܭP�4Q�!�M5	��Ic ���r��ս@������f:-[�;A��H��ē)>�zÓ6Q�!S�t�VL�K���0b�/^���u(��q�@�1ZH[p9���b�ڼ�|��e��@&4�b����1������;ʇ��*�l������k�K$
�}Sj��j>WP��}Đi�s��B�Z[S�n���*"�Q4:7	����oE�B���|l2�qr��6���[p��Mn�@��#���(�N9x6��1���F�
R���,��ޏ���d$u9�{A�̴��nsfij�
�ԯB�(aL^ӧm5�͉���/���.�)����c�k��9J
�4H_>C�H%�P�����V����6��N�Q��룄�4�*�\^���:$�x�x��!� �loo����):��V����rtp&��c@2��x�
}Ԯ��7�W`o]9�c��2'_2�z�$�LU�/�C>���,ΣV�+_C�R}�#"�UQ�Hg��f;�C:��l�2�K����EQC�H-_��h���!K�9��!��e��c3����JI�p<F3x_'��P�sx,�t>2�Q^���c�;�o1��o�J��-�d�P��O�4���L`aM�P'qD��73�/��:6��#�z�DE'�p��}d�5��W)k��~~m��d0���KThP�,{dv뫫l�z��iAM	(t�$,�m� �� �L#����ğg�EQ�sunb�$��x=R�wt� ���$I�$���vT��j�I��'5�"��enTTe*t<�J�fʓ�R7ۛ�Z3���c�����H��CZ�zf
�����\*��Kf/bhT����>}�V9�A5E�>���[�
�J��c)��tL�}ks����p���'�|m|-�1ݞ���4��N��T�J
�}*/K����!�u%���Q�߄;�>�'s:�Kۺ�I�߇�T�|]V�R�1�Q�(f0J�*�VQ(�W��u�V����2�B�NL6(C�4�^*w���dq��CV_����*ܮW`a�-�7������U)!Eq�FD�r{Gu0�7��Q����#�h:���Ĵ��K����P_��~��s�`w{�#䈁�uR���Y�����*P��-C�V����q\:�ȭ5=7�4%Ǆ�?�S�x�Cb��M_k���C����E�u�>Xٳ9��s|=T�Z�����Xc�S
�d�aQk<.>w�pj�|>���4Q��c˪?��Bat�w�&��%5�n�K	��
�"+QS�������T�_���m�G�l�$7��ukJ2�����NP�n��|t<b~��{�S�P���JG�%tȯ������vu���kz9������5*G�WkJ��.U���5U9a�� )�j�ǣ��檊 ��gd�v�e1X�p`8�Mt�L�ܚ0	ݻw�;{�n��J
I��7 o��mrPc,4��t�)�0o�V��F��2D%	PE�3Q<Q��Y,5[�ȑ.�b5�����r���Ĭ�X��zh}WE3�o��>�3�ә�&3��9��asoے�tW%�Q�c�r6�9H�r��%�4���T�m���1�)�4��;��rD��PL-���1��+��\R�/���,�>ڼ&��V����u���.�C�O��������Tf?�l���W���X<^jwL�Hi5�-���!�q��ӮkA�VY��-��m����>�o��)��5_UVPs�;�@_�L��K"Py9�ַ�E垇:�L"�;Ȕ&�ى_��@�G���&��o�������� ǅuQ`��cML*fK�rs�)3O���$H"�]�G�QxC�1����A�+#�݂`�r_I��%�o��XK�c����g���ǝDP'K}j)�i�����_¥�@���vP���-���I��r��js?�9R���3:��rt+a�U���h�!���r���6A?3�1�T9����o:8����Ҋ֐�6��㦃2�3AZP���m��0,Ƿ��J4|��7��{��g�(LbN3������WI�b�s�qMK��X�-]�,I�Ծ�P�T#������t�_���1=69���B�d"8��W����}Z�\�+�GR��fG��Mi0u�,�L䦳/���뎹|,���nY]�<��>�g	y���ZRɸ��.Qd��P�M}\��	ҙl_�&�*���N�v�I��V�d��JD��������H$
�qϔxñ�a��<���"��35�@k*� hs�Ө.@x&Փ);ߣh4�	�/�;���-��i�z.
�0OC�M㽋4���T*�V�q�������V>�X���}�'9�p��@C	繴��f}�Zm������rִ|9�tO�<�z���m���}���(����������*��Z����4:6�q}"Ź1���ɠ�
$����X*��i\����Wwk(Ba��{����D*���S&A��I���Q�[�O��tD'��t�Et������ɢ�8�F�s�.���C����x6��.]��,��|�C�Q�M�Q'@1����^g��r���$��� ���vE<dMFyfω��u��Yɷ�$����Κ�A5�Ƹ۝o��5'L���kB��ŀߎ�>��/��7�ph����\��f��ko��?�I����4|F�G����y���8���o����[�=�8�fW��7ԊN�����Z�Z'���t$"��L�J�V���r}���
<��"�&�H��I�˷"-%�3F�(,��FzT��J�PM1�;�Zi��UnY%��o䀧m�F����0??��n��k$~*�
�*�G�	�
������q���S8Q��#UY���v�2�[i0�.M!�2�A�(!@Hc������lg���%������aM��$�~M���Y߂���}i}��i绩7�e�P_�k����l��=�Zbk��p��M(nm�mP�]ͭ�|"ݾ9�C������S�W�\9�ª�g**�󆞋��X/����J�����q�~F�ʋз����,��
?�71+�����b%�@TEYt�4>����[���� t_g�SY�9F�jH�sA�^J�=��i������j�r��j�I�2�&�@�]�&�N��x�������~�g~�E"�L.\��D@������O����ҥK��� I�$�	�����ƒ��jd��f�s �*@��8�C�Ÿ��ğOr���Q�5�}�T����$�gv��Q;��_k��~Qa���7�F$�Ҷ\ΐ'����UQ�U��P+霒69G�MT�ku���6���®�C�Gƽ�͂���l��l#�x�b�����W��G���/��/����ԧ�][[�\�re����}~arr�gQ�II�o�Y1Í�=�� `$��y�U��>�ܲ�a���R��<
���HL�����e
_=�$����.0�\�}筪~~�ypf8rė%JKq% �����׆ױw���p6"+��iː`#�XC�'X#��,8�ȖEb{[�	)G
cّ��I)��9$�������=�����ݹ�]���Ws~����W����{�eLᥠ�ۋ����c�y?�s?w��ӧ���v����o>��3�X��!�~�����֏_^�aTipO\�z��n��;�}ǎ���p���r�{4N6�R��N�Ba3�&�M���m{���/M�z֞�p��I&Ӑf��ǖ����t�.*蝀��v�y��C�;��(������'�ﾭGy�&X翿�;�;�{�����gp�'O���x�0.G/�<�=�� �_J���[��O�g<����t�4�ڨ��y<�x:�=i�������*����}��:w�����6���,����<��_il6�x�����ʎ��Uji��f�y�&�!|6���c�A�x8�n�����j��}箻�D�Go�������֥nغ��u8�s�̙����+���ѣG����E���"�;���!z����T���b|�{���bZl�0��wTq��:�(�#̓G����S���.d�w��a��#���n_��qv���(�V�Eq~��G�3C�9�g���^u�jt�9��q��J�����oz�gև����︡���8_Z^^~����_��ؽ7ƃ���S����V��o�v�m���-��@,/�������E�qB�^Hl��c[ă�I}	�y��H� x�{�3��U���tl/���_�-eJ�����f}|1z�!oa�z��z|�Q��9����~�6�j����ڞ%���?(���7Du�+#_ݲ����5��V_�F=僡#�ECyb��-��r��hz�h��iݼӃe��:{������B��R��w��	E;,␥�8��/��R�}PJp\'~�ua��ܺ(�:
��{�Ah�I�L��J\t^���(k4�l_�b��!K��~�����1WQ�˿����&%�����|6���F�ӊ����(��� �����ꙥե� ���t�Rk�۽K��];vLa�\_5[w���n��j)��u"(&��琌A-���:y$�Q�z
c!�T-��71�(o�e�P7����d&��b��o�l�<��u��d%묏'F��\���;1Q��3�W�q˷^���JDe���71�����'-�����5\G57��c�U��N���ݮ�G{	�X]}cMm$Êz�,_���ⰳ�j��!d�ѳH�M����Pd�<(��)E�}��xHT&"�^���h9�����I|LM�I�h2���ϡ^��wqʾ@U=�0�ZO��<ԗ縦c����Ϭ믯��+�E���?����K[�JOq���[�j(S�x|?�n���N����
�����
�C�?Rs����ߤ93�J�x8)����v'���Q���CRA3�20D��7�M�K���r�ɠ=T�&��x�0�B��PH.��'�Ⱥ'a2�������\��0�v㌢b�/'����vP��4�n����}E�aۆ�e�3�PL� cZ�M;�Yq^���#�i�mMX�����;�.e����)���lW �Ԝh�����y*�dМacb,;I����f\�? ^��T<�����6�o���1m5����q���ñ��D`��{�8ki,2,=yY��$*�̔���׷�:/=D��R��q�7C�M�OǎE���?�΍��XT%FiC�}�=F��i� ��f�U:5��=�j���3��b�
�M䳄�o�'�:�O�9،~�犰u7(���t]�c��?�O���r�;_T�cl�S��x^^0���^][�^}�2�������l���D��7Z�8ȅ�f�2�4�5V���^�*����)�i9�wVe4�/7���f\Ċ��i?�š�g�a��q�%�i��""��:1�i��uQЗ�uJ3��K��+��x����ocZn���uL�'M�x�n�<�%M<�x?Ӯ/�;��4L:�Z�6|;X+�}5'k����q���v;�?6T3t�q���wF���^��V����#ul<)����w���Eq^�!�B���`��m�_�"�Q8V.LT���=���!���/�.@�)�(>�
�G�&C�����.&6a�j����ĲN�R�4�fܧ1iƹ�/2߶ߴL�6/����6|��Ѽ���%*6����L�9�����5үWں����Gi����<�d/�0�UUb���9��׍�����V�?�;���~r8��խ�8ȧB�Q�B��W��R��"���7i��$}M��Ӆ��Bʆ�1�D	��[��}�B����I�����8|��|l�k��Ȭ3��>O��4�li�d�l���Q���ZU̻0Q���<ˋ��m�;f]4��0-����y��d�L�Bvm��5կ�<\N�� }��S�ZN4�?��k/���+�7���� �O����q����&�Q0���X��588����S+��� H�7_~���<$��Ѥ-��$�[��f�oV�!����CT�Dy��+�&/%k[i;϶Ur�� <�"�O�DM�Ӽ2�(�y)���c�*me�:�N����D;��B��LR�,�� ���	?��[n��;���LR��5���E�7��p0��`�3��O�����.,<�H����
����7�o���d-7����3U����ڮeފ��z�����۶�h�{ބ�y��d�����vEßi"5ͳh�>�>ټ�y��l��9�i_Iy���u~̳ң�Y��;����V端�|�Ol�ܿ�~�J\Qś�ѓ~(]��M���}x (�8���#����xQ@6a}�gq�Ξ��F�BM�0%� ��������׬�yF6L����W���f��t�<ǘ-fl��t������J#:�u慭Dk�����|bѵ=;y�>�T�L�^?��ᷪ��,����o�2��
v:{����#<�w`�+�'((�K(�g%g����=�yQgw��y�pi��H�4�:���a,"Q��X6^]�����y����#��r�+z�E��{>Ӭ�EUe"�q9(L��@"7�>�y�g�kY���U!�v.&[��#�@1�B;�����a�L`E�by*�o��_����������j뎫C���\��K�b��7U���F���H�R��!H+���o&��J~��E�z�t�*ϱ�����{�Y/@�mm��Bh�ד��G����
&Z��6���{�wUϯ�����.4�eݠFwp]�����T)$*����~�x5l_��亱�
���}`M1�<JQaI���c�k�WT�R�N#4e��DY�U�G�gp�F�E!��gt��?�yz�
�z4#-$I��Y��s���jN8a�����Z��mDj�U+iZ��]0o؞W�Nz��Mó�� e��i�n���Fm�4	�iߺ(ٲ���m�����{���i�)No��Eb���1�*H�V}���QW�<�b�5*��
w�����o;��^�&l�A���$��>7a�_��"+?��x4:F�X	�m	��ε�~M^ �^n}2�o[n��<|���m��S��������N�����Ӄ��R��Л�)�mm�U�['���=�,��pU\Ou)&��[h)Zx#���(��E"oT���J��X�&���w��T��}�Rop�uS;��7}�(GaAw=�|��� ��!�����2��m��o������ ��MH�M�F�9��4L���MT��i���d1�:�<���@��h̻ɲ�<�z��I{�L˪x��2��_d�y���Mj�B{�'N�X�:����$x&�_YY��K�.������6sC���@S�aG��H�����4a��!![���Ť=�&a��`J�{[�8&�U_ΓhR�̴f�6a-b��K���8Y�#���ͫ˳o��F����./{��{��������{�Y�`^O$���������hZ�&=z���la�5'2EN̹���om��xwe�#o�z��5��R���&�T׆���$��^�($�l_�.7�4�dLh��@��'E������~эՏi���Y�JÇ�C�FM_�lI;�%��$8�:�2�/{����V���o�}W��
�y=���G�ն/Sa�F�H�i�jS!S��v�t�<��bm�ӵ�y����_��������7���v�
N@��z��j5n��Z��#N���_|qO=�q��D���L7�Fg$�1]`2��E�sq���E�������#Hr����'���/�0���^�,�*kty���� ̂����"�����W)(Ӭo�^�z��6ͻ����l�-��u���QS�e��ɖ����^�ߨ�#;����Y[[���׸�-�~����z�88�G�	�N7t\��n�o���}�s�g��Z����7�[AO�I0q��"��ɛ�!�8}3�߬�0�y�\`��FE�Py.{����h�?L$P��%�ԇ'6m_���˴t�YS���e�"�R3����Pt�<F��:����0y(6a1��3�GG�sH	f� �On���`�Ji�vB����Ν�_�����Sw��ܱ���EON�2bR�j�r���8���B�9��`pDn����3���ޔ�0�yp}JM��P���	}d�<np��YzU�AW�ϒ<Ϗi�n�Җ�Ⱥ�E��"!�<�Q�/�M���i�<�]�9f�τɖ��·�bOz������3���FowǸ@����Q2יL>��jz��Z��ƙr���WV�"/�_4rḧB�/���X/E�^ :�/4��tM/}�Kl:6��V���J��1�B��~m�~�뛎��,Rh�:�4����/������Ӵ.��'Ln:^���^Z��%�}7�W�c%z��7�u\��V��i����~�q�z�P�/r��Ѕ�3���̜��;����ͽ��F����$�|;@��<��"3M	\(N�BM�v�E[�)��i��GZD@�	Y!�"痵S'����'jhdڏ~�M��WR��`^_͑�m�xG��rq��9����fÛ��j{{{���aR��{�'������}b��������fu&tqx=�o����<4�c��-��E�����WV�3����w�F�JO��R��C9,Te4�l��}��L�M�"�������ׅ�D�1n*�"��T��֮`�|��ۨ�H��ѣ���p0��9-'rN�1A�6=ouy�{���a��F�(|D���[^^���͐� �՗�e�����x]]\�I�M��4��;"�>MM2�P�=>lL[���:�S��IU�0����sSxj���.�1L�y8^ߗ����˅H�q�J
�(*C5G?��?�����w���y��>��*������ool4�(�q<�߻���o=ǻ��nް��r��y�/���������
"�~�-��mll�1��m5��ʕ+'Hy���KKK�"�E�e(J�\�鞏=��tT	��`��\���$<����d��'fi��T]'���x��A�<Y��bC�M6ӾU�e����5��VQ5�ޘ�Y���-�x9���i�?������{說���E8ٗ~�~��|�����^�����'�0|O0�0\���3L�M�w ^�ӗ.^��#��C�k�z���(�h��ɻ���P�����t��!6��'N�P \�رc��y�7�D[4?~<��1)lE-x�7���R{����U�bYx�C� \?��)O�=/�_��s5*�Ӵ8�&iA2�;���c�����g���7�Ap�x8n{m���h��v/|�s�� ��������ڷ^�t�]�k�,/��YY�؈��?�J��p8��:x8����ﭯ���W^ye�{WWWbkk�
R����̿�$i�����|���萗B���$A����n���P��<�x���:��A�=�C_e;'�;slN�J(�����
^I�k`ގz��gw���;���?�|����������?��D�#���7�no���ӟ>y��/^�Z���~����p4�F���'��|�q��{��O��;;;;{�w))��^�,�.����ᡲy������ ����H����%6e��y,�Q�}o�SO=տ�ԩ?
����~���ɓ�>��ӯ����o�F�8�bwk�m�p@L�y��b���?����O��\>{�쏁x,Ӿ�ΆB_(*(.z}	�������2���[�	�0{���R��gQ� �W_QI�ٵ5����}<
~AQ@��|��'�����߿ϝCo����_�����K��<}�w�J��?�K�4�͌�j����|Q��n����ua��詀ݛ[�bdaD%V�sIc�W���_{���8q�'����:]�f���"���z)��P���m����6m����������?�<�7%��՟ $*�W1�>����"�G��TY������Lf��ٟ��J��+�������蝲(5�A��A�ޅA/�"|EU��<�=?�^0��סj��h��;{��5�G�� �!�����+�hu*>���YQ_pC|S�w�Uբ�K$�'�S�3n���<��+�~Ɣ�e��ETʀM�LI��n�0�� �ckuJو�.�
[��ˎ`�R�R�!{��+��]a�����Q�ޡ7�MT��h$�JIB[����"y"v�P_xb>D9z)�A���� �/�e���!U�fE$!1A8��i���ּ���/㭿�"*e��/��TQ/B=�{��X���W8����`B�f�)u*e�3�7Cަ{�Y�m�:_�e��L�m���P�)�=|��ұy�ɼ�P@���}��.$�4�B���P���E�sȟi>�����-�LJ����w����o��=���Q)\ؐߤEG���q`����m�0u��女�vi�%Z��p��3	�>����gIU�O�>�V��s^���MVc����^yx�<>�-�o�B������PR�R��u*���ddkpPS[y��t�ɻo}?��Fޤ�_���Y1���3EKԇ���P���7���3_E��	z��1��V�%�J�N�0�6I�����ଐV�H���!��C ��,�mha�Ǵ�2�3��*�Ƣ���**|L#������S�x�s>K/\/bIBa#��/	֩&Q��!��{�&��f�M1a�\_f�����e!�<�<����A��������--7}r/�'���I�(Rp���OyyY<�2����f�dά�UL�:A#\�/ ݋��B��Ĩ�9���ƿ�%����+{NU��E��l����	_rQ��[�o�~E¿E
=<��$����ښ�J�fӔ���:�Bk����`��Jq"Qх��P�����Rͪ;�wP�gW�6y�����gM�n�O�(��]�w��|�0����@��ϴ�K�T`��]"l[������gM�D�c6�pfEه�f��*�D�:o�ȯ��HLۺI/���~y�K?n�����ת��yޒ�i�<�1�EJ�@Z������<=�m�6U4����e%�v��y�T� 2��1�i��,���y�v|��������tC��LM��ۙ��4�BY����E�fQ��cI��ei/j���yE�,m=�y��������G﫥�i��4A�6�Y5i�JL�-�ߟvO�¿zX߿���4d:B�B�U�~$�~��g����2�EEQ�L�-�м΀�t�c��+��8��4?O<6.zd�������^E<1�9���Kɦ��ut#��>?mi�/�-t�E�gt�uҶ)ڙ���Yy~D�;f�lb�ϳM�1���Q.*<|M�����g�ߏ�k�۸l��G�Ο?��E�De<iO7��@"��T��п���~p�\@��MLޗJ߆�1��c��c.2Y�#	��9�W@�f�J��Y�U�nY��έ�
�-
�~&��&*���"���=]T�>�9��)�1�bQIR��a���ȏ���w�����$4$��發����\2���7I,��~�8zXfV����p�5��k,M�m��?��S�БvNUn�������c�Zt��ע���˳m�;��o[�,m{:�M詠�t:�����F��3�0�\�!���<ֈ��Uy'Bw?�<����������-[4�
�H�*�0��0m�0�wZ�4��;�'�v�y���1���T��T��M���ק�>y(1�/EH�g��z(�eg2�׫�\ZZQ)ܔ��p�O��`�4�(t���,�����6����������'\�v�M����t�m�$�KI�Y��6�e�h�����e�ݟ��}�<�"��Өj{���Uh��}��.\4���z���u�]l�s��^�w���S�N}�駟�9S;Qi�ۻ��������-�P�Tt��J��:�#M�<%�i(j����v��h�<)�lӍC�a����gS������S*��>e=?z�V};Sx6띰�;�lh��y��b�>+|�T鹤�wll��Ad��ce<x$/����������?;~����?��Μ�R�ډ
��A��:\�.��	z���p�J�:� �R�i�~mƬhh��C͍AV�$���ǛR�Je.*EJú8�zL�'5�5����>)WT�~Y�rY�e��m_�\^�C�A���n����c��ͅ��u�Ԛ�/������jp�����]��ں���/�3�m�o---�ۮ_�pa�br���ډʳ�>;:{�����/<7�]p�o�a.~�7�c.;=]|u`����Nr������_g�*$�ö��x9������8� :�~\�?�.���s�?�Ӛ8��FB��6|t`j�y�ti��mY�p�/�m�i�Д��x��A�R�,��v�Y�&[X���Fƴ�z�Gx�2�-̓,_��m�_T0�>W��^�Ԙ�S�ύ·�B�'�	����@D��_~����Q@^q� o����>|�g|�,BX�v��\�x�*|�	����Oz?��?������pӋ/�������$<N�Ws��+++_F��;;;	U�����ƿ��F#�2�W�&<dM�/
j6i&���<X+�'�D�H0̤�����#�L�w�h<��)��55�tX�f6۟�l��<��7����o��<6y�:�4L��T����d��U�ɖ������{t��	��) �Q�M�xjH���"r��1g��k����a�?�y_���_{�'��p�"��N-E�Hn��{N	��ŭ$�����[�q�w�=�P�ҥK���y���dx။K�z(��}�E��R$t8���/�?SSB���"=����Rچ{B蝜<yR��꫿������g���SO=՟��:Hj-*�tT\�7��Ɠ�w��_���|����m*���:i��7 �FLfMي�,f�������A�0Ց��;�1�}S(�i蝼������=��/�zs��U5"*B-����A��u^��u*Y�|�d��T�zO/b��U�^%e=��=�����������L�B�������}�k_{�9D������~�����~�Jt&OFu��Λ��;��gE�yO����F;𜽡j���P0�7����?����y�c:dt��>�eZ��(�阎Y�~ښ���{�<����TMQj��s碇~��ӂcx���gB��05�-C���<�6ȳ���}��æ���h�=8�H��.`�졩_I����/������S���-Q��V"��Ә���	N<Kw�k���Cw��57��7�uq�X��';�܉�¢��ׁ�a!*�a.s�<}?lW?����z��i�|��ߜW����Y���n��i~����m��N�ղ�;?d��� �A�9sf��i�����KX���7��1M��4�3�������*A�����Ńg&�CY�m��/�'��J�{��C����t:"*��h��۝&��n��>$��_��<�@�e��|��s��m��s�����Y黎��Ҩ�ߟd����XLM���� |����C�7�#�"ԉ~ђ�^
���2�'��(�T�63�����Y����h��N��uL�
5���\\Pp�uLBe���c��9z�h�j���P�݅&&�k	M�*q�S�o����f���?�(���4OD�V���>O�P�&��TgdZ�+�i�$�y�}?�����Gt��¢�n�����1S3�.R�z᯼����}h�D%ﱧ��1�Wȫ��~�Z����?y>���qt�����%ᴫ�ϟ?������ub��>�U9�?��ϛZ�V����Vy�CȰ�!J�{�o�l�lU%�YGѿ�*��<��-���Ͻf�8���7ϝ;'u*��h��;�3���n踁���p�*�!#���^$*��m�fgE��p�RiM�u�0m����H�wm�mU#DT�� /-8*�.��HLk`M���j���$�B����@DE�KKK#����y��H�k����֢	g�
i��+r����-U#DT��0�L#�ñ��S�x*�!oc��XBe#xfwU�Qj��___�$�dK�ӶV2�I$^���HTu��:L{��!�"�l��g%�<�x��#�J%��N��5��c�b�VT�Qj���G��ZFF�z��~;�lX���F�������\]4Q)S�n�K�J��b�OIk�>- *;�1T5BDE��,��o��������xP�&�*c������u/�O�2�R� x�y�k>\^���o4����S��2O�WDH��<��T��x��"*B��R�z*�'�a�V�fKV�Ȋ�;h�۵KQj�����yQ<�*�?���|����m��D����V`K�EӤ�Oe���h\A}��>�S"�"�
xQ��Ѩ������#��|�u�j<���ի�¢��
6�TQM�D"(Ǭ[	b%}�Ѩǃ� �"Ԋ��%Д�O{/Ӑg�i�ˆA�3+�� ,*詄a�E-���",��������ϛ执2���~+D�����s���O~��<�ꂈ�P+vww�N�ӣ������w��5��x<���-��Z�V�������3��߅�CO��M�s��-�:"*B� /%��z�r)��HOs<I�2{���.��{�ש���"*B�h�Z�����0�"��A�	]�Tu�u���X��s�j���P+>��D?�C?�7>��0���Oo���ŵ�����ԫ[H�V��ѠGi�2�Ҿ)��4�"��31��,Ԫ�7��Ze(FDT�Z�-i(뫄�����@�gS`���� ,:!�[�����u�_�sB}���S�YA�IL�T��{곂����ԩ�!`�\S�V���^���*�DTa�y��g1�U��)�������
�T��ԩ�! <$�s�����2M�
o�A�
V�A��j�j5>="�"ԑ��T�~���TC-�0�)|J�K�Em���x*��A�PT�c�l6�"*���<��ѯ�����f�4�/=(�k4���"�/A8,��L�4U88ʌ��[q���W@TF�f����*���1L��t�_�@_|<�Ti��V��k��P=�gD�х�*�_t��r�Z�%�PT|U3DT����oB(x?6�꣏><�䓪N��B¬��5�O��Pų�C`�k���/~�P4/���P[��y�l1S8<�y>�Γ�粁KΟ?�ꄈ�p]�f f%.�i��Q���s�����,�="�"ԑ�U��O3|�JZ}�x*��i{��^��J<�-UCDT�:R�8�ppT�a�V`��ümUCDT��/�B�i�������Ǳ�����<�v�$�v�K;�>&��	��/9o�ɩ*fڿm��Y��0���EԔ��8��A��<A8$d���`��S�-���P+�5�ѣG�y����Я��J�|�����q��@����K���8��X<���ä��b�2ʎQOa0Г~��Q�� ��{l���8�&���I�n��{��aR���Fנ�
DT�:1 ��J��\?Psb�_G�OEؤs+Q˯4í�:/������X����x*�ph4>e���<=�<�����*�~O�S�Z�Z�d�v�!����E��߂~��2�|����	�0<M�}<��wmm������P;���e�+�*��NL��|����^U7DT���y�GS��{��T����᳿��]�SDE�ौ��`{����<�	�"��P��Q�𗈊 �S���1f�m/eQO(�C���~Ν;������%��U���+����l�=)%_�qꄈ�P;�SA	��
I��P�i��<���"�P"*B� 1	�0R�A
S�|��TMQjG��b̚<>�
z-8��f��[�p}��4OB`�?z�t["P�>�:��>.�G}mK;"*B��x5�XƗG�[tD<�<u*��iٱyݺ!�"�l��#�a_�����e����Fe,�����Ïi,^��Z�8���!"*B��t:>����2a�k^C��؄E����t/���)�T��!^�x(�z,;-F�K��4�6!���p�Lۤ�<ʖ��z$�%�����"�"��i�G�ςPx!�A�����ꆈ�P;F�֩\!Qэ���{0�4�z�/	o->Y�H��㙈IPt�9ADE��ԧ���.�թ�Л�V�)ݽ~l�>�:=aJ�� ���/b˚�S���C�&���S��s��(JU{^�5�O���9�:�d惩 a�\7��}p�g��l�#��5q�gSDE�>�h��Oz�6�J^c=/�A��Ë)�E�Du)�����Q�����n��f�"7l�O��fŋ�Xt�@1!A��sOD�W5EDE�%���AЃ�G������ ^�b��4u������$�#M��0/��������c�yE�<����E�Si�Z��G��������IUMQ��=[�<�#�$�r��=�G�Jy���.����aHDGDE��0S�i�"r�?9�Px���nǟT���S�X���KA8L���J04�����
yj>L�*�J{��~��ԩ�a"�0��)z�>�ޏ�ǿ�|Ĵ�,��x��4x	זi��w���gI^��s�T8Y��e[�[
�I"��Np"A��7�:�T��j�F����ue����Ph��776uJ��/BZz>٠橼w�>�XeE!o�������)�fھm�߶���osQA1�_��C`�
8�<O؀DDE��F�ѕ��%k�rSɟн��}d��q=�qM˜�3 �i"��!9��eȺE�'m�2�J���B�x��W(���3�B	
.Kz��t�]�"���`��67��5z#6cd�Z��$.E�$ne<�<F���״a��"�'��S������wAu%ت���=�\��wL�E
<���%��#G��7�n�Qύ �4yӒ'�ŗ���iy�_Y!���[y���)Ms�M������<}}1�B_(*z�:w����J���"������a�����~x/���ti3`��FI�HE��[/���1U
����0m��2�\�1���_�>m�.2��p��S�~'y�^�7�&� *W;��ԩ�a�ܹs�C=�N�TZ��R(֍p�΍�L�4�f4�O�ZLcqL+
y+�g���s��Ϸ	�>?+���׍=�7����hO�D�����=�|�;���z���A��uIr	�!^����ӗ� ���nH�m��H�l^B�1[��-�@�-�l�9��}MV�i��	�MC�i�a�(�^qϑ{�iBɗg	*|fj6��k��LL'����HlR�ů~���x�UGDT����"�����[y_43��BR��ۖ��e�j&�}�u�����
��碋-�	����)����c�S�x���e�����Q�����9��]c�x�BӶ��x���G��{@c���ֿ��F��x��suuU����9�����_*����v��z��o��-o��V�u������n�2�T�K}����4/��~h?�b?;�N<a�] u�H��Ϭ�pS�9�����L�3�M���x-QX�\�������y�ճ�o���`!�ɓ'�3�e!������2Ɩ\@���~�<��>�D��������I��"�"Ԗ�{n�;����	/�} 2�����K�����������:.��$�~��:��WVV���ucc�Y__W���ה�u㦏&H����=	������0]��c<-�t���p�E��4������}�zq���y�	�}���4�o��7>~�OS�P\������ �����Ӕ����N��x�p}C�w�:X��'~��ӧ
����kR�$H�`�D�wH�	ca��z�W�O�?�m��`�7qr�����Q4��|�7a�9��H�߇�ԇ�F�������_��_�=���Mт����^x���������[x���o��q�Ew�px`0,�ǒ)��	ֹ�������X�B�`,�J�{!���7l�L����=�'N�p����|	�mc_	X���D�GPpИ�� ��B��yp���o����"� B��B0�������g�a����ˑmdM��p��ma�{����>�c�<i�~���E�Ν��{���t���ѣGfggg��)�΋z�S:z
����z�p]\�W��7���z*�b�Z��Qjσ>�%ɝd��'�x�/>��m�9s�{�-S���i�)d��t1AHT���%���/��T�x��ǧ�l����ޡ��&p$�W<��Hp��#��^��
̿0A�^Q�)�0�=���(]cx��$
�%�&�F=�y�H^�O�:�G�YS�p]��z&~���"���H`h����f֩m�y �"% �=�v��T�b3v���~�M8�~w~��~m|��*a\���^wŽ��ܔ;��S������⥔@DEJ ���wh���"oD7l���i���uB\��W��ס�z#l��x_=�bu8�t��B	���xii�Ob3�}��)���,�7Q��6n���~�q��j���`�Т�Q���{6��N,�&�RA(���&�E�j�`Rr����-�(��~���ބZ�A(���
���S�����_��8�%�"��l�����ST�ET�ADEJ���9�t:[��d Y.����_�;�ǈD<�����>	��ǎ�k^A(��?����7l�������SI�_U��\��w�)�'����U�w��K/�5/��� � S������~O+5�aʻ�T>o�9G�4`�x�a���a"z�b=���O~�����}V��BI���l��08`[	���3،����)��$�XA(z��zk�~S�%�|��8q�-k�P�;�6��"*�P(��)���Q!Y��'_L҄�ߓqѥ��6����<ōi �?
���=)iqWA(	�����i	ET40�r8�З�^���*��� ���Ge�6Û'C؊����賊z	9�DDE�ӟ�I�� a��}%\C2�W������^�0ADEJ0 Q�3��A�K�<�Z�8�L�����>�S)��� �g�8���"M��S�����h�U�'��\󒈨BI0U��^:z�d�3KK$c�XS�'����J(��� �D�ܭ���p8��t$J�G���S!������zBDEJ"2���$��F��F&$p$�d�6�G*�5pTF� ��	�7��� ���	A(	V��1ω2c|�miR|-�������^�G�P'iV,�RA(	��� �.h�'�aO%	��W��k�������m4�i�CK�JyDT�$I���Uf?\��p����5����'�Y��LӬ[<�jQ��@��2�Ƣ�׭d��SIDe'ɖ���|&z衇z�n7�]&��Nr�DTJ"�"%�1�� ��ǀ�l///��������_�z#�")�M�Q"%�WIDT�$(*8�9�8�L[����- ,"*8�	xq�t���R�����GDEJFn�S�ӭga�R�4)��C�k�@p7����<����u��� �=��:���ߦ�x��`�;vL�T4Гx��߽�j���į�i\�Z���B�x*�Q���g%M�U�\�$0I�d�Ae`��&ń���ADE�!� �f+6�˒��+++b��5]כ���<hc�ucJ(��� �=���>UD�����h�R�bg�p�5jVѤ����^*�"*�P�DT"�ER���&*��>�����W�~�z���-�F'L�R�[���8�J �"%AAi4!���M�)\��͌�O���S���o��T�����_R�RA(I���>*!��ˌSO��L쓡�k�qf���hZ�%�UA(	z*8�RxZ���-b��F��Y����c�{@��$"*�P(5��~2pLV�����k�j�K+�\�\�+\TL�
�SIƞ�&'�r�ŝԩ�GDEJ��tPTJ�}B^
V���"�}3A� �W��v����3�������?�^LD�$"*�P�f���C|jR\�τ�t�T�˨��y��������e���tH�P�1�)Y��#�"%���XI?�����p�&�C%��Zm%B�0y)<ܥ��#�b ޏ�JIDT�$�Vӱ�zo���
㠊pZ]���=�ܳ��	�yY�a��������<"*�P��&Y=����Z���@�\筴�_i�+� ��$)Z亗DDE* K����78z*XG��4v(S1R�3���

N8�'6WB)DT�$���YZZ��@M�P�'��x*���鑧R�ӣ橈�T��� �d49G�q�s_����!"�����{ �%X���
f1Ї�!��@<7}�~Bcا�JIDT�$�n��R��MؙQ�/�gȒ�����<� �SD%�n�����wm�ƈ�c���c��|�Q_A��+^���кZ�S�TRh�ۣN���8\L�ښ�;���Z��Gļ$"*�PzE��3�qB�'�"	Jޘ�E�TRHDw K��A����Epy��r�&��3����DDE*�W�S�/7r|��M���h%f	ä��B�O����uF�f���QT�����vDTJ"�"@�,c��8�7��H�i�׍:%��.-�����7���=u���/>��H�[c�c󒈨BI0��J:�q��>8������mO����)�v���e�k�_g���ē4?i��W�E���l��#�J!� ���ѣ8�S�M�ш!p5pBC���;7�[Au)hаY,z7�����h6[�n� �1p�]L*��Ebii)��x�X�r^Y��}8��V�O���v�����3J(�<��P`�B4N�N��K�$*h�h�R1B�e4p�� �<v�6OV7�x��nI	Vn��hee%P������^g�B�B�ɣA?r��J,B��z�
°�onNߓR�Q���x  -,%SF,A�@���y<���^h�P`vww�uϜ9����q,��/�7 �h��������j,�<�Eb�[~!x�Q�z�^|N�8�F�~��)��@DEJ�a[F�E�K�8������lmm���	<��~���2����kp��:�v��8	o�^y)��uG�S+1���~�^��:����!�5/��� ��ȑ#0Z+I%�$>�g��8���S�P�C�˰���M��?���Yv�v��V�B�b�b�ך�r���u�z+���	�1�����^�=X�fw4ZVB)DT�$  ��a����S�E��ӄF�ҍ�o�<�}�c7o�]~K	��v:m��]q�
�D�(4I�B;QXp�M8�*�4�.��� �J��j��"O?qb@��Q�S�Pop*]�o������cJ0�v�8��$�|<�g=�Z��w���u=�O	�Q����`�:�#�3�Ә���Il�wTjE	FB�s�z9��D��zOz��]g�\7WM�>轐��� T���Bﱍ�ϔl����]%i���
)�h=>���,����Ҥ�$"*�P��Z魺x�KO�ν
��VJ�m)���uc�:-5�ʏ���'�,��y��`����C��?�a �½IE�x) �"@������Љ��`��X`�PЅi*�"*�P�؀֭�ж:a�;�a�EH7ځ��T�������(�^��P��)18.
��	&�3��}8q��PA(���&X�5N���*�k��
<�A�S)��� �$ZQ��F��$���Z)�(�L_���ղE���SS5�y4lC�p���F�:�ׯ�9fM���ݻ|��!�*%Q�
)"(�6�vP)�H�#�i��r���b㺮�S)��� �����sݸ����U"2N��T@��)���J`"Io������iq��s��T�`F���K�|U��� �v
��rE��"*��_1���q۹���4vCQ����BIp�.����itG��>Y��pO�O�N������UgM-���T�Յ��xy�֘�f[��/���X����p��j�1��}�OHܕ҈�BI�á�y�L�=���dØJ0��w*U�u�4.{=��i;=}�PA(	x����A���DD��i����8+�h�{�
�.xu]p@��c<6=x$.\��h2�@�/�M4�cEM�V&�WD�ZDT�$�n�FQv�!S4���)�E��M�0�'gJ��FR
|����dr$�X"*�P�����퉨�u%zh�D����J}2�M	Y	��$�Ҹ�:�H��ՍZq�/��7���5T�lĭ��K�b���%��x{�TphI�RA(	f˵�N���ݛ����Ux�9������x����w�xM'����8��x��xܠ�&e��$����A�⭔DDEJ�)������T�bc��]Z� ���A�(����Ӫ�4�wܳ�����AP<5h��Z�-���k{��+����9O�?�\����B5�,>�5)����Ɔ�aa芁��M��#�P�u���;�jkkK��NB���j|��j��߈=����xp5�%ޏ��Fӥ��Q������i���$���n*�o���?	�4��p�8Zmpq'���wc��o�Y�j�5`��0��7�!�;��N�;�������q8VֺC�{����)��psH#F�o�������:�>�^s.�����/���,�RA(	��p#>���QL������!PB���?"g/�������8�=���#C��Xpw���&[��&<zH�>,|<{�M(�RA� �1
��P5_9�f���aY��0�.��N2�#�
�M�[��q,���{����tI�b��E���7L%���:+ԆX?WI��DT�A։<O��,"*�P،�J�h�PP0^���x�'�����oR0���ԏ���9P���f3\GcSoz[���˞��P�R	"*�Pl��a��ǽ"_�á
��j7�����KR����S�Z�T�	"2�OJ�N{b�h�:c�T,,��t}'n���_�3ȵ!4|:�<N��C��*��� ���&	'�����L͌�O��G�^�Ȥ�F�0������J;�6l˯�@�>�FDEJ₧FK�g��� 
M��ɘ���-���T:v��Si;�x
��
RR�G
E鲰�:���)*x��hDɔ�xr]c/g�u.���;�TԗEDE��� J���0���Ҹ�#�1)@�>"S���,�㋨�EDEJ�M�M/��ߏ��SJ5�-|i���m�T4T�3���K��qu?�J��U�Q �b�r��v��q3m����=���]��+���6��w{���/M�S)��� ����S�M�y3Q8�l4zRQo�,�w������c�i4�IqYDT�$�7�br+T^ %a?.{�/W�඀@�K��`��H��
��qR����G�F��AG�[8w�\�ۿ���y3n��D
;N�K��4"*�P��8��T{���Qx���L(|���q�nK9A�R��$"*�P���;���'ؾ���HɄ�qRq��3)9�X4�ɍ��t1w&��p��q��?~\D�N(g��<�����|r�w��%z�HIȱ$"*�P�F��u��n��M!׉���s��l3��c��J�0�|�m縻��#�#J"�"%	� �D^�F-��6L��O#p;�0Up2�L\���\_�<X�C��*M(I��8�#����]~����f��$�W�>�5��M�1��%Q���A�Qۗ�˖�ʰ�5�츹�R�XW�_��#����􌟂@��Cϓ�WIDT�$(*M^�����'N����+�T�+7�+���\��k��qծ;PQ��j�
�=X�%��Ɨ�F��0�koXfZ�.���ל�X��7�Sa�am��e>�e�^�-����BIZ���D�E��"B�����İ����p]+=nR�='�p3r�W��ʎ�o,5��_��9f�������}^c��G<�}r���^�[w�)�#J"�"%9w���O���+�64R��p�X!���4ף�07X�u^RcM	�|��߾�_X�/p�g�:�N�eo���W�C�qM�O�:N�����=�8�$"*�P��>��g���k�Ap��{�^��6�e(�G�L�W�=�F�:���`0�!ع��{�O|�O-wW6����.%�v�ƐX�-��$�eDҲ=�b/qy�ۡ�����XA��m�N�O��J�},5���dP�$��z�7G�u�������e�E�o\��w���z8����]�j)|����-��{��dML��D�c��8ts<HZ��D�G���{�PA����]��o��o�xl�]`����}�/��K�h�p��v�O=��ã��JH�W��?�_��#���[��}O�2f~���gn�yx헖��~k�=۹|^	eQ�
���W��g?�S'�������onm���Vl��*����h䰂ǩ�)\>��+o\>%͉����g��'���3w��rd��}譨DН�%XH��%b��WVV�ɥ;�O��_�}��ux@*�+@DE*"�����8��u|i�B��^om"����(��j��7ܠn=����F�O��xK	��:��녧�;���Ou��b1�DA!q�*��;0酪�ݮ:v��:~�?����ֿ����e%T��� T�����o~���++�a^�Z�����2���ʩ�+��v~�o�����L�?~���/�o9�ԫ����dL�7�c�k�h6�ɓ'ն��O�������BDEf f�ϳ���������P��L	���������9��F���
tEB��"�"3`�����l[��.�����eO����QQ��%-�$֫��;�j���4�t9]+"*�0V��OD�~�u�[i6[-��W�vC5�YIVx��H��e�UB����hu�`��J��ႅ뉨���V��^�#�L�����T�+��Vm%T���_�T�v�    IEND�B`�PK
     uK\�4%2P  P  /   images/c7b8e0ca-67ed-4237-9266-7527aa3ce92a.png�PNG

   IHDR   d   e   ��F�   	pHYs  �  ��+  IDATx��]	�Օ>Uo�~����K�o�DTH�d�LΘ�I��/1�Jt���gƉ_2ctBb �� Q@�UZ�l�fm�����K՜s_��v������$ݟ��U�n�{�{�v��§�wE��=���O�UU��r��(`�Z�A�8I��u�$�2�F�E"���ba��7�Og:x^<=]��t��:�Fy�i)o~��7]]�� �
�����v��x�	عs'<��SI��Y�`477�ѣG!�
�����#�<���s��Ҫ��4BJ���x�
&S0���k2^ch"T� ��5��O	k�跂�bi)/�N��t��N�SIOO���|u�С�1c���X�`�|�Q���0��l���������Y�X�����o�}pҤI�v��ﴴ4Kkk�",��/_>P��¤v�2�	=�1�@��1P�4O����݊���ԞW���^���|��=�CH�5z�:}�� 2؇����� m���:Lw �э7�Lƍ�@����c� 2w�\=z4c*ugaq[[ۓx�K����DI����E�ō>����g�!�� �B[�lك��뿅�����L��D��7�������رc�r8��C��dI��XL�$^��4�{�KO�:!�#�PZ<���������K�^RXXEEE�W`r�{�&55�V��]J����x���� ���<t�2�=����&݂|��\+��⫨{ډO=QҀ2�@gg'R������\�%B�5�-��+*�9�[L�G��(�P5�́�z+)qQ,��-545L��-�{�/���)���p����%H{{;3g=O�d#*����D*�-i @le��q�5 B���WB`s���*3�
I��X&:�h�����"@T?�����˿��W����}_Ҁ�]�x�b���~:33s�}����ZU�Hl�I��
_���0jD)({�%E�P�}��� �SY��+�$1�^��A� ��رc�"󺱱�0Ϥ Y�p!SN����Ì��nL��V�Wu`,0k�l�V9:�PQ�Y��6�ɖ�06"�l�7R��E�xo�u��p��w�h�z��]��GR�ضmL�<Pg�Cg'�X*$����;���_��wv��Nb�
��m��S �++��(�>8r��)����hi���O�d�"�Q�dUTTa���/��e�b�M
rvHN�2�Ez$Q��L�� C�-��h���f��d� Y�ദ��7-�E�̀�]�? CF��o�N��s?��X�� ae��0���x�0]R�4551Ge�d1��H��K�#��7.�<L��g!+#��\�:�75�_7n��l�@�|�̡v��]�#'�Կ@텩�HD"� (o����cK�� !{z���2���D1뭛%�X���!=�>,��˖�˾
)+��翀S�k�d]��8ʇU��a��W!�HПaonc���Xz�i�*GII	�2��D���O��������>f��i�&Xr�B�"65%��`����;n�/}�K �[a��#�|m ���O��f>R�ڵk%�Gńi@(�Q�F�����>=�g�UӟD =[� �����wv�G�����K��}UU��/,��Kn��<�
ܾ X�y���#��!��3sss�H��"Ӏ�8��]��ٕ�3'�Y���&�������0�rL�>>�9�_�F�`�FQ{�Ԡ�咼��C�O�Z�/Z�Y�D���f��4 �?�<̟?�l�b[�^X�O"����,<���PV6�����}�/�e^:�%2�áxn��(�����X�2�o� IA����yLr�u�1�
{Q���m���ުUUw[3Դ\�0z��VX�1X�W�`,x�hkb���ʥ�ȷ�:E�Ӊ��w���W�1��녬�,�	ŉ�+J�C$}C��#��ρ@�7���r_'A�C�迕��?��1ә�����L3I/��{トq��HT~�X�!0l�0���V%�!��@�x<ׂ9 �nw`�dl�1�x�K��@���'�r!���Ǽo����%��l�P�K��|�[CJ�!ŕ��x���f��9A�\7�J[c�
�s�|:�.�ۛ���GF)n��:��c&]�(4n"E=�+yji�U
S����a4���χcǎ�L�����ʓ&M*L�x��=Q(���u7̝>�y�	�,?��1y<��cp����~"�3Ӯ[ ˿r'x����p�B����)�*ZV�T$�0�{>�-K�3YXf4م8�8&U"A4�H�E�f�V<���_�n=�"ӀhÐv��zbtoM^��U;w�ޝ����jH�o���
#
� +�.����Ul����>c
��7@qq�=N׽
*�R4��33����@*'T�����탼�a0~�h4��C��#([�`��a�*����y�PQ^
�O�Bm�I����K�r�J���RKJJ�1�l�I��#3�H$}oL^��U�ߋ�a�Ca�(*̆��UPWW��{�A��fB��߽�Gx��`��ɰy�c�(()�k���;vCi�X�6i,�ݳN�k����CyQ<��'a��j���&X�����C�ѱ30��E��.�s�>�X�E"�dz�:�"'���B��u����J'j�&K���nA`Eŗ��2x���/~�K�D�n�����|T�Ϟ;�� vW��w��� ?'.��Aͱ����B�K�?��8sG���Z����3�@]C;|�_��F�����ǵ(��B��:x�~'?i��>�i��P��a�U��N�6���)� S�<���,���f��Szq�Hr&�!�I!����Z�����gVAͩ��p�PEGU-V��r�`��	p��0c��d|P^:�����M�ܨ���x������`���EW =���c���`�ֻ��Z�$
4\�$�sr� ���	���](��322.�Jg
��+Wo�Iʱ �7gOL��؇�����spì)��'���OA���`Q����U�Z@!T�&OG��Mm>�Nw��S�P^<�N��?<xŗ�i��#�QQ"uii�N�s�Q�qFc�h0O�c�8����bd�����}�~A��Y
�!������5�?Q�̄��n�����^[[w�C?-$2Ym)�����w`��_g�rz>,�?&��p9!����dI]�Cm��l�n�J�l(�d��;��3'����a>���:��b
�s��AAAU&�q��:�4�j�-�@NfdN���f�)5 �ۃ�E��@��g��LF+���ZRi�(PVZ
C��`��yP�DQ� ���a�!�t�� dd�@��0jx9���������	�rL�9��g7̻�&8�ql���*'Cr��q5dS��C���\�D���o���oFq�M~#�M�����?��5�E��N�S?�!��>����W�D������Qѡ�*�?�$X�4����>
�=�(j��C!صc�z�F�����!gO���x�up��hmkӢ��I]��{���h�"�������g��89j�;sߩ��N>���(!�O��h:�0������]2S�x���s,��^6!�X%hhĿ��B��Ψ�ol����~�'6'�V��d"�Tlh|R�k���CƜ9��~�v�e�O�٦���>:~�ő���SH��b
!��ǋ���Y�q�ar���h:	x��:lѨ�$<&ws�l�KY�5�]0|h�'�!��ʇ���Љ�e��s�w�����X�5��A��^�Ƿ�� �S����Ǎ�O.|���=)��N���BlmKʔZ ��4��{�S���*���t�|`����VdQ�nY��W�w��zZ(�]i�j�.��C<��V���l���ܯ����9���CQʅC����uY��e6�5�M��̌Y��C
' 4FBgq�?�i�=�"nO�2���n���Z�h�`��4��t�_ƕw�����p�tqZ�5|��g+�L���P��.�`uyʈ �2�����9̯�5���6�3�Z}��p5h�ւĢX�b�_|o��{z_,�AaZYY�+�Xs�"����?.�u�������
�P \N;���&�DL�ݎO�C��f��h�'Q���x+�����M܎���(�鱘��).I׍����\<H��^�Ik(�?������}����I�j`G��h�АcNG�K�C��ⓦ���X���W"$�¾)4����>#�l"--����$�0*�u䞭hZa��r⵿�Ѐ �%#����K�8�K��h��#���B��%���
k\ŨLF�2�Fe0�=Y��}-�N+��u)D>u�3 �o�P(��ٟ����VQ�'������ ��\,�o�Z��iW�$�F=)�\|c�bK��[�5)��[�x捕|�����"�*������x����(���|\_Й2�J^[�<�,"V�*13VK�I)�3��b�d��������%υL�Q�ֹ7�0Pq�ٳ� �Gv�,K�1�&d�d�xZt�i]���0��r&wt���X�D*�쳱�&���O������U�-�c��1<w�փ�a��A~F��-U	~�o�>�7t����q}�����z��F`hS[.����� S�ՇٱAG�A��xf=R]�~̬��Y�FßwU���(-)���|=��>��{��.�A)4*���|�X��{"^OR��zӶ(�CFz�K��=z�"�����7-cC=b���f�i�wU�A �s�@$�!�`0��Bѓ�𻶬��b�D�B�?�`�*tQ/$�{�!14D�Wǲ�:�d<��!V�v���fꕙ^���q��u�Hh,e)���FJ�Ha�
��e��wbYx#�[[��FE$q�L�:����H��!�G��v{�e��≶�x���G9���'R��h��{���y<�&��n�w��&ca�(#?B++��92�)p��t蘋�-@dts,V|^��i�D�L�:9������F���O�>�-�� ���9�<ۏi��F�И�[���^�:���x;��,̸+&- #i=��I�k!�س⳶��4�5�1����A��V���!a��V~�ػ��9�s(=9�?��e�F�RpU4c��4��=X�'��{��k9rdW4N�CO� Y�jˈ����+�[/�N��g}:���'V�*����'
2�+T�Y=������kF!�X���
��&�hm?�GtѢE����,�)@.]�Ď�����n��n�������C/牌�q�� �h$&s�Jcn��C�E?����+)ߤ���ύ��k#cH��{�B"�Mo��alڷQ��̷���߀�^z)�z@x0+ߚ�N�;��D)V 1�I��M:靉�A4` �������u4�����J,����Pd��hy��̀d����n"%i��9��!}��!A��<fGL ��	&0���F=9�}Eq|�H�B��5�b*�ꉢ�͇C{"�$�OPLn£�]/u4` !��B�R�L�o@�D�C�c�2��3c;U�G/m,G�?�:����s�\����i@�Q�P���=���!H�gΜ�UVV��s��H0P���U��2����z(�i�&Sy(@4]@5�}"6���)�>��s��Aӫ� Z��5�[ S��L�I��~���G{2K� �cѦ%12
�\+�*N �M񬌌���wр��>���iׂ��!��>d�ԩ,�((@���Z�E�f��kIZ4D����� ��Q�d��lN�^����K4
�<�Ç��s@Bu:�T�n�p]�+�+���!�Qz�Um�D���((@h0����_[[�ί%2D��PnoH����f�9@fh@Ba���ׇƍ�)��%bU%:���>��<��?Z[[��&���D34� �/�M�8����C�|N�~l�~�cF��8w��|�?���uM9"=��״��4��(@HkKª����a��EӍ��o2H?*��xH��g��tN:�٪ �蚂����i(���R|��O� �c������&�a� �<���юy��w�}7TUU%\���2�ټ��W�6d�L��(���z�G�V��!QA����t����ފ�I��-	 �H��U����Q��}��K�����4�y���޻}۶ml����Huuuh�̙����>,y-����#CȤ� ~Z�)2� �4�WSGQW}�ҥ��y�hy�?<�I���|��Y�<`�L��Y��P��׼v��pIII�����3�ZBz͚5��8� 9y�d��+V���{�8>q�f�PSo����Ғ%K����`"�ZCP�q0�{Æ�4� 1�իW3eOk���y�m����7;�-��[tͬ�l�ô�hP B�>}:1���(زUa�3U8�Y���c=�$����dhP B"d���,���&}P�D_Co���e|�*���fP�E��g�4( !Җ���-�a����7�ڻ'��	�2�G��)|E��q��A�td<��X��0��d!�<p����[���ؾ�A���UAA?����W��!�;4o�1�,D�_�S���/ �z	����UQQ�|�rR��G��g�5a� ���M���A��z�B)ݬ!� ��3'�52g�ʻ��������H��0@�Wp8wڸcH�Z`J��)�q뭷������ny#�a|g�/�[ �~]�{b%H��m�ݚT���;３ �666RS&����`�g�قA��P�h� B��$teZI�ɢ�X�nw��+\h�z6l0:!�S"��OT�U�L_��m��4�mڴ���u}R�A��\���VT�,"K��ԩSMMMe���Ǔͻ �^�ZXXh),(`��v�ǎK��А�����W�4���_�6��t-��6Z}m�͗��x�:oP"�����*��"K�>�*�E;���2��t������[�*�Ht�sEۦ� �-VD���7h �(���mNf0*�H��k�D��h��vf��*�Ȫ��P)�Ac�SO�*�d+Ȗ�EePD����ݩ�8SS�� b�m�@	�T��ɝ#��YP {�H��	���-�bCP}5;�
��t���ʎ4ER�����Qa��R�A�(�t�[\0�f������"�ݗ� N�r2�j�Pc(�� ����0r��p�X(,�D��P��E+}� a�Qjɟ:�Wۆ�bW��N��wK
�VBR��T�CM�y��m� ŧ�� �ޮ-�`:E���ArT���5
���Ƌ�XXu�6���mI:�0��6%�Q>�}3T��W�*�@>���"�6W����g[¡H�M�~�3��ַ�v�/mͯ���+;`�]�7���;>�����>D���/.�Q��/W�Y= R4U���(x ��[�*v�0=�/��c��&�����>��g+O�����q��ˡ���?]�z�2�ܚ��4h �N�:v��8n�WO�x�jQ����ٛfo>_[�[�+[m#�u�4H)��Ҟ�v�D����s�L�G�?�K������"
8�i    IEND�B`�PK
     uK\�|��*  *  /   images/fe816bc3-a1ac-4496-aca2-7e46c72bb630.png�PNG

   IHDR  �  �   ynN+   	pHYs  �  ��+   %tEXtdate:create 2025-05-07T18:50:54+00:00��P�   %tEXtdate:modify 2025-05-07T18:50:54+00:00���o   (tEXtdate:timestamp 2025-05-07T18:51:13+00:00���  FIDATx���{���}����{��j8��X���x��$�c�gNc�D�$�$ 5�ͥM4st��L4�K��1Qm"�h5��`�**�u�%ފ.�%�m����Ӫa������f���Of�^���g�����_ �(����?��K�,yꩧ
@����8�]�z�a�V�v�뮻������?�S�����=_��WN9�R�*�ĉ�M�V ji޼y��z�g�y�-���Q��)��ߔ)S:::���T��������N�Z �t�M�'�|��eԥ�_�җ
@�f�}��j�P��/Z����/ 9�Ν�t��8��5ԥ� ���?��e��� ����?��W��Z т�]���M#F��v
�J�R)8@*H�� �R>~��aÆ��g���6m*9R>s����ۯ l?ͭ��ŋK�Ԃoذ� lW}}}%Jj�����vw��Ԃ�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
��'�\�jՀ�8��ÇV�ZR�H�7o�<y�_��_���w����.:��sP?
�����[0h�ʕ���g�:aԌ��뮻Z��������N�y�P'
������Z<��^[�h�����ԉ��1bD�<� 5��y���
���Rp�T
�J�R)8@*�<7n���~����v�a�4
an���K/��^ؾ����>6u�ԝvک�C�!�����N�<y �|�]w���s��)�Pp��aÆ��;o���裏�q��GT��c͚5˖-�����Qp��h4������nĨQ�
9 ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � U-
�h�b oM{W���-�[�l���kkkk�
:::6n�X �t�)��KO���7�<��wl-xOO�/~�իW7�nooo�JƎ�dɒ��ʋ�-ϵ|��[�)�㓍�{�ܹ/���N;��܀�MT��+٦ ���/}�����~�<�˖-k�w�e���R�оM���LX)Mߥ4��<xpU��m�/����ֿ{	�o�!� �\��J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� ����===�4�_����Ϻu�
 Q�V�z��߭� qC����. ��N&@*H�� � UcӦM�* �i����V�* �i�;��g�1bD Jc�ƍ����4��H�� � ���Rp�T
1������t���dQp����6�#|�t�cƌ�Ї>4k֬�1aB�7�x�A�iӦ�8�����?��C�!�>��p���.����ێ��c�=>���~�ӟ.DQp����z�6l؎����*Rp���45:;;]?���nݺ�C� �4-Zt�1ǬX�� e�y����@�F{{��$r-
@*��ꫯ�~��͛P3
��N�2eJ+'�1bܸq��FwwwGGG!�g�q��>��#-�x�UW����ưaü@�3k֬I�&�����@=z�^x�Yg�~�Ǐ���R����5}��f[W�Z5���8∑#G���^M8�w�`��ߦ ���|7#^ H�Z�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H����mkk+ �i4���gȐ!����m����{/_���ooo/�l���/������7m�4k֬����_����?~�����{�7v��������;�|��>��Ço>�[�o>y4_x��{�{�g���<���U����9mڴ�mmm����G����}��{�g���okF˖��m�6wöw2��g�f��;�m���tvv2��[����{�7�|��/����Ts���w������n�4i҉'���ުA]�sd��[_^-�:��ע�M�Ug%�j�7��[��}�������z��os��_p���G�/F�I�}�����wZ>�����Z��p5aU��5�f�~��_~���a���?��ѣG�}�ٗ]vY�7�mHi�"_��ӮE:{{{�w~��s�=w��7b͚5��y�=�\z�'�tR��Z�O���(8����4�ޭ��|�8���<��k��fĈ�J���e˖}�#Y�hQ��N�2��?����_�)��%��f̘��|旿�e%ӗ/_~ꩧ6w����ԏ�S_�]�I��^E���0w���o��@�(85u�-��u�Y��O�^�]S�N�:�:uj}���f���ھ�����v�M�v�g��i���Ə�C(8���SOM�8��խ��z�1�|�S�*P
N�w�q��&L�0~��#�8�@����'>��/��;�3�}��USp�b�̙o\�Q������/���F�J)8u1y����+��0aX�:
N-|�K_��/߶I�&=��#���T�W^�ꪫJ�9s��v�m���'TD��ޥ�^z��o~�
N������4w�%�{�1WR�b3f�X�vm����}m�̙���T,����u�ֹ�Pp���+���G?*ɺ��򓟜v�iZN��Rs��%u���
N%�*�}��%������>�@k)8�iV�(��l���3�z�ZK����ի׬YSv���WpZO����ٳˎb�ܹ~���Sp*���]v>l�J(8�y��ʎ��_޼y�������S��m�7̛7o�ڵcƌ)�B
Ne�Zv���ZK��L[[[�Q�H�/Qp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp*�~����ؼysooo��Rp*�w���(�nS����\x�3g�,;�.�`�ȑZK��̻���+������/�N<�ċ.��@�)8U��|�	'�|�ͯ��j����}��O.P�b�z���__��N�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�S���M�6m���:娣���?X�ZR�HO<��i����3ϴ`��?���o�� ���y���c�=v�ڵ�7}��1c�\}����s�׶,�o��k>�����^�ϳx���]�l��C�(x��#G�~hWWWjF�R)8@*H�� � ���Rp�����{���{��I�\3G�!̧>���n�m����/��~�����C�!�7��́�wӊ+>�������,�Pp��v�ڋ/�x���~��뮻�/��/
!b���k6l�O?�t!��C�A�������܈#Fr(8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@�Z|Ȑ! Nc����W�W����okkk�
���V�ZU ��j^�0����}��-�O�Z�W_}uѢE�_۶i�J��{o7W"�����'��k���Q76m�4w��-[�>�TaРA��� NǶU�~ea��g�mF|�ȑ����#Jcݺu�-�|��/��@ �H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8��������6l(�Pp����5�#F�Uȡ�c����gv�u�܈�}�s�
I���y��=��#q�;�$Qȡ��dȐ!?��-��r��wo�Î;�����X����g�6��z
�J�R)8@*H�� � ������i�����Ԍ��ٲeK�vtt�f<�ĉo���VN���=��Ԍ��y�{�;�o��L�6���� 5������op�7�p�ʕ+tБGy��~���Ou�6�����N6lX�J��),�6Sp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� ����mmm�4�����!C���� R�����������݃qҭZ�j��6m��O�����������9��vۭ@��R�Kc�]w?~�ҥK7n��|����ʖ-[���
�]�-z��fϞ����lŊ�G���w^w�u�_�����c�~�����G>�<���ӳ5�eC�{����_��͎/_���giF����y�m�xV�^=u��{���~KpÆOo������?��#?�я�x��ƍ+��OyX٫�s����*�s֯�E�y�R��V�����t7w����w�-�͏��6͔�s�9��~���[�Mz��e��������j�-[�x/^��o}�;���@��m�>��n�a����[���v~-
o�W\q�����<蠃�������F�O*���?� .<��sz衖M�ꪫ���f�I�L���;����Oo�ܥK�w�q_����������ڟ����_�U���k�{�[n�eԨQjF���I�&M�2��U���,�7o��S7
NM�$�ox������8u�����ɓ��74#����wΜ9��K�zPpj�sι��K�<��SG}�ԃ�S/�������o������|����Ԁ�S#+W�<�3J�5�`����M�8�@��I���>��SN�&�Sp��K.Y�tiI���}�i�͚5�@��ZX�j�e�]Vr���w�}�I'�T�:
N-L�0����D9��?��:�@E��-X���?�qI��K/]~��\rI��(8���W�Z2�t�M
N����Y��?�aɴr��3f��
HvT
NŦN����]b]y�
NU���y�%�c�=���Ͽ��,�r
N��}��y��p��{�y�W���*͘1��>}�9����Q���*���?-�z���׏9�@k)8�Y�nݣ�>Zv.|���_����<�쳯��z�!<���
N�)8��={v�Q�0/&Ȣ�TfG:q�~��-��TfΜ9eG�x��fć^����̟?��(�~��_��W
N�)8�1bD�Q<���V�H�� � ���Rp�T
�J�Rբ�c��Z x����^zlSoO�hyӇ4[���t5@�l���O~qޕ���/m����Ne������|�+G�:�lXYF�����^ �e���[�8ѭ��e�q��w�7��Z����
��k<�ʒ2xԯ�@��΃�/+ ��Մ �
�J�R)8@*H�� � ���Rp�T
�J�R)8�Y�v��T�͛7���h-�2�~��9;����sϑ#Gh-�2�\r�7�Pv�^{mWWW��Rp*�뮻>�������.]Zb��N^xᩧ�Z���*u�QK�,���;_{����ǌS�

N�N;��u
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�4hPqo�@���ח�C i���9���z ��� ������ �؃�Rp�T
��Qz�K{[ M�t����@�Fy����@�F�h+�}�͉�0���/� �\��J�R)8@*H�� � ���Rp�T
�J�R)8@*H����7��F{ J��x��=��jK Jc���� q���]� y' ���Rp�T
��Q6n,���l( Di��?�^�zu)��(����{�ҟ�Qc Q}�0��H�� � ���Rp�T
�J�R)8@*H�� � ���Rp�T
�J�R)8@*H�� � ���J-�^{�U ��δ۾�����=zt�~���%����sO��Zp  ���Rp�T
�J�ަ���j����-�� �uttT��Ʀ���߳-���,�9���� ��c�9��4&�����ܬ2l�ʖЬw�@�1c�T��������|��{�N{���R�Z���˸���Z�� �1b�GQ�m�s��F<���75��>��Kh���i��z��ާ@�ɓ':��5l�eH[�e�u�A�{��������/��S^:b��_}��P{��˥�^Z�*��Մ���F���}�1����:��
@�͜9�����U��z�c�=�G?��E]4o޼PK������o��C)5P��7�����~��w/Y�� �Ƹq�N>����6�U�7|b������Pp�T
�J�R)8@*H�� � ���Rp�T
�J�R�_.4����I    IEND�B`�PK
     uK\�|3�  �  /   images/559c8cb2-c573-4147-bde4-a0b817dc20ed.png�PNG

   IHDR   d   �   �|�W   	pHYs  �  ��+   %tEXtdate:create 2025-05-07T18:50:54+00:00��P�   %tEXtdate:modify 2025-05-07T18:50:54+00:00���o   (tEXtdate:timestamp 2025-05-07T18:51:13+00:00���  �IDATx��OhY�����[Y{Pt]ť-(붦t��vY���Ez��R�Ų��*
b�Td� �����R�Q[)
�V��t1����Mf�gf�	b&���vf:������k�̯�}3���{LUU��ٳg�O����
 ~����>�O/�۠(���Ǉ����x��i}}��ݻ�nՕ%����,���hY�N�\��g��[SS�� �G*IROOO8�_EQ�˩++�C��&	�K(���IY90$+�B^�5�8ѥ0$��*�"��,$�B@��,$�B@��,$�Y���`WW�,˩^V~��?777WUU�31KVoooGG�6]�3g΀31K�e�����z�x�6l(--5�,�dY�������=***�%rS�����n3�rv��F��޽���靜���&�lY�ؒ)�V�ކyV�A�	�$I����%�؊�@"������t�ņ�����zĿ�@�D� ��wnY{6Y,+��5�%�� o%$�B@��,$�B@��,$Kv�a �Y�ӫ���߼�%g�,��U\\��XRRbRqΖ%��[����R����xMM�Iř���/�`��%�U�<�����Y���]�v�c1+����>���I��Bp,�ƬT(���-�d! YH���d! YH������5Z�uY�7mڴs�N�F�.��mh���M��r$IRQQXH 8{�l?7�L���hii9z�����D�퀺�Y�g���$��
�q9^�_v._�|�ĉ�NΉ�	������;w�_�ޢ])���e٢��|�����رcz[?~|����d+�F��q�?���̜<y2w�����W��>�����߿����%�]�~�����0�����~��lo޼�!l���`�˚��6�-�~����e9���d! Y�e������u�ԩ���ܯr�۠�k�z<��e�� �����B@��,$�B@��,$�B@��,$�B@��,$�B@��,$�B@��,$�B@��,$�B@��,$�B@��,$�B@��,$�Y�FGG}>_$I_ŋ��ֶg�p&f����զ��Ց�L�f�[���^�z�>O��(��Օ��`ΎY\��Ç_�x��������gFqΖ��%)s���g˂lol�7+��,+'�YY��l���YmM�dY�
��>��!��2�
�����h'P�u�'j��+fn�� e��ene�i^�=����:�@ٮ|ୄd! YH���d! YH���d! YH����#-�
[)�-��voٲe||<53�,˛7o6�8g��ܾ};���TUݸq�Ie�%KoE�e_��`	f�jhhhmm�"��?755�c1K%����_8>fY	�B@��,$�B@��,$�[����V*d[XXYY�$Iڅ�2�˶����'O����&{Z���m�f�>���VCf]Q�,���x�^��p8l��IW�\�p�����S)|���w����[�Z�����ӎ���@�+�1�jo�G��y�fFz$�{�n x�����fg@,(�e���;::��R��������u��Y�;�=n���/w����s��]�xl�~Y����BKf���}͚5`��4��Ç��&�?�,��F�)�2??��e��xD�Z�(
��l�u��s��Â�/������z@�+S�i��fFTm��	�
�Y�v
+ݒ�FH�r�hM�2��m�]��l�u묬Z�
l�~Y���/_���^�S�
˺;�U� �����Aw�!a1��_C�Ȕq(f! YH�ÊA��c0�Uơ�������=���K�2-..���y�D\.��ϟ��g���~�ҥk׮��;T�Z�I��d%
�f�A n:I~%��@o�4��m"4-
�ףl�f?)�Sf�Z������bd-�����?���鯔�7<l�ر���J/C� ���t�޽@�]g!�@��OP��    IEND�B`�PK
     uK\ә�CJK  JK  /   images/a0bdb5a7-9945-4126-87cb-dac9f24142ab.png�PNG

   IHDR    �   
���   	pHYs  �  ��+  J�IDATx���T�y��LhS���C��P�(���"�Ԩ�4��hR��qe�(U�$��j[���(%FLI��(�<�- ���)!��o_�s��2sff����[k��9�59������FFQ���RQ���RQ���RQ���TV�Z�ۼi����oEI7_��M�֭M��=3��o
V*[�l�-Z��,_��|��'��>3����O�?�k׮5/��R�m�v��;�r)X�`���0���C.�3��ٳg���
R*�֮�-]��(�&�L��}�q��\۶m?�Z)H��۷�|��GFQ�p���Oͦ�'��Q�R�\�(J�`��~����wRV�`
	ДU���Q�d2���*��Q���d���)�������t�G~Hd��f�g�ʿ)���5�_�����C�U&v��\��)�R��̗��%�g�g�Q�F�
E��"J��?4}�����?��?7�'b2F� Z�ɧ�ڿ��W�U>��+Z���?6�r�QG��=z�V�Z�ώ
��V�\i���ڵ[7ӹ�$#��={vn����o�g���U����g�ɕ#S�d�"�k�+Ń2��S9�d*&=������r)�JY}*��%�]���%�'���CR.iHYQ���J�R���F�J { ���)���Q��U*Q&��QJY����(�_|1WSS��p�e_�fMm~��ϼ/\��L�:5���d�\�l�)>���A�ՍzR�ڵ��߿���+�M�6�n��&C��-��cy�f��fРA��GFO>��m����ɐ�3�<Ӝp�	v�!�iӦ�w�y'��(��/����U\��`,X���hK';�R�c��_5ݺu�ra��{�n[bNF�*��e���������bK��.W��;v،m`��Aŕ
7�I�=/?<C�*r@:t��;J��rB},�����l�2*���={��o�=�GqQ����J����z���4o��>D�[*����)Y}�+_1͚5�&�*��q�e�Zse���\!�JE����Ʈ���R��{��q��f�ر4��4}�t��k�َ{J2������'�-ZDQ���~�̝;����5�|�1��u���T\�'#��]F)|UX�n�,@� `p�lL�;7zQ*қ<y�=�jF-,n^�n1�W\a���jk�K?�pD���[
���:�k�v�rI~���9s�x�no�~T���9��E2|�p��s��~�+��o�H�`�"�گ_�H�>���B~|�wM��g��0�x���S���DuCʻv�2��[@�a�ࠬ?���h�!ם;w�5��?�E���k�<z���7�
q�F�#aO9�K_U�������my�{(p�����T�����Ew��]��;��r�駛>}���Undm�8ڷo��Q���'�D��T}�Q[��o���I�J�]����m��*�í�P�Y�������n�8$��{�vW�$���̚5K��J G�	LӦM�gd��O��_=��j(���c�=�h�E-����y�4i�Ĵi�Ɔ���S"WB�$����L֠�2)O��
����O�*�1�ͩ9����رct��н{w�@��f���(D��T���kлwokJ�>�Ry��̆�~�WG�d��R�S*�X�*�ʨR)Q*�P����Gw��O�xM~#M_��Q��γ։�TfϞmfΜi�1�)T8R�O�)GH�  �2j��W���G����3*���f*k�A?hFm@zeP�V�JE:�)uH����/�U^�ɗ���\������߿ݼ`Ś�Dyh{(N5�i/�?�ޢ�/Q$D��W���h�Eoiәf�J[�l�-P��W�2p�@m'y Q �黡O^(��$�Í2�y�T�:/�����R�m۶�S���Ϗu�
%���ZX�n�Y�b��RdT�ʚ3,@7���J�V��B�iF������?�����Qua�k���8��m����]CQ#א���q�^-<kFmr��ܹsL&}����;g��Z*E#]�I�w��t�I�U�VA$�I%�N������ڣvȐ!�1)�BƍLФٽ�xʶm��rW��p���T��?(�l6����~��t*)�����3��q��\%i��������v��!������<xp�GF7���N��hFm@�Z%�ŕ�ll9=zW�p����PR���;Н�p�ߣ��OFt�ʫx����U+�;������WG�C=d�A���r���/�Ť�0���`D��NB��gz$K�~��*�-��b+�}��Q���(�N��`�ь�V����ߚ�K����(��\ټF�msU�!m�����&�]���wz���|��!��K�.1��֭[��4�-9$��� �hC���VY��T��5M�1�񩸣$xu����7�>3z�)
�+�}�3��S�:G�L ǟ��>�>�j�����/T��P������i}�Q�R4����'�۴˕�d�P�j����I��J-,~���U��;�~9��� �J�h��kE�)�AY��R�J�Jŷ����㐅�C5-�i�GmrȨ���lQ(�AB�!�k3��Rqs/��H4,�e�&��+�P-e_�Y�W-��^�zEEsJ�4i��x�9
��F%9���?�\)�9PЩS'/�Sq��ߴO���q�9�R�\�?�e�*��4iR�AZ(�ʭ��J�`�:}�t/ߣ�u�ui�Ϊsiʃ�xW��A�J��x+��N"����Ri��4�|�Q��(JYQ��(JYQ��(JYQ��(JYQ�� �讀�z���r��T �J%��˂�T����^�ʦM�r�D�CB�Ν;��;�*�y睜��$��A�2I���^�zu.�uH�E�͚5���W|���!sS�L���Y6C�1�?�iz�dƌV��Z��*)`e�=s�d �s�=g���D?��K�4T\��p���fѢEQ�����=�\��x�y�3g��o�>�$�M&L0C��
���7�Y��SE�U�Zq��C�����hȠ`�Q���9�/e�R)�U�2F,,B^!��7Ǒ�f_�˧���.Ǟ{��v:S�R�;��������K�@���#m$���{�e���|�;ш��"�dp��7[�W����f��CR2�yv�g��c�F���6o���y���MF-���ab_|�8p`$���϶4iS�R����{�g�8,���|�� +ё�L"K%�\?���&�}��_Vg��%�t��;Ɔ�㥧���Rk�pD�qd���vĈ�!�]�r�O<��y�o� ���}�BŝOC;I9a� +v=.>�X��:�J�>͈ҬFc*���/4�\r �ɫ{���~�ʕֹ��'�VJ����Ν;�v���k����6���b@��_j}*r�۶m3J��Q�EιǎU�ْK(�/�o555�V��x���=����Ʉτ�%�G)���8`��6̎M���z=�6��,�:��$$E_|M�����J�x�!��f͚E2E�2v7��'�����[��'�,n��/�sn>��X#fd�.��޽{��z��p���R�������´W,����J�"Z��k����D����_��7n\�}���K/�dǞf��)Q $^s�5��O����_�¼��k�ߒ ��=Vcī���](u�	?���e4�T'���G&��lh��!�V�D�U���ǐ�rt��9������� ��Oq�\)��Zq�^�j_U��*�Һu�G��T(�r��#�D��eРA�O�>�ZV�?E#No�������O���|*�0����ݶ�W���w�m�!�C

���y��bx����^�ߒ!�\p�9��#���w�3�/���֭[����7L1%N�&M"����c�3X\�ߒ��&-��]�]�~�zM~�0����.���NJF���6��)/xU*���)į�2+�k�|�ϡȵ�K�i��s�ϡ��R�Y����L[�'C2jݔ|�^�А���U�_"��sU�Z*4x�4�Z$IҩS�(B�{Ϟ=m��Š&{qHH�u֪U�X�r߾}m�!��$�<}�t;��'^C��^���R�E�����T	�b�@FJш\�J@�*�ĳ(j�%����޿�kHyҤIF�8t�3f��袋�����7�f��v�%�?���ԩS�����m۶�&ƅ�Ȁ�/�$Lt*�9�*��q�w!�n,@�`y*r��:��������[�S3j�|*��=��9�cwXȪO�(D�˨=����Yg���y�n�¿�ۿ�x�~�ǟɓ'[���>�[���)�?��S��Dg��[�T����K�7~<@�T(/]�4����'�(}�5�ַ��"�Q��L�X�d}��ɴU���w�i����k��:��2jS;�C�Xӣ�A�8����J��D�<`�T�ZY�&��|�đyɮOg6�{HQ�r��xG�\?X�ڴBC*��㋪8j���?�iӦ�$�Q�F�SN9%���T
G�̈��5�z�y����J�\�A��e˖y�n��Z���:$��EN��;��J�i*r%y��ۨi˖-fӦMA�?�3W��W;�׿��Q��� H��[o�e^}�Um}P(�-Zؼ@�h�={vP>��'�IހRg���J�@��L[vی�B��]H��)v� ���C�|�U���O
k��7~��k�ȭ�Y���RnA!��\�5�b	����_�G>�xu���9�q���4G"��R�4$M_�R���ȕDJ�xu���?��Q�@Ǝ�؟~�i3s�LM~+|*W^ye� �\��X�J5fᄄ��;N�EC�IV��ͨY���^�
&g~%�RE9긹+r]IF~/9jr$
1WJ��>��R�ԩSf��}��هEK�f�Ń��8g��G^J2��{�g�)r��h��C�+��<Z�li~���U���X*}��QM�9,X� �jժ(�hP�.]Tf%2{��ܻ�k�F�
:v�r�0�A4`D��1H�������H�?T�4 �bBy��q�*W�Ri h2��&T�(�RVT�(�RVT�4 �1��	U* 7�3���J����r��*�*�k׮�d����e����]�s���R�5kV��_��z̝;�f{��Y�|9E�9�Y�C�x��푲�RaBAHrKM2j۷oO�����+�TV�^���׿nP�>T�2���/�
����3p}O�KԚ}���6Æ��������mW�P�U����y�o�؍i��N�8����;�_�}��Z�A~"W��Cd��t�dc�c_j���1������m��&{Ղ�`�K���`�'Ɣ�R8b�;������ZA�R�0i�${Ėk>�ڤ��;�j���^�'�x�}*Q�g�}֬\���ͨR)�J5�#L���#�>��V�b�� ������ϛ7/6�I�{ںu�����o���m��$_U�~�bǟիW�5BH�SjǞ�a@�4�V�R{��o����0[���X*Y� r�wBOZ��?��Szئ��ŋ�;vx�n��
]�e��*��6�8ee��@3�J��H-��8�r��TJ�J�"�
�B�ϧ��u"g���;�SI�X*4eb�q�F�b�
�t28j!�
����Ja��Űf��������O����oI�GQ�M?�	������US��P+WN��*��C��2��\��j��m׮�}X��S�~�����.������X)�d���L��!$��2ݺu��u�uB�u�]g��d�P��Y��TF�iN=�T��Mr�%��e��3�><��RHy�=���z�n��o<�@d��R�)��e��{"�BC����J���M�=�cЌ3�Fd-@�{^�n���������$�����l޼�:k5�-r��2^@����Y���j��*rT�8�$?�N�
������� W��;2ł�d�a��.L��S��;lM�}Ll��;Ǐo�����M��9��
�K/���܈[Z�ÿ�˿����{�n�>�iӦE�\U�������0 R",�?�O�Q�C�a�c��Z���g���o���y��!����O�������W_�����B�ڵ���\�,Yb�બ+���7�>�����/� ��q�*�o������ZT�T�JE4�G"���UU^ɑa��\y�&WBʩN�'KT;�ׁ\H~�Ձ< ������>�/�m�G�� �Q5����C�+�Tv����;�����C���Z�^����BdGͨR)��+�(�s�9��3������ޚN�"7x�E%�)9)����}��Ǭ$ͨ-�?W\q�:th$ן��綥ħ:T��xϨ������\㥋?9���?���ڐ�J�<���o}+j':�@�I�O�V)4ȶ� M_à�!G�&>�v�gؖ��N2�>��Sދ
�Z*r�U�R���w���[F�J�������M��1�,������OG}�ZȦeW�tr�&��7��&M%@��j���
��=�4�����U�lٲ�(q����,{��5555�]I�Z7$�;�脦i��ūOE�	�:p��'��'��+9��o�&S��T;jG�mT=��"=>:u���S�����6����A��3�>����p�ݟ�z�����xuԶi��F|kΆ
r�"��W�l�9����0��H�7���mڴilp{��%�ž��Sy���u���45j��СC�WY�h�����E�J�H�_�s����5��gm��%|s��j��0&��|��8d]��޽�l۶M3jK e�=۵k��Ԧ���J�{��ZP���կ~՚��֭[�N8�>���G
5� �V1	�4��$ _��|G��~����Б$-y�űc��>�2�0���`$��I~��gYK�\�7�~�#�ㆽ�d��AA��k��� �����B�����O~b}U�T����.U�H��,�L�9+šz��i�����E���5^�y*�6iB^\��*��H(�m��q�6
���/fť۩S�̔)Srxݳ��2�Y+��8�;�<;OY}O�A�����ҳن��?z�T/*����2�zp)S��q�F+~|�u�@4���a��رc���b���+�uȆպuk/7�e�6m�4�_�-Z� �DȎ=�X�Y�̞=;���k�V�T�F�����#dGb�q媎o�Ri ȹ?�oE�"�JEQ���JEQ���JEQ���JEQ���J���|��*��;ۇLPm�T�n�T�TU*U���&�iӦH��"�v�Ν�&M��ɒ��۷�V�\)h�Jw}��T\�l޼9���جX��(�ajc߾}����mr��w�u�Y�j�2d�&�$������ܳgO��°�ez��믿��Uŕ
��ҥK͜9sl���Н���Ҩ��: ���0��P�ٻw�h�!Wj�,XT�3�$>餓�|�����ۿ�[�X4c�.s��ެY�ؿQ�yꩧF)檈G䊒n۶�}%2n�83|���גIy�7�0e��|�����S�i���0��??<���۵V%!�/���h��~�t��T>����5xu�>��F�C�z|�,e^�z��Wm�f%+���J{����K/�~�!�=���U�0�%���E�t~W<,�]�2z�)�(JW=��5eDGre܋益W�2d�{z iq����r�W׮]�����aQ>�u$��U��=z��2�1�r�g̘a�m�ěR��֭[�U�R74�Iz.Xt<�jެ|>���2q减�^֟��[o�����)~���4J�9��qGt<��Sf�̙�S)�#:�M�fSB�PX*�T2�8,��0I'W���+G��?��T��Z֛��=�`8�`�+�#r��E�(��� V��d��+�G=���#G��Tj{����$?<ra��謟Q%\4�=��cc�h�*�sI+����_6Ԗ�ī�����3�Th!
��� Q�\#�,Q
�p��a2�D60�kP�iF���^����Ӎ>$��B�"A���oo����?~T��Qk�`D1�iݺ�}����Z�pa���\��A�U�����$�(����{�=Z"شr%$|}���k$��C*�F��W�r��WGY��S��&:��찼�fz��y*	�B��;.vmԨQf��&�<��׿��m����o�i�����,~��k�X��*�d�\��	3Y�i� 箥T�T���O~b�8RPx�FIZ�>��&����������O��<��R����HR�$��IZ��&�I��P�G�JD�U�w"�l���(��:e��u�)�!�*n;͏�׌Zι�[ԁ\襊Y.r"܉��<���ˍ��#兓���+�t�>$�џ�S��Uw�Z�9��i�'�*�����\{�V���8�"�ā\�+���믷�%�Jo�n��:�}���ĉ�t����2J��ώ| �'O�]�ɨͨ�R4�Q;~�xӿ��~�}��%K�X�\�n���;��>�]��E�q�Ʊ�1�ڳg��U~��R8(����]�vY��R��ɫ��j\,=�����J�CW&4k�ܹ�}(�z�)
9�P��υ��(l�Fi��l��ׯ7{�����^��g�a3ECW*r�R�ܾ}��:/�/�;�:kǕ+��-[����M�6��V�,W�7�R�T���Oq���R��4(�G�t��1���իW[GcFJQ�b&��01i~�9��Y�&���ϩFV�ׂ�^x�(qH��L����.[�L���2=���mK	�![�x�M�i�O5�T���2���)��*��r�"$�V�ˢW���,��E~h��x�?>#;ڴic�3z�)q���`xar$
�M'�c|���Q{�gF��կR��ԩS$��ݻw��F�I&�a���S@�}��"mi����|��'�ڵk�~�WK�p�N(���O4L�)D.|�cO>EV�JQ�
�w"reǦ��8j3)���FN�W���c�%�oгg�h!����6�Z�ߒ��K�#���Ν;�h?���U�䏡Tje"��)|S+%9�O
5�-(ħ
�z��_��>��:`�sr�	����.3&L�PBD����������}g6���I�&�0�O��v�m�,��Ŋ�%G���O��t�k��zԺ+�+i��G����Y�˗/��a�.WdA��o�>��\Q��$�#
�ſy�f����o���2x���,�6�5�O��	��R��(��w�w���̒s0�XfT��/ˬ�J�$f����(�t

�H3!��Y�Z����i޼y48g%G!��B����d��T\��l�23o޼�Ν;S�P,nIp�'I�β�U^�#r�C�
2D�cƌ�ZLfS*�?�ux9����?�_0K�.���=�J�Tf%2w���ƍ��<X��i�F�Za4� �4wC�!�QT9Rb���'���U*��Q��S��r��*��.~勌*EQʊ*EQʊ*EQʊ*�HFsS�/0�T n��&��|9�\��J� ���R:��h������2mڴ3W��~�ҥѐ5
�f͚��ߜԭ(�!E�L�}��ؓ{�7W�Q��q7&)�ݻ7-6*�cU\�lذ!w�uי����~`��Ǧ��i��fF�5lf>�hOreH����k�!�'�x�h'�6�J͓di_~��^���J�pݺu�EM��R�CvTyɘS1�ݶJ���?�vϗ�i���=d�/��ݻ�|����r�2d�v�?�������/%�2H<���`�ԗYʢT��B��0�Z��駟��Jj�������y�*�Z�KiݺutY1����&3�� W��H;N@���A�!�S+-_>�T8�*q�9Q,��e!�z��tDG	�N���2�^F�舎��5�L?֬v��q��GG��npȊ�eJ2h(���y+ǟP`x���^����x�����7?8g^�T�˵�^k�*��A�X#<P�U" 7�x��Uq4ʤܟº�G���_���ގ?<,�^zi�Pj�R6l�m)f����#!e%X*\p�9餓�����S
Bh�%�>$�x�������Ì_7��C�dA�J2�`���C��v�!V�ǁ��4�*#։k�g2�)�r�jx��|*�CR�8����Gw���Q�֚��54?V��r�J�k��E:BE�ӰU�V��פ����#�Q��u�q���:r�H&;Q	.>��{̬Z���w{�.^xU*u��`�@�gT���5��m&Ҋ�I��џ��5J�c�9Ɯ{$��ӧ�ٳgk�[	U�0a�i֬���\IY'�ӀF�T#'ǫ��[�n��� ����#_ m��|�A�z9���bqw�6m��5��!�
W�QD��o�s�u>j�[�)����B�	}/Z�h��R8���c����ҡC{-�JE6��S��S��n��-�>�h�������B��,4Z"Wh'H�f��|�r{�I�(�Gn�o�&��yK�â�s�)�D;�+̜9s��u�xH~#��k׮��t��W��o�E�ߪL~_Z�?�Q�$ܤB9~�\��J���2�\����7�Q[�i��k��+9�s�VP2��B���?�V��T�����~��D�:u�%���ի�m}��?�'���"A!Bv3j���g��[&��v�Lfx��w�~����x�}k����%�^�l�iӦQ>EF���Ō���)�Ƌ�֠X-!�Ud��Jϻ�]�"B��:Y�W�6�-���\���T��5/��o��v!e!�!�w�y�(q0���F0W)�4��`���ͅ5��CJӯƽz�T�;�<��8H7�Ν;��}����+�T2j�2�엌Z�FF�T��]�J'7l���^��k�>s�h�~-"������i׮�ѣO2$�A�k��v�	'�����I'A�{�T*�5��o��(q�HƎk.��(�zFthFmrȨ�8q�:th$ׇz�f*눎��է��ٰsJ�G>��JǕ�f��C3jE)+^����;ER�y����y�uPy���ͪu{��TPȤ� ��Zδ��ꨭs���#y����m.���|W�R8�\��$�]y啶Orڏ�ro���7�l��|��Q{�M7i�쨴=1bD�@�M�f������D�h�I�+��#�<b�B{�n�:���է�r�J}H��7�ʑ���$�c���[�l�	��GVT�jD���T�?�����Б$-Q*"�Q�#��Jq`��ΤM��EHB\(�o�e2�}��R���!R�RWP���W��\�|G�hAaq��$�u�8jY�2^6�_EZk���7�2,���XjwT"b(ZR����1��R�JB��/V	���[�l�Y�pa��ߎ;��W����!��JR7Ik�֭�I�f�&����.���8���6�+�Pr1��P}���O�.����cmМ���j�\3Z�d�JSq�B_�SO=՚��8�5t�En���;s�y ѡ$���G��ȕ�o�a�ʚ(={|P�E��mEr�m���N���ꫯ��r+��n�)�a��7r����;Z+�������� `�֑���GF)vg�T���z��*� �=����YI��A�T�~P�� �p��EF���(eE���(eE���(eE���(eE�J�mĤM��G�U�~P�� p+f��R:���j��7�(�U�V�(���>��޽;�M۶mf���9�Wr�+��R�C�A&?.X� �x��v���Y�f^2�+�T�oߞ���l{D�G�\w���6j�> �>��ٸq�N(L����״m�6R*�?���T�Y\������>���U\�`�<��v��4#Rꠝ$ʄ"BY�����}i;��Ч��2�e=k�,3o޼`�Ir�R-Z���^ZHu2U�<4�1Zס�o�.4lz���m�&��ȕ�y͛7��!;65A� :��1�@��/>�/���c�R��ŏ\h��B�Z�C�M��R�Cp$zԲ�!�P�z���S� ?��j�8t(9r�7n\��p��L��Or8�����G���c�� �>\��T�{�א��\UK��L���Y�R�A�&�R�/ Ӑ�J5�Gޔ
��n���tBa-��3ݕ�9�cd?g��S4ݡ�5�\Əo��e��=?���6����Lz��:�C��O��e1N^�b��Y��-
�+�
�#9^��i}�W��b��g���K�G
_���bmܸ�}���/�\���+�D�aU*�#rŧҽ{wөS'��.^�؆�C���S;�P�6���GϟC�5^��09�4���R9�*�t(q8�;��L>��+9�܀��LC:~˔�T\����Ç��~��5�o�L�$-
,��}�F�H~s�)�p�	V�!���F��Z2�x��\x�6�T�J-���"���7�V�V*��q��ș���O>9�ӌ(�]�V�p�W\q�Q��3f���7�e�>��C��^3���3J2���ކɕ�ҹs���R��T���>T��t�3��.�� W,@ٱyg�!�jDD���;ΫR!�H�Tj��EN�S�>��X����y*��)[�j]�E��o�u6FA!�8�īOG��*��ŏ�%OŅD8��ͪR)
�+2#WťM�6ւ����{#�6uJE~<~�����1�v^2��B"@��"�U(E�\�:�([P����PZAa*3j]|k�/$b�;E>JmMM�ٻw�Q�A᠛9�\�'�M¬,���ʈ2q-�NJǕ��U�~�T��S�C-��	U�C��M����U�P�.�͕���oD$܌Z����Ѩ�k� C|*n�����6��B�?���}�5M��3ΰ9�O���F�o�>R&M����U��L%�O��ٳ�U�UK+�q���3�ׯ���ޓ�xXT��)[�)�8���p�C��F�*�����Gr6��~*պO�J����7JL�s�=�t��%Z�3f̰}?4M?9��'L�%�![��0�$��r56p�J��Q���?>�Kv��Q{Ԗ ~���U�
Y��}V҈X*Le��9yͨ�����O�.�󿴃��K������O�r��8�/��R�7[6 �
�z��[��'^�����:����N�g�رv$�(FIP�LFm6N��\�P�O���|����?J*�<y��R%��=3��7^{��ܹ�(q�M~F-�i�{ｪ�lIb��ʃwdJ�zH�$S�S	�,[,� ��b�+�8�Ä<�T/JE~`LR%	ZR�,
FBʡ���=jK���!�������Oŭ���[�,��q-��nF-���=��R�\������_���mm:E�����M����E�i�r@���6m)�M�6�-[��ݡr%�ӫW/��2K��AQ�R����>�)S��F2*u=j��ȇ���-�߈��k��~F�3g��G��0��?�T�;�(D�J����ťE��z���R��]~�7�kY�i�U�kf����M~�!C�DM�5�vA���s����P�T��-(Yk�A���`Ѷ����y=��3�V*��n�#t\��B����L���|����J�d�ߟ�Z��^���?l�8D(Ȩ�)�$�͞=۞�5�-9�Tx�?E�J�&�iDG5�T����E-��s���L�>*_k�K�>�F���J-8jɛ��
��86d\)	%�H
7%'(D��U����:djjjr!�[r�y��_���m�JH���#y)ԉ\��N{����D�~���U���l�͛7��,�ŋ��{��,��;��JdΜ999z�TP��ڵS�V�� ���4�S�H)�ET�~P�� pC�Z�\>�����*��.v%M�RQ���RQ���Ri ��Q�haYP9VU*���WZDX���ޔ�Ν;�7Rw�:p�~��Gv6�$d��m۶�&�%�^�:R$ȗ֊;v�ȅ�\$ФI/�����&��_�2��V�Er(�t�yH|��E�*I�Q� �K�L�+�
!ɕ���}ƌ�aÆU��+�T֮]�c��o�a��Pu�9瘋.�(��y�G�ba����_����YB�<`�a�y@�����|�K�M���Qr`'e<��SAN\c�g�R)��4��>�B@�b��w0=�|�z�T���.k�k��Z$�<��\`Ǟ�s�xdmI�(^��i.����U�7���;�0o��ft�ޔ
7x�=�h9��[j,���N;-ZӧO7˗/��_
�\�TF�ez�������2+W����I;k֬���^�pFt(q�t�С^��%K�h7���3p����gÆv����K5�իR=z�m�G�Z8���v���~�����F.8g�J)i(޶m����N:�6�!�&�GċM�'^�
�(t�X-R��������V�AJ�\�kͽ�L���w6�*9�U#��K;Iњ���Q�c-�<�"�Z�ܹs$+��8�>��M�/Q*(f,f��cvٲef���	�Zٱc����j��Z��(q��k׮Xp���fݺu�M�#?קB�N�l��ie�T�J�2��1���ǥq(�q=$�V#}��JŽ�nݺ}P�����_A/U�sR��$?��ő�e˖v�cH#c�x��x�Y*쾷�v[�C��,t���ŵ���ۗX+���ȐP*9Q���ķ�[�r�F��r�-���7�:q�Ī�blH�
+�	���e1P|�ꫯ�< U*��ʕ��+����"Wj�̙c�
Ӯ��9�w�^���էR�l��J�A����x�����*��p劕�C�uԲ�xI-Lr�F�W�ұcG�=sz��vT|*�︾�-Z�p(�%�ǟ��RL�l�/�ˬ�B�r�6m��էr�e�ٜU*u���cֽ~��'ہ풤�Q�R02:���\:t��۷ot4Ȥ\� G��K�z�n�>����w6�O�J-ȁ$�����f͚E��)+V��џ�*����#G���Y�:o�<�XBK	9�������g�6J��Z�nM'DV$������*�'�xb���/ɗ8j5���xk}��|S<�>|��U�I�67Q��xQ*�C�"W�Ed���˝�,��?��Z�\��"Wd�Y m:�G"]���^��O=��(�1d��%�OEZK�NؓprIZ�ĕ+�?D�܄8R�%�6H��?�>�R�����(�P�����]"b�:�Sl�2Y�U*E�LE��ș����|+��+���?�iz�
7H���ķ1cƘ�/�8�N>k�,m'YDH�'7E��w�}�����N�xu�����T'0�wB�2��E�2+W�����kP�Jr%��wU���ύ7�e��4.ʨ���",���VqĒQ+պ�}r�g��&�cD�/~����o{�~���\�A�H�k��P,�s�]�ּ��;��V)��+�?����8v�l J���ݻ��׌Z��� gR�ݚ��=-�z�2�:u���-��{�{b�o�c]5֐W�ʞ={��H��h�@�.M�/7����4M��xU*8 3�t����b���g�w�W2D���P��5��dh��߾��o��䀏	]~x��Qi׮��RdT�2$���G7�gРAv
�]��fx�gl��O�F(�'��J�Y�n��`�b���B���e!�f�#�]��4�1��k�����A$���Z�)�b���/�ͭQ�C�~��ߵNp@��?�����J#��O�,ev�>$1ɑI���g�KҒʬp\���MF�J�ar��xU*��<�Z�^��մ
�ɖ��OѠ�9��m:�K�.v��X)uc,0�.(��w<��(��6h�޽{GŬV)�[�)-:��$C�K�}J��^�m�fR]Px���%�$��s�F>�G}Ԟ�u�rrH*d����_ e���'��Tc���T�L�S�l=���m'�N,T�!r=Կ������Tk�S�#��n�&vU��T�$�c6��!��Z�ځ�*�T:v�y�r;v�P��A����y�ַ�e_٬:i��f&���\���*��DBAf!ᨾ�;*�}^,��#G�&9;w�̭_�ެY��*~|�'�p�ʬv�ڕ[�l�uT��B�q���r�0�)�.*F�&M2�-�ɱG¡Ji4n�83{��X**W舎��S@LU�tD������~(H������CVI�Y*���NV�����?9ɥ�]UQ�ϡQn�̜u����O�ʭ[���#��(���FfȐ��/Z�4���Mn��(�r8��sN���+F~B�&V���#������d�4�\I���ٴW��D�*�T�~hdn���/�����,?=e�IS��vӦM9:ć�]�L����d����+r�j5�i�7n�)��[�2O)�(�MR,3�>2t�kѢE�͵F�+́o>��+����d�m3��?H��7(��n��NIS�>����Ϝ~��Qo���߬\�RGI� �Ç�%�I�����!B��}�(Ӧ�a��K��	-v��������9�cL�����R�"M����Հ���n޼�nn!e,ӏW�i>8��k����H��~	�?�~��h��b�r|���ѣ�СCu�rB���e˖����R>묳��H;��~8���������sh2�I��#�_=�9�k_3Gu���&Jٗs�-[t��qݐ;S�h��.J� W�&tw�0-8B&&J_�{����Θ9�w�բE3r�3lذ���?��?��cƌ��.D毾���;�o�>�$�2a��T��/�hgTWclE��J;�w�}�s��O���ms��(� K����
4ln۶�������� gH�K����i�#�d|iot�0�tk+Ǐ0d�{����n�ȃ�]���,���T�F�h(���G�V��૒g����Tz���k����1�XGb91�j������6+�G����$�|�OM�2������ب������;��p�ɓ'%#:�;�<;�Fd5{�l3s�L�Q)�m�6m"%3c�+ېFtT,�ê��K��H(��=b��R��ֵ�
�W�t��sj�G�#Wg 2�׵Y�X�*�� Wp������E�����WX;I��j��ǩ���Z�� NY:����3ΰNEI��ݵ0d]��pxK�/��!ȕ��:u�-�����6l��^�T�
;'�^�u���g��*�����3����v��e�*��,W��j�zV�Y&%��+�DٵJ��C�|
,q(J���)Ł\��q�g����.]j�|�M��3X)���5�{��5��đ�ʄȏ���4�r����p�����^��5�\s���8[�js(���}�G���GZt��)vmԨQf������pϏ=��Y�j�����T�I�素�7"ᆐ�>Q*U,#rE��Q��B�⠮F���J�}X~�ӟ%�$���/>�g�}V��J_ՕW^iN;�H����o͜9s4���x�T2��Iv�h�_�䷒q�%�0��TG�JD�U�+�U�~�Tԇrh���R�����x?T\���κ[�!�T0�EN�;q&r]�A�#k�IN��p=�~*4���@�k���G�II���ΉӐ<7M����2�^{�U.�(�HP� _Q��_�U,!ȕ�C7�p�u��ěRᇝ8q���?u R�ir}��gG> �/\�P;�%D2jǏok}�~�}��%K��������v�֕!"ٳ�4�FVڣ69(k�>��ZR֑kH!��g��NR�������,�:���ݺu���Y=�r%y���.�WI;�L �o��z�-;��'^����eԪR�[�$�	ȅy5�P�R<��@��e����w�{ԺYش=H�Rqo��>�Zd�s��Z�NEd�~�z; J��LF�*�"rE�(��!#O� ɧ�g�����Ra�+E��t�ڵf޼y��_���=����:���xU*j���m�> +�S
�`�MC��g%tmL�w���i���'S
]G-&;���(�!�Ď<�Ș\�V�<�~*��(M#�x˨�&Ǎ��ġx���߾}�kYu���L8V�$��K�np!����~��_�O���/���Z*���n:x�`ۨI������ŋ���J�xP*l^�VJCx!S�Dոgߑ�z��I���Q�?cz���f����-���>#_"?o���~*�ūR���hxԅݔ�B�eUV�a��Y)(�z5�L�����kA�>��0��bB����̄	��MJq�\ݮ�\�G22�Y�N�4�v��W��m��VoWQ�(Y�4�����O>i���Q��pD�$��=����+*(�6m��WI_���Y����O8��J|*�M,�͛7[���T��O��Vyg�k0T�������Ը(����`����2K������\��	���u䫸R�1b��Ȫ��A"w �ډ'�h�>�(Ebpʒ�#�*�{�)��H[hm%ŧԧO/�Wq�Ҽy��ʕ+s$�}~m���o�����g��X��+2�_���3f�ʹ���*J�Y�f^�ϋO�K�.���	X�dInǎV����v��QeV"s���I6)ʚ�5�e�r�0�i ���>���(*�)eZ����T n�*m`U>��r��*EQʊ*EQʊ*EQʊ*EQ�Jٔ��[1J�s&2���T�2���*��''�O�R:1Yft*��@:�Q�JE*k�Xܵk�ٴi1QU0�χ��ݲ%���P�g�Y�vm�n7J� �O>��N%p5w�_�֯����F��G����e���j�,�
�'���y�&S�m�Q
��	;��@]���Ǝ>՝�4(�����+,�J����Cj����!{�R}M0*����_�n]Ԭ(��E��5�E�:��ถr���Q��V�#�1<�c�X�����s)�e\�����	q{��A)*W?�T����/*j���Bz"�T�8��#��6����)�+Gy���0�r����CE	��1��p�Thl�`��sYC�C�(Jz&}�Ѷ����ۂ�}���,]�$GB�4�Q%�p�YxӦM̀��r��ѳg���&����f,*��R�h�0�q���͊)b�(�.��@Q���JEQ���JEQ���JEQ���JEQ���JEQ���JEQ���JEQ���JEQ�����Q��Nr�    IEND�B`�PK
     uK\;b�i�  �  /   images/68998569-73de-4f26-b1b3-0b6c45f8499f.png�PNG

   IHDR   d   �   �Sh�   	pHYs  �  ��+  YIDATx��]	pUe��ｬ/�d'	���iDD���D�5%.���"�0�4�RX��V=Z*��ڎ��*�"(���=	KV�o���.�0O*y�"��35ͩJ��q����}���8`�����FUU���z�k !!!FBb�q���W�^F��L�$H^n�a8F�����w��t&�4�@hAAA�!���~nhl4o��tyG�q������f57_�����1JKK���[o$.�����;f���e555�8�� ���K�?.�xu�������wٷworKK�� ���������r��]�����D�?��Q�S�1n���o�$qc_��a�硾�[���=� ����?^w�uFzFƔÇ툊�
5�����ƞ.,�^���2���9s�a��D�+*���vWwNK������ĸn��Zz�����g�wX&/5���I���.�ҥKŶmیjkR�i<���gΜi��hX�bEq���I�.#�r���%k׮��i��L�:ՠS�8��h�w�>FAA~�jK4�M��j����>F�%�^X�����=���ZD����:����%�:&���W_��ETVV�?�Y�]�*��x�Π���Ν;�s0'���l��m� <<��6��u�ֽˋlH�淚��8���8����Z�OA������e˖W�.�p�ٴ&#�����_������|@�ैΊ�
�gI����B�K��j7��J� I �e-��w[� >�������亿��&pc}����J�ĳ�6��3-	�����5�2�t�U�	"��a\�p�8t萹 � p#dt��a��A<�cǎjGVЀ�W1$ �Fl�vVV�6� �����nR*	�'Nuuu���XTŃH�R!���8LN�:���J7��
��}q*%��1��/��"K@p��	&eeeƎ;]VpC\2�;w*���Io��-	��f��&��Ax|A<"�S����9ڳgO�VVII�Ix%"g�N���p*���M��T�ς�hii��y[��f��gQ�u:���U��W�,K����l;~���7n�q��y���� 7�^���g��nCZZ���m2D�C�!D�d�����^����j�u��1uf/ �T�:a\:uօ������f�]�͒ ��.l�g���?��_���R��l��pCd�J�@L�;:u�Bϵ"�a:-���_gdd�$�E� t�<d�G'%%}@VN�֭[g>��455y����ߣ�:2����i��x�/��HOOo@,�����;Ll��СC��F��J@�~��իW�mܸ��d�����-4�Eh��O>�Ĺ~���j�o߾i���ƹs�ငb�\�̖��t�R1b �´�.����7��X�*�/���˕��XG"���@`Ix���rKOæ���DT�l�Ű�����:JOP`�&�L�Ci���}p#x�px;�&���'e{Ǽy�!�x$e:��СC����z��wst�A��ɓ'��~��9�G����?ܛ�ee Ί "D,�}Ni�"Iaa�Sw���-((p�6{�TӺ�F�if$I/��yK1D�a;]����o��u ���H]�^%�bt^;�z����\q?��vl?�q��CP# �1���(`gd�t���V���C�C%�<��i����d�	������o�-v��NH��~a<P*��b�+4��:�����V�ԑqU��F�l�TꈶN�6�<M?���֪{�J���j���G�jR��}K�1B\��(III��Z�\n��HLLT����e=�6�$C'��g�4{��A
���y[�,83�f/W~�w�}f@q���Z�:�ܐ��qs�8_i�	"��~6��g������7�N�N�9�S�N�V�N�㩛D�u��0��l��	S�V]��v�^o�4�0W����~�^'s6��A@��f.z��{�>M��jء���	BP/��cy�%:9�ֈe���EY�wff�+--����=Of} H����{�����䑅i�iӦ_�v�?{���|�ג���6 �ճf��2.�.T��a�-,(�!KބB����$�^��^�zU�� w?v�ؚ���I�������ܻw��C D!�b7�8�$�A��@�#;��ڵk�/]@����>��0`����|͚��JP5�x�������<�C �C%�Æ����1q��=:����l�ȑ#c;�X��I�&yU�&�w%&&��'?v�ᨶ�� ���<x+��f/�M�����nt*u�F|�&���:tr����V�AB4�7���f�=�tT.bc$C����(|�����اg6�J��!�C����C' ^^g>�qb�p�9�"��ǫɇ�E�Yݺu�|!�\�=uƝ���<ڋ��OY�q��;�8|���1�n��	�;`��
mҡ�g��\�6�V\�"W�A��Dӧ$`3Əo������� ܥ���7�|#�Ci�܁d�!dxrr�1f��:�Q��z�x�ѣGM�ZIƐuN��������Pn�U'�!vE�m�H�!��)0��K��j��L$k%a������kvӝ�p�RǡP�N<�����h���Y �n��G��z4���A�v8�|;t�J��\��ܶ�!���:U��t��Ч"cx��o4Ξ=+vj�S�������{ll��u�p���@"��*�n�1!sp�믿>�~��)�¥h!��k׮����E�f͚�k%�
R
�+|ǎ�3g>B?�(ƍ|�i��ȊV2ȁ��S�Nm�.�����,[���{�-H����q���;	w����޴h�"允�ӹsg�A͖JZ�x�9�@J��୷��[���_~ٜ��+�?��s� �>��#�_���5�}�Y��Z��TTVbsr�<RJ}���M)))}H�F���%�y睃ׯ__F�]��:|�p�����v�m1UUU����6�E���n��A_MD�cHG�awxx}}]��KJJ>�֭�G��d�w��ݮN�:!s�TXX���#�	�*���N�Cי��@=�W
�*(�ڿ�92�3�}��%�>���������f/X�F�&���^��􈲲2�ĘXZ���[;�,�󥃋<�R2�n����;�a���Q0,�!�d����srrڥ��8����,�{�����C�w���y�<[Re�yz;u� [�E���?��=GJxˁp��bܪE���%��RB&Mr�5����6��[�N+A .�����'[�P�g�жD�i�͊G{y�4p�·��D��j+�L٘Xv����f/�q��sF��2��#�v��'�P���R���@���3�j�pF�ؚu��>���cb�v�
tV.�ո��>���P��-]�Ȧ'��q;p�U�W�l\����ey����q��V�Yd�_��J&6R��^���5��3�!w�鶲��� �SSS�i��nL,=(�N���S��Yy1/��B�'������i���U����>�&��			�3g���~�t��d�����ԩSC�E��rLlhHHy~~�,�Z)(�?��!7n��8�`�ʕ��~�}~�2�˖-�3:�D�	&̘;w��R����b�2�Nb_�觤��Y=pKKK�}Γ�믿6�{�93K)h}�3gN��={d�:�o�s�NFl��&�a+��O�࣏>jHN����ʣ��2��o�]ך��-��-{KJK{<��c������Cajg$���'O�����fgg�F�{�̙o����߫�Q�S��ŕ̘1c��'��铜��999�pDT��������m��0~ո�,��IVL�2%��,��j�$h�Љ4AXl�m�+���X5A|)�M������͐:�>��D��vpb�`ܪB'��[!Ϣ��/�F]-m����8��:�ȕ�J<u���]�Ll����x&��;�,e�^nG��}�?�^�E{�27Us;�]�bkL,^RǘX�8�-�� t9p��,	������Jw�u�x�D�ŎÇ�Zu\��T]u�\r=J�>�� fi	�g_�GAx���fE�
�d=��^p	�,:�^�Py�sp���y�V�1Tn������^�ҝ�ǭZ��Xef/^�9:2��������שz����
���^��yY���1��ƌ�6{9NF�	2����	�ˬ��TEDD�%��^P�x	��m!�a�_qA�#j�Ґ)<}�4p+��"c���Q�ڬ�0�_I�����l}饗ҡ�������e���qy���^xᅛ1SUS �-��a��ݺu�"�\�駟6��I_�7�6^��^ �\+�z�և�Ț0a"�rss��I�oD?��>�رc��W �@��=zԫr*#�#<�����%�p*��8�Wyn&�	�����2�DE��4�!$��đS�/q�Ҍ%�c�Wu�'�`KpHHd||�L�0T�H�){>��c7�"a�$<x�ϙ�1=�����B�$c"d�ҥ/b��J�E��Ŵ�$����	B���СCw�Z��%i+��@K@��͛�Mwpc4ӦM��Uu]�9�կ��ʟ.TU�GEF��y+�tCەVq_	\~b�����	��ĩ��!��.��"�e+����o���:��nv:��N�!�s��I�Op
�HLjo���{��J4}"�� xQ?��MM��F��O���B��Uǲp���J:��>��-�r���P��X9fܪ�!�Q�!8�|K�d�g9k��a�1i�$�����~R�U;��� �.OS:�Ε<sQg>D
7����
l'ㅤ�Ϙ/�j�� ��*n�At@u��,���.b����KI�4U�N��b\V`��ә�uȸq��t'.֭C$q�m �)�:�us��;��@\!��v �����j�x�\`)3{�Gt���C�s{�o�Q�N.�����Sw"�#�s�'Lϼ��v���U{������p;YH˦Oz��ӧO���)ְ��O29ͦϧ�~�#CO���M������Ϧy�������tL,���.]�4\�,�>I��۷o6)K�,�/���fӧ��.X�dɓh��C%�Y�V�B��4}���O�49U@"�����7}����")q�i�B�2e�y�����.�q�ښ8q��W����Qh��(qG_��������>�6%��z���×I9���޽{wHqqq�[�`�r� ��h��<������y��[f����e���!=�񤒒��͛7?��S�<y��1��/�čgA��(�|��?����������6�&�/,.�!k�bk��l��X����fC�"Rp���/�;��[���=�������!������`TH�V:&/�b9ՙ4`o��!����! �n<��Ҍ�t����$��pgU�Ƴ؄V^� �e����>up�}%5�OY����TR���mѺv8��%�����3���+N�קO�;|[4p�.rPZu�o���˫�d�*� 	�WJX�C�#H��� !�}��i7{7���!\(�$cȣ�%M���t���V=j�B��]�Ӗ���>#J.VkO���PN�YW����S�,B��S��Z�7p�T�X���O�V����+'&&��:cH'5�^t�=���riii�Ԉ?\^����A/=)**�x������8E�5w��1-!!a*�qcǎ}��V�4cH8*����-��zW�0��~k@]9��� �˺HUҩ�\� %׻v�j̟??bӦM#bbb�l۶���pH��vѢEA6l�'66��ʕ+�N�6�T�E!b�փ�����C}�����Y �d��&(� ��.�����֬Y�E�c�����<&�����b-H����\����SX�Ѡ������� c(���L��#B_�%��t��{hu�N�*�>D�$��c�!O?�=��;��}H�]Jg��4��^�x�_ϟ?:�3g�%ueeeE�={��g�}���{
������}*���%�H�L�4i$1bU +.hNEş��q11QY��=]$���u�d!�޺uk?��ҁ� 9r���.p���Ѽ��ު�^��XN<x���@7��^���'/�>�:t��_`F��o��\���	\�;���R�N��7�����YO̘���b�~}��J���lt�`&]���p������U���!P���K�,���<`�1��{�,))���(,-4����n�=�3�X�j���n+t�d��ڵ����Іd�	���g]�Qf)�W9��R?��������u��޺u�D$.'��q�$���"��<x�Q�F��0nٲ��	��ƥ5_~��e7}"|o�=Z<c���cƌ����f/�J���	��XdA���������%�	+�n��:��k|��n��*���6{�q���������SIq��t>�'��u�C7֩z*)�se	*�,�$����<ZC�{��r�(Ə[��P�E�V�l���!��n���:�й�ԊSbninv�]^��iQu"]t��w]��[���G=--->NyYY��N�64�UWUm]�p�m�`�d%��=x]^^�w����ԩS�	'ʗ�b܄�#�]���f������ Ni$���@\bś���Td�vK��1@T2$<77��^��w�ى���
Dʰa�\���~��۷�v����
��m0V��w�$X644����Ԉp�I���K��޵�M֎��E_,�D��3��s�<��[�~���&�[%6�,:wn���p�[�m&rx9x0M�^�'u����Z<-)C�>��r�ĉh�Ȱ��O_�ܾ!�B���j�>=���� �O�%�{�LH�>�s�/'�@x�14�&����͝+���`����$�y�
��XC�����xR�@�PȚ��Mk�ԕ�����Q���f^� �$׺w��������Ki,2��_(""bݠA�N��N�I���G�0v�������^x���@z��Ȥ'}Ҝ�����ǎ58|�	� ]�t1H��b�߷o}S�5Z�qLk̐��BDp���ۯ�q��&�\���` 
]�    IEND�B`�PK
     uK\1y1�? �? /   images/a003a845-706b-4c0a-bac4-0f60a60b44e4.png�PNG

   IHDR  �  �   ��ߊ   sRGB ���    IDATx^�	�egU.:W���ש�T��*U��-�!(Ābs����UA�wqؽ瓇��W�\E쮠�D�退H�`0�44iL��RIu�ow���7�?�Z����8���������^�[�?��O���"`�X,�炿{��E�"`��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%t�,��E�"�	���	n����E�"`�XB�k�"`�X,� K��&�K�X,��%��<ϝ#G�x�N���81[{챣���%��j��j��,s��>��J���+"ǩ�T%�9n^���={�d����##��z���������8�]z��E�"���L�#G�c_�zդ�z������ԡf�##����ONf47���g��%��{�ǯT��\:==s�c'�����t:a�R��8r;ݞ�q�!y�GI�wף�d��d���F-�d��k[�nyzrr��##�����v�h�a�X,_���;]�馠5�,��Ǳ[w+�U*��[�~�N'Yd���D�٘��ٴO������%�K	��wܱem-}�����Z����ʔ�u���$��<''Igqq��$��rr�����|xd$+A��I�eY�l4{�fc�R��Z��~�q�{��c?������8k��a�X��#pϝ����عx���Wgǣn�>>�ũU�N�:��fM��ZX���Ɛ��n��i���rw-���i�I�:Q�I�ꤣ�ۧv�;���f�쁟x��f����������K�>x���_n6�^R�շ&IB#ã4<<B�n�X�G����j�QG�!�������-|���߾��R���0Vk������O?��ַ�5�̋�^�E�"`�����;��ٵѰ޸1�F�Z�_xEgueoޏG�����7K�������Vk�\M)�Vo��Q�ziBy���Ki7������m[�o�pPk�{���#�of��������ٱ�}����_�һVWWu����~@�F�FGA����q�?��R�#4��s<�(���E��� �<����ё���O��ݞ睽�;�i���-��fF�o~�����wT��k�~� I&��j�Y�{ �8����8�Vۉ�eIJI"iH�G��D�F���U��T�6��BJ{1EY���|��eOg��������ڿ?ڬ�n	}�N�����O���G�������y��V8��Z�F�f���%i���'�ݰ��h��(����)��K;vl�����G~���Oo}�[;�y��k�X,����ۛ���W;�+���Z��C��ӬՉ�����9n�Ci�R�gD�Z:���*�*9A���B�P����B��-dݎ[���w������w�zæ�ZB߰����?��ȑ{^��������%����:�
ժUJ���!X�A��1�(������ ���TCڷw����7�������[��i���-��fF�=W�viJ�����Vw���T�<
��</��R��R�J�B�j�*a�(���e��=r�u�lN��x��+�6�w�h6�Pmr�����7�w����3wt7#���7�Տ|�����ٛ���/�����ų��L��� `2�s���l���=����5�G~�-��]
=����������?ʲ������+�qQ�k�X,��?��փ��|_>�t����l8.yY��r�#/ȅ��\j6��Q"������!Op3,u���$�����9u��V�>-P��������=���O\�����|��Bz�%�w�������w�g_~��_�����K��������D�B����,������v� .����4M)�R��>�۷�c���o�3�����i��s�X,/6x�U�<{���r]���)#?w�͉��ʁ]/�eD�j���:��K��D�,�c��s����рet��i-�i���ر�C�����O���~��6�w��y\�w��ɗ}��������%�v�]��ti���E#?x<Msv����U*k�Vk��cT&�#7�|�����;��ι{s��Y,�	���y�!�u���־��ڮ�yLr�s<j����s���pS��$$��%�QF������r9S��!�yD�yD3i��S����[_�?�<���ߺs�B�����%�H}�C����W���}�痗�����<�5l�#!øԉ�w�2g�1vt��sl=��w�=��s�_w�Gs'�����g��X,����q�eeZ]�^�hu��r�Y�E����P&dp��!N�.wJ��ir�PN.��8�����E�C+yD�U
�O||��7~0���~�onN�%�;�W�}�=���7��?|���;[���$D�K'E�EN��[=�2c��2
G22�j�V�L�i�P��PFSS�����:��?����fܠ��,���A ��~��7]�v?X]m]Q]�x t�J~��/��}r(t}!t�B<�iBn�P�'DyF�r��a�t�F���Oo��ʻ�,��[���7�w���U����⫧�g�x��{aqq���F�^W��L�:��Oa��ek k;4H(� ~��k5.uKc��Oi�Ҏ�;�����y��>���}>�޾�"`�lF������{Ege��*���յ���0�Rin�����1�����DX���3�',z�jCM�}�]���U����5�}��;xՇ�;�񴄾ᮾ��?�]�+K?��c�޲��4�1���qr�sy�`q!��Zsq��Վ&�9���n�j���G?��ݻ�i���#?���&��E�"�|@��_���������p�\>�&�="G<�<
ȥ*�����A�|c�sR\ڧ�?���+VkT�zڧ3���c_����:������3���.��XB�p�n���?�j���?}����j���E�A89[��p8����@�\���\7��@�(qjjj�S�\j�+����g/�c��"`��X<���#����V�L�ً/�r��|r�G8��w�xTɉj~@հʄε�ILiң,�8���2AX�J�F��a��O��(�~"ܷ�N��;?��S/�5|#�'���ˋ������7Ν;S����h�N�6��덼��� Nð�A��a���0Ls��$I�~��8A5���O�����۞:vt{��A�h݊�u��t�cy�ˉ�NF�R�u���V+�2B�^�G���vNM����|�};���fmM�����X,__�?��_���]?������l���d1U݀*nHJ��jw\
�\=��[���	�Q�R��;p��BO<��4���
%�������v������������u���'�~���q���_|�e��sWy�ߨV�^�����z�Vk��뵕Z�������</q]'���4͢8N�2I���̧>�����ɓ��8~,X]]u�4&Icn�
�\�֘��~H:,t�������ㄺQ���&�[�md���?��?���m��mɑ#G�݇��o�o�ݤy�������:{��"`�:!p���|ۓ���������%Cb�)r��*G�v�<�8�\��~E��a��,�'�0d�{u�I��P+��\{��ѡi�:���u�����_�:]���^Є�����'�x��O<���N�<wv��OT���S	���x��0;~�wrRǡcK�I]�M�<O�4���]=s��%gϞ9t��3���@�v����u)�v�8�
B�{�xi@�2��A��G�F)EqB�z#�2�e檫��������i�$I�qw�	P�
4|w�;9�Bs�[�<N��R�AQ�u����q3|D��s�R����7���#�����=���=af�τA�����'~�O\׃�#�}'�<7w3���,�r'pq��q�����+�*F�澏s��<��,�j^�B��$I2ǩ�A ��Y�xcf�w%���#�gy�V��;�b���O�i���	��{��f3�WL��f3��t(����4�qF4A��˼O��F�$��W*�n��a������6�8N�Z�ɍ(�d6XI*~G��J߭T�<�V�8�AR�z~���aZ��3�O���Ĝ��N-
�$�yQ�3�&�*���[sFhd $�ݎ;\8�f�i�y��i3φ�s`��EJ�Q~���:����:ccſ���FF����Y�m[�{ş?yR�;5��O=Et��~v?��I��9�ٽ�hf�sv��8+�,���r/���{�pN=D�_�޳����A������������Pz�?�xݛ�������۩�O�����G�������_~�֧�|���k��8!?�($�W�������S�2�zU�
�^�=���I�2]�����^5$X�,���*��mwj�c�W^������G��;��n�m�5/w-����s�^��t��Kë�ku����FQm�:�D�μ�?���xs.hB��|`��<�{���z���J����{S����6�HRCg7����Z7�˝޸ѿK���477G�������.3Q;.,oX�x����˰ y�}�^�܅���|��x~�1��M7���h4(NR�u� M3��\�����mh�ߎ�z�k����6J�z+*h��������2(1�Y���Y���`㲶ĝk��q�����u���Z�n��>�'u]/v]'�<?r7�}��y^̟s�}r�8���	��u<�}�M��M�e�U%srJ0���g8]�!�C�gP2d
CƟ����%7���O����-�7剓�^��yJ	9_W��x��n�'hP��'e���p�Y��y�e�ɜL{��ż8�2ש��a�yy�{�V�#��
F�qJ>���xu�1Vn4�⻮��bʠqey��oQ�u27��I�nF� &�����7�t��qC�'�XE���%����Z�����Q:	��5&='��8f(s��}�)s3����J�<2�P|�r7ry�GIVz�e^��~7K{��O �s� ���uRh�Ne�������x��!�Hn+��I���EyVp��e�<��y�zy�BP({�K��b2C�2/��{�/�o�*��K=nU"��G�DPh�����7qB
��^���u�A/4���M7�`����n�����Z�V��jf�b�%_E���c�#�����yi��*O���<O���?������?�s3H
����g�ͱ�EeD���$ͽ�����^7}�翭��6���Fqt��k���,aK�˘r6����ݎ��#��2��}�m�%�(����۶P�wϙ�ƫ��sǗ�����=?���SE
}��n椕0�v:��nw<��l������u�9��_��>������C=�5��&��������N~����v{�����C4>��j�bR����<�p�$�_@��s}ii�ff����4-�,Q���3X��	<汔�y��>8�Ԩ#�.�h��$��8�������8]w�Y�9�_�y��&v�5�|1��'	A��9��`t	s[�xt�B�prV;�+�n��1�������$X�" 3�$����o3	*�I���@R��N�h%89��4|�g�^>W�]y������P[L�*�xL�P� N��q�ͤ&��s!�qxG/]��C�#��.��;�'t����s���H��Kf  �.MS�P޸er�ݹs�3�u�3�l���xf��>�C�Riƥ�$�.V��IPQ�,��Ô����q�NJS����q�1��ļ>p�y�)�0�y������L]g����d�06\�!e��BL�{pN�_p��-Q��Lf}��U,<s'YE�3�3K)ŸL�b�7��s>r��V�)�b�(���Bc�XW5+����CCI���;�oV�Y�狐-�:��z��8</-��8h��{YJ�����ۭ�����.�{#0%|/t�T $`�a���v���c�u^�� �p/y㭮-�#�8.^q_���R�P!�ϡN��,2�B�N k�����m�[�?\!V��͑ֆ��s� ϓ0�� �C��Xmyy2z⩱�ښ?�$ɍ�v�:x��D4�!�-v�A}:�0#�B��2�yc�;��R����[�P�oWwᢩcg���L�$Y?k�S����h@�3�ìl��2�yZ��ϧg�e��KQ�Ry|��ħ�<��#G>�U�vA����ް0�����W��ߏƚ�&:x��GF�B�~`�(���"���lH�%�:pqi��|z�,[��^���st"��h��$����*��7T'��kM�E�[^}/`B���+ٓ��y]��x�G�k���VH�����SbǺ����=Y�Y>�nג$W���x��Z3�_�{�7��9*6�c���W��x��jx�� ������m4��|�*=�0_O��{�:)cDs�����E_B;w�0�R�eԏ���0�C�+}YF	�Ɯ3s�G;LQ� �j���VX��<Fh(��xM�Xe�����m�)���YyP�x�T�}F��g�4S<S�Y�3���a��^-��o|=���@o�\O��9(��"�(ا�$��1���Ƈ`c�sY�$���QJt���e��Ɂu�$�:�"cY�>�9#+I�Z�߳ց�R���F�U
���3g�gO��ڭ+u����3�?>��� vv�n%�'��(QE��z�Z6��UfX	���L���6Q@�&���t�F���(��e��{�P�r�
�hQDw�������VP�i��Q��w���j�=�TWV����33�?
����*�L�>\?�c��������o���2&�������IJ�Ne��n��xc�S���N�R�CHH������3��K�K4^�����fGF��p��e�����Ǿ��o���}A�����?��v���3�/˲�1<<ʄ^�7Xi�a���pA�^�Y�<�1n�eܸ�i:{���-S���Np���q=�צ8)M�Nr"�����0��]���1&�fs�	\,~Q�E����H�$�X�懖���d��D�L�(�^!G%�@���0�	h�l�(0J��)Ut��T�GBk��ԋ߃�l[�����=����OdaBI(=�H�����y+~eBR��-f&69�F�I7�p:|�vM��{�j�iye�VV��V�    IDAT�r�k���C^�����AE��h��ϡ�Q�21N�
"�Xu[����������
�gE7�wu�R��]��Mq��*��1���=气!�8Ix
!ּ(�Q�a�9蹍�,��`�3kӬ7!_�p�0#�� 
iAX���Lه�w��( ��XL���(7e%�9�ќ���`rܘ�����ao"$�iw�\�+���?N�<��9{��Q����n�41���='b0l`�W΄��-Z%W���Lw�5�JRyo��Q(��*p�.FQ��(�P(��H��D�/s�>0�c}��Oc�{-I"n�Q��1
�����Q��y��3H���a�W���a�� �s��[���J��Mj�%P)vl�d�M��A��.�&�^��$ǽp��-�<)5N|ϥN�M����̳'1;��*�o~����W������� �&�����g�(�����q����-t��aj4�Xx@�2��{j`M��}����-\#Z[[���9:w���.Q��^�fBO�>�J�J� �
�K	�Rln<���S�ڀ����q�sv���]s͵4:2j樛&
lI�p]$�:Kt@�j1���\˳Dʅu�8�!���,Y1�N�~(6j�������U���7���]\��P�jF��`),���*��B�������F!�_�|���l`��7��C� o"c/�+n~<tm۱���Z��D;��_�(�y}�8�m*%��fM/44b����1+�si��Iھm+ի�Ʌ"У��2�WV*@P�҄�~$�&���[�ne
�@�{��u�aR��`!t9QI�>�{}���LR�M����,>�����q�Z��Ǩ�|��Tp]�$Ble�ŵ� $(-��3�������sY�pM�k18&K,�A��U�~&�D��z���O�L�?�7�?g<2���;��֤�dB�J_�җ����3g�H�g��֜��EARrrD�x���*n��>�>=w�M��^QX�s��X�ŚCB�/�N�J�8�G���=����a0�3&��B���]jt�T]^���	j�Z4�;b�F8�h,��99�Ȉj��;G���P`��Y	��x� \�R�W��D��벅�l�h�.Z8���<�I0}B���IH��<"�r��U�%�j���'�Q���&c�oz鍿sɁ�������q_�?^����󱱋�?�S��g��Z�W?J�qgǎ��w�>�7*q���c�]��+[�FCFfqi�c����Z�~�KI�Nq���i0&��@�0h�rp�qb{<�X�&B�c�8F�.�k����F��"��UJ�\J�ۮ�&7�FE\]$#�\�^I�pN������_vf#���@�݃�:��-Yz���k���\�6��.Ic����
_�l��p>��9�����z��y����OQ��@:�f�ixx�^��o���柳�	.��w{=ZY]���5a���N�4����A��v9�~���>22D����7�,������s���.0�<��(AbA����2v� ����gB�)�A�B����@l]����e�!`��d��~�هJ�,tu��Ks��}��-t�d��Tk�������*�C�A�f����(<-�_����������d�l6����=��3��k�|.�Rd��sBM��_śT�5��SR{���Ј�YN�5�_��� �0��_�Y��zO�`?`�1s#�V����\�P,�}J���T�{Tk�R�0O�3'��Z��$�� ��q��	s�������p������&v�co��!9Հ:YJ-����'F��{'-����8!���8)�o��Px'��������yX�K\���Í?�����|���_yA�o��]���\���~�O������45�����Gc#c�%)�}h�pU�\Ņ�7����rc7��8��yD3�����S���@�.F��(�uЁ�<_>o~�0!���[.b������<��X}H�#ct�5����8�&!\�$��T7�(&P�%f�S��<67O�+\�B��RPv�o|��2֋Qx�s���E�$ߘգ�S&���K��f����WD��J�.��yB��%�����>L?�x*�V�d<%�`��$BOI�D��wgtt���կ�={����0Xf �N���kW
2�:jw:b��D!��%�<� �J��\j�kT���rGl+���0V x��׮�9r�3C��:��<�T��3�`���s��(�L)�3�x�A �a��Z�Pb��0U�	��ȃj��}X��e�V�QK>}vR��?+�c��s�ge�*���)Ǘ88�U b�j��rM�B<�h B"j�ѣG����ǏS����(2��C �y_�1pl��z�W?�rop=�����1�аGc`�����D�����f��Y�@Ȅ�5@>��L�h�a�9,�q�*������:E��գ>����H����A�А�S���Bg�X��`-�%�\d�W|��w҄:qL��Q���A���Cg�T��5>�y��l�u����������4;{�z�N��m��j��z��?�{wމʎ���$��������m�����w�����$��.�K"W�ϰ�MB/Zwb��� o,d�̌�wBRs�3?G�j��}4-��A��l��h�
����o��Lc&t?��CP�`��μ��2t�W����T�&aI��dK����Z��L��$(�JB�qC�]݋,\G�%�$�����-�ϙt�-�Q�)�Y�O��D.��J�h��Bb���Xl��A�-,~A�r�B�*t&C��BQ)��ʟ���_;O��ؒU��	���3 ��u��ݻ��V�Q������-,p����m۶��;\ .\X�p��XB��8;�6�[-��ܱ�v��i����iuy��e�V�~�� %��<H	s&<��Q�׸�a��"�416N�z��	X�%��iux��!��j��hq�W��(��p"�tppXh�&
�t-!�@IG�b�SX���=�=���3�d8���CC�
kʒ(6/����R	�P E�Dɚ���a!�������l�q��+J;�G(ΒY8�ѣO���E:��S|?E��3NdW�T"X�0�ǵ.kQL�"EMy.���07$1�R�XY�)�_�>ϊ��H.�$QD�&����G5a��+&m���é�9yPT4s����S��	[���2yss�=G�v��	J#S�&g���S�k&I�j �0����t�I�U<�"�$M��
�>���A�.����!��*+�\�n`����#}��>CgΜ�ť�t��h��h���/�~�'?9��F �����r[�8����Sg�_N~@���<HI�ǃ���%���rL�%6#6-'���
ʅ�ϝ��y:&���<Ȕw���US��Y�bӪ�MX�� x�= t��&'�+.��&'�J��*) ��ycH��n�"B���lD�@!aRxk���ֶ�w�r8��D��ͪ^.ۃK�7��x$kڸ�٥g���|�~�&([���� �a�4H��$I�� ��s+<e)J�Id߸���p[���nH}?'sr��IlbA*!�6::F���u�kj����Z����q���av�c��D@�H�C����(,av#s�:�m&�.�TȎ�huy���8�=곻�)ޣ$K9��¹⼪��c�\�q�#Oƣ��J�;M9��>���tʠ�Zq��\�L�o/�f�=��M?����x�`����^��:�3���[��y�,�n�(pL?�������5V�qb(	���"^\\��8w$@��G�*���l��ǬT$��\b�E������ez��'�bar x[�������
�`!ֿ���ZT��C������(��ޏ�2��+�>��6L��`�ּIޓ�G�<�/��3'�&�,��]b�Wӄ3ڃ�%���ɛ��F�K����-�s<6���U�ݎ$9��E��1�y��������(���͐�R?s��{����}t���t/&/"חPP�cXC[����V�RX	���駏�ٳ���P5����{��V���q�/�K@q�_�g$����yg�o}�/���3�k���e�_I��?@q�3HB\E��3�`��I�P���+�Lss �S4B�%ԇ��$=�
&2�a��IH]�g`�C����q��������凯���mT�7��!%�}V�WK�֑� ��ҙ"��et��d��O�l��m/
�Z����eM�Q�[�8B~ nYwA` �W�d7(��+���,��/,`�$��'5�b�AA�\*�R�H��S���A�oPcD����\�	�w��>
������k���O�5$V�:[nqB���t뭷���.j4j��q�^�V[-&x{$C[2�{=4�%�"M6 ~��5�Ԭ7x��e��n�J	�5j�1�&��c��w����?���3�Qb�4q> W|����qA�n��Kp�CbPF�Z��ZRG�h��n�>�=6�/WK$	---��������n������Yڶmx��%I|1+�Zu������!�"�� E��D3)�U\7�V���w(	��47?GC�C���?�nC*k���Iz�+�җ��ej��)�u%j�d~�"*{S���TU�&aQv��F��x�$q�H���-�t�ҿ��_���o%���m���=��SD�{Q��QIZC�G(��>���c����-
��34��S���ÍNY,.wzP��W�,w�[��C�ZJ5��	_f�Äށ�ͅ��S۩u��t�2z��''"r>g��5H06^P.̘�!��=�ԓt��Q
|�v�������7�����򶷽M�ȯ��$�����0%�O=v�u3�K�7�Gi��K�}���Y�Ҹ�I\���3lq� P$��s.��hn.�Ӝ'�Ljy�B�M+��M-�"�je(�C  �^�t�bLr=N�By�NvO�n}~�V�)m���>I
��x���/�~BjZ֣��Z��$��,�r���>5�F������g��u��'nUd��6��AҒ(N_W�E�W���l����B��̻�V�&C<�P��;�pUP*jҷ|k�S�k.�7~�w�˽�JZ�Ɇ]���9�*ʍL,�XZF��$7��������r#�S�$w�k0��G���evE��"a�f��=5�yJ)���l!�D�fmI���AC����f��3�%|&���r�ܔ~��J�ƕ!;v���y�����[���u��kS,}��W�U}x�)�PVR�b�?��Ϟ=˟�CI�����1��B�Z����:�
-]k��Bެ��r�"�[���6s!J��Ey-��uv��x�Xy1y8e�q� л�d^>n��y~�Q��GB�!ԲD#g��F�QbP��Q�'TMcj�z��/�;=K��jv��L���֐�&J �`.F��"4t(�g���ȯ`+�/��=�K�g���E�J�P�X���۩s�:��L�W�[�,�h(J`291�/(��'��'�x��~�vO���7~�w�������Ο^�:r�(_�x!���W߶7����|��k��:��\�IG۶n�Sw�xP�#�:�G���:t���MD��9�A?��6��&��T�\o=%rN�E,����u�^k6�����l]�v^Kդ���er�[�)e����0Z�FW���U��S_����(6�qq��-�r0�����dyɹ�K\�W��u.�;N��d KՀh���(�)]��P��(�)��=�ЋD�U�n���ȶQ�B	]�����C[�l�׽�V&t(�P �"ַ'���"�Ѕp��o�9+T� 9%Bs&�#wpt��M,uC63c\N��^u�����ϡȋ���t�d�K/��M$���!	�w>�����s��(�cQ$��������ƽZ�Rs��V=�
1��|��/M��g�����.��u�ax(��~���k��A��,�� f�B<+��1�����hvv��x���|���AY���k�t�3U	E�+ӥ`�ka �:�)Ǔrٲ�o����UTF�A�JT��S��ZGov�x�C52CC�x��1�p�'wf�ܳ�T�^��n��)^O�]Te	�!�
q-�R���NDY9P�"G{b�7t=NVFH��QD�(�^J����6�]}�����AX˫Sw;��6��C�U����T������䓏���4�ڵ��ox���,�&��;�\|!|�b~�$��nz�E�,S�|���+[��ޫ����o�A�z��~�3A�1��L�h= ��4�KԔ'���M��3B?s�]p�v��$6ZXP s�~r]3)��8*,L��`�M	�����]|�~ڹc�FG'�y��kSk_�p�����R�j��3�7������D���V���n(���d�K�3�<s����Kq�A\֭f�n�⚸�)�JU������Z�VU����8PL�G�e,!v��B�YO�帙\_�lX|FKu
�H�E	�����f#�~�7r�G�x�n���� ��|�-��FB�Qr�QK�a��yR��Y�B��qL��3"�>����7�hS&�}I�x�)KG�J�{TA%�.���%t����`A�P�xf�H�E��I��ۢ!w�!-�y������㵂�&6�%���&�%<�*�>�N�(+�8�$މ�a��u���r�c5ju��nu�7��������Cs������!��|e�I�J���X)$�����7Y�ſ�äT��5n���^V�uo��F�W�#�Wك��h0U/���^3nފt6Mfe}��M)�"���F9�3�>G͙%������*sQL�\�c?��P�	���j����LM!����z� О&���n�O�(�N�I��(��2:�=��S�)a~ 渇B4��0)[�R����'�ӱ���;����o���i�7�zם�/&9��c]�����_q⸿r��S7�u�/{�-\���:�d ��Gn��I⃰;���*�:^��iv�g��ͦ�.�*��Ee>�EK�nhB�ֽ� �Lx:��HW-l$�wO�-[��X����m��,�b�oa���.�aل&><�ٕ���]34�X��� t-�ᅏ�e<�R�֥&�a����fZ��U\d�� � L�����Q"�._��b��J�J�b�n�@�X�{�^��7fƯx��L�8cIq#�ԸpÎ@�~ƹFa�DKI��R����p�K���z ��
�p	���DC�[+4\����X�Gڅ�P!|�Yoi�9
(�D��h�BtR��A<�O�%���;c���4c�梦�ĎK5к>���{���t�9(���f�-%�Cߋd?M�ԤD|7���e�����2���A��oQv�7�"'
����s����P��8Zk-Z^Z���e�5�;�xK�J�(�����6�H�_a���/��IE��U�T	��
y���Sɍ0�^x���+v N�a�ͺZ��'�i��?�I�w��=��0Ϟ#��Y]\��~LM�A�.�<�
��4<>B5䐠&n�Cy/b%eg��́��TkԨV����}�v����ԩ֨�m���q/�c�.�C�o��L�/+��DG�;≄܏���f��}�}�&�n��o���W^�?��;-��%�^v�7�'����3/���/��F�FD�'9�Q?w����*����ei��1�8�q�^:F���a�k&�����"1	Ma�tY��5B�$�<����sm��!��Eb��{Yb|�d-��N��8�x�:=HDSPU�V���ȍ�.��q4ḾU�6�RF�dn�g���9�)
K!�8�]j�SN~�M��_�9�����eF���R4�6�$����w��ʭY�/=��ŨP��w�Rl�[:���B�N���B�����M\^����S����Lf�Mܴ��`���P�d֝��˞
�CҸ6�e��Q&��qL-USBg������^�K$Mc	���`9�K]��Ii'���{bb 2�5ܢ�^$�C(�b6    IDAT�j%0]o�`,����nuU��l�|��:����2��}� �|I��Iɤ��4�%�G�,�r��z%S�P�{�*-�^/ɲr*����}[ｒ�m�h�G��u��uًUx�4<Q�e���Υ��O�͎<x��v�112�`������iQ~�9����J�F����?�=߅TѲ5�ڮ4<6L5T"$99��>�Q��t��U�*�
����{1�� �ڕ*u1����鸗��n�za��0�8�I��P��#�:��Z�U��Oݍ�˟�����w{���|��"��C��~���.u����N��ܯ�\}����ER�7��T��Q�
m�#y ��V�ck��Ytifv�Ν�/R���R �,�$0��P?���i�z_�D!��(=���S�@���U˷Vi��}�w�E�}�.Ѩ3u���+sS�nb���b\W��Z�<W,VuMn\'-�r�Q5w!�"�Y&6.36�+f���.��E����/�yZ�����]3پB�災$&�	Pj�p�B��Ӧ�U㤪8&F�� Ӿ��-<���D9�^ƭ��
���8�'��,��}�	PO��������lH ��5`��> (���l�ͬDH	Qh���9��}箺�`��w��nz��k	�����q]�|���VTMq^���u�{D��J��9���B���0�A"��W{���9��=��*�7u�@�b����:2	y��P��~��|�(hBh��w�l�R��dU�(Y�JE����7�E�g�Ɗf.������\/����RiQ�`h�_]��Cgj�z.�5`�\���2�RB-0P�I�(l<ٙ��ET��To�P��)ʟ=M[��4'��d �:&�I��Ps�NU$$G9�]�ߔj%��2�ڊGaU2�ѡ.� �Q5�B� ��+蘛��N�:a�z�G1��ԻD�Y���xEخ�D)r�����y��o�+�㿰��5���]����c׻&�^vŵ\"�ٰ���X$1��U�4@��\� ��� ��0_F��OY+]�ʨU*_:B����1����J�:t%}4�`�sl}j�ڷ�ڱc�g�r]�Xw���m�&MҘ�zY �0��7�B����/P��q�xf�pr
RU������,��')BU�)��X2k�E��F�w]���}tP-ø�?1�@6h���M2�v.�&mO�%k��%v&��VGًQ���z�
+/ՍU
��(:�qa�����ɋ��VrP��
��A�X4H��1�F8An�H%���{�B@����(�z��K�]]�� 'kB�ִ����* ��$%T�I��6�>���Wpϴ;#����^R�'kǖ�w4H@�܊�U0%���e%[{�C���k2�p���Ic?�����"�K<]0q�#g��\�=�5QԻT$��I�0小�Om�RV���_�Y.{^2d�?˸ɱ��ۻw�I�C��xτ��P��h��%�Cׁ<��d���x�OL�7$3Ԙ��
y�:�Bd�Ch�Q=�Rue��gOR��i�l�4�r��P�O���&9K�j@�(H2�vD������,���{����c�Z���&ȿ�r:�$t��F��B}t��7��Uo�b(^S���u�}�'��c_�F�z���?R	*��_�s�Rڋ���B����u�K�>y��������t�����Io�ν<.VrƱWuY�[S�LA���P%%�M�&̔Z�e:w�4�9{�-tX�ju�Mo���!�4IF]z,ܹJTh�&n�ϛ�F������];w3�qƵ�<b�c�R�$&����+�����F�۰L�*H�o]fe+UK�=eR�c�d���f�iee�}�+l��0��k��`ҝ[�Z_j1�1��e:+���v&\J������Z�b��/���C�`)9Pr����T�S�(g�;�\ӯ�YE&~O=7���ek����e�YpkXS��ǖ��MWjߩnX��R��:L�#�Ib�צ=���4w�Xx�:�}�-U���ؒE��d�2y.�d�����&1b<ט�$����k���r���J�#S+Z~D1��HlY�W�.U�������@���\Y\�8�	�I�gN�@惵3��P��,L#�7*�8.m3%��e�і-��l���L��;��9�Q�t.S��KeO����E�僈"Ө$ȡ0yꃹi<y-Z%!����P��g(;s���SIRj�b�K��>I�����h�J.��J�Bfaf��o�IX�v�IJ�4�V�B�m�T��
:��t��J�0d=fP�eĭ�r�2��qOwC�(]sݜ��Z>�u��_����_�yј��!�?���&'��3���8����S�^͟�t���>DI�P�։ɰe׺XI��A����\$!�D��A?�\L�+�t��3t��3����H��!PC�Z��VB��/ھlv,.Բr�8X�f�4�r�޽��?Ŀ1�Ef�K�.\��,%�@y��X2�5WPE�X��
��f�n$��m���c�1Bi����,bGkĝ;w���$s2�ֱ��7�I��5��TL�SW��]�ZCr"2�!�_��ײҠ�eu������!�C1�yJ�&h	��yp7@:�����[����n�I޿�-�����f��"�+�j�`�`���	z����3^�Rx*��FӃa��'�B!nFu�r}�q�b�J���g�멥�mG:Oq1�v�G8c��1zUF5�eW��)��{h��b�1=Q7V$H��Z�� ���\KC)3�؂��^VR	߇�:r�s��X(Ju9�}+++�H��T�Y֐1J�꺗�=f�Z�s"��g��]3Jٌ!E����-.-�W���_��h^�E	�y�'1h|&���U�����y�TF��c��Rp��At"x£'��M�RJ�,�z�!on��Ϟ���ڒf4��3�A,��\J�Ǵ5ף�/��C�&���q92��sVV�4B�AIS��)�~mUC�M�Q����l��3�.�|�Z9Q�BNi��T�<��e� yɮ
|�~r��J�����wN�@~�>v��/^u�E�̓��^m����O-Ԫns�^ݳ��J��ܡ>6��89���L����&&&iێ�TC��҄Ξ:EQ�MIԡ��z��'�ر�f��ch����@�����F��%i��k�̔�/�s���A-c�v��E�^N��]BI�Ӗ-[�,�u���}n�u������[ɂ���&	�Ҥ<w}(Q�5qxe�p#��ߥ%k��8�7���E!j4���*֘ڌF���ר*Eҟ�p��]]��ε��<�[@��z+�ہ9w��_�x�r��b)j��,Lv9gH�7GʈT���[�Y��N~&��S��^L�~�j�+a�E��]ܝb��}QV���4�ֻl)������R�U��^e�|��`���XLR5�,�-|%1��5���g�e�q�\���qL\z����&)��_P�4ɵ��%J�$Hjl�G3�3�5��ײ�Z�����>w��ky�K���A�����'�/�������g��z�JG���??����B#�� \���A���5���|�|��U>�Nk�=u��\v�0�ؾ�FFG�'�nc�M�����0�B�JZ�yʉ{�D��1R9Q�f�� E�8!���t��`�����1�j��J�sл'O��SOR��34'T�\z�����D@�z��p<��!���>�{�H7P#O5�_�c��g���Aw�ܡNR46L����o��4�����U�F�rR�!���Yl*���#��Dp�R�ill{����G�4��{��k�П�j���@��I�э�(;��n�N���)qC���^A �[�\�0<2J�[hdh���U�u�+�zÐ�ǿ�%Z���ng���M�;�qt��e�K�kM@q9�M��H��F3y���\I�E6�X�a�J��w���N�G�\r�.;t95M~/�	b��S,./�{R7��~�+���mĵ ������>H2+%���h����Q׋�z�������zb���L��J��5QJ��!)�]��}�!��cuu��{���o��o�C���K��e@�1�Č�Z�(\���tZ�-m[%@��˹��A]����s`����)����b\e�=)����F����b�8ȝ(�x.M3�>12��ِ-�\FPʱK:��eHG�0⁘4��J�L��s@Lڌc/�!�r�]�N4��3��Ӝ�����s�·XO��/��yZ"�d��k�]�8�'Q�Kf�l��>��,��O~�'�8p�]ግ�"��J�Y}hi�*�xH��'�yc��v�[[[e��Сôs�.�>!59Uۉ��H��RB�.kc}��,+Χ�<Bfi.7�bE�G�K���U����P=M�G���F����;Jk�NR%�Q%M)�ׇ�u��<�����Uj«
�Ɂ�t:��14鿀�r0�*Ր\ߧ]:�1���P��Fh�K�z��'��l�C�Q�擄V�V�J��^_z�sސ��uo��4��!r�q��.�q?��w��f�?_B���_�?�鷲(yi7N&��2�FǨ�{aH=���辜��Q�Ѯ�)ڿ� ]��brr���>�=�=--,���O��}�V��s�v[���|���)1A�l�L���b�p	�{^�v"$�?�&��A���T�:�]qŕt��h@���7!���O<�� C��)�~�U"eYA�I�l�l$��-,��e+j=q(��z�7Yx��/���5�uz��o��	qkѰx�j�g𫆘T�
���w�SO=��~���J>�y`\&���l߾��c�������D��Q�^��"�&0�Nf�լ���R��.�s�l��gBWK�X��7�]�c!�=�>�o�ٔm�b�L$��Z�y]��X�lesS��V"��T(����e�J����Oi��D2�E�)��	ܘ�^��|���_�)Q�+�~:&�A^��r�j�M�Dt�b�j�r�{���+��B,��iv�����upC��f5�A�a6��{?s���`PBCj=J��T2���@��=#<VV\�(7,����҇7lyi���Ү]S���S��Jb�$�i�+!;�*{�ԓU���$���8r)GC�~�(oȫ)��!�������!5��ZO��F�+]��}�YjO�!/�q�� mz�q
=Ĩ�*�!�dᾣ���`(���M��J�
�i�@�Z����a>p9[�Pw�Ng�u�U�5�@9��)�Ew"�vzܔJ*0�}�l�3��Z�ih���]���Y�R������Nqϗ���?�;ϲ�Y]^y�R�}�30�v�ʶ�M�<M dFʰz��@��j���OR��`�s�A���K���?ӳgɯ{����*XH��o��С=K��i�J k�������>��2#�c�Z���F��Kѡ��ht|�]�0�MO���S��C� ��z�h�,�mo��;�D-��b�����_�d�����ן?��C�I�W����l�@L���"d4<��%�Qy��,���1�駟f���C�$�c�[��s�.?+]��$f/1q���R2�E�O�z;�:��/���]^�H�1�pSkHs�{��%�m���".Ϯ�D�D�5�c���*���A��aB�&эɍ;$���w�J�IP�d�.L��˥ٵ8jM�����f�5NmH����]%p7��l���UEވ��4�%��t�3]��`&�i��R��M�B��R"]r����e�S�Ӧ�|�˼��Y�8.�������D�y &��=&@��V+�/����/V�ò�ȑ#<	��5��	}�֭�#f�O��C#Ʌ�{{��Z�l��׋���q�H���L�ŚF�C����蕷�BՠBQ��1�:���
��?���LyNYF�~���G5�(�^5c���.�L1��f�\�
�4�1Q���^�HpF�ȼY��^���($g�E0�<�ᆯT�\ң3Q����%{h��K(����t�n�O��������R�@�^��	���޽�?�oy՟QJ{�;~|���ٿ��.���o��y�%������7��p�R�R�^�r�n n�.Ō\��
���V��~Ef?7�T���9s�iz��G��3OQ�g���9$5�������jϰ��4g�se�j�J�ŏ��e;>�I���W�9ܟ�A۷�k���_~�C#D8 �,tL��]S"1;�|�%$]�e��׋�`�5j}�1���Ȋɀ	]b��>���8q�{з��[n1�Ɍj�����DXn�b
�&5�5(333���"ֈ#�7xgii���+��Rf��6�Z�6pE�z2�P/�F��
�u�j�����Xs�-Cރ��B��-{	�q�&�������8�Z��[��\��s�2�d�R�Ou�3�s*��3jŖ�W�+�e�{��_b?J�){4��z	_���|4�X�Fy�<��E^��PeQK��\�|���k\��ɴMni���mF���'�=��O��F{�c�"~B��N�C)Y	۲�PO����}н&�\]����{�Y����S���Au�����ue�-縗��FLx=�P���
+����k1	�<�r��n����:Ǻ}��{=ꜛ������3��4�:����.��R�j�#��,�)��+T���r�F�v���1�M�jB޻�On-$�V����c�C�Z�ڝ���z�G�z:uh��Ӗ�hە�)��^�X����SG�q�K�Q�41�hrr�����u����?a]��WS��w�yg��?Z��ސ���'B�c��ju����͈�ٌ"�� {=��H�9��)ʒ�	t��-46:B�ZH���8��x���>�_&�$	�;&k���*q��y�*/'��=Zf�
6�G�X�:^Mf�m�NW^y5�d���47?����=꯹�:!,n�\O���#龕q�,�&6���w��^k�-^/��D^�RCC}ꩣ����:XJcc��җ����D�������P�K.H	�������:��%o�K��C��S���o�>�(y�oq��]Ky�*q�k0�*׸1v]�G�����"�,���>��f����3��u{����{T�a,
@9�����c���.exoLR���
�����+��ȔF�I��{��נ����eΧ6�\'�����g����a�jU.O��" ���[�6���*Y碨��A&���P�$ck�Gy-�_J����֝K��*$B�����������Ō��X� u�X�w�a�׼�5�FmY��p�ڦ�X���>�P >�����+4S��pE��q��6�=w;zK1��<��\ꊎ��^����������C#'�X�C��QY x�=����ɇ���:=�3�
.�� �^�q9�>���jD�[�{w�������1a-�r*!�!��^�k�����B+�.�
��)-�	�jM��&.���z��Z�R�g�1���E��.w$ �����տ���~�g�[��|	�W�^r���=aP��j��.�C3�K�QD����hTh簱Q��7�o�)��4;;�s�!P� \r�y����~��N��f"$d�c!+��,j����T-]n�Xj���`U��d� �٥��Q���Ϯ�Vk�����׏8�&��C��[�5��491I�e�% ��|^��Ll�\�z�̥�[�KMR+F��.��i-��T8�I4a��юP��g����nX��_=:E��B�U&F�$ũ��E�*IF*�hq͘���:6�7�8��/�qe��#�1򼜉�]�$�X|�ߍ
�:ׯY�,�4��D(jq,r&{��e#J��se�����JZ�Ŗ��b7�S0+�c�v�w`T����&&��Ұ��+)��1���9s�2̴�$M֮v�� ��Aݯi[��.�,Jk\	�h��9>wyθI�[�����lL+bͦL>����{ Kӫ:��o���RU�UK�-�������}<h���61��&�V�,�DG`�hF���0x���� A4B,�GH-�[�R[֖�{�2�s�=�w�?_V���	��z�������r���;Q3/���LO���G���AH���Q���:����    IDAT�l���#!1�%ʐ�Z#�6}$!Q��B��G�� �@��������� S�J�{���5B3�����Q�V��ȋ��DP�r��HF�Q�r����lq�
���g�}�\Yi�/5�KW��~���i`��ᰙk�ZCŏJ��K!/L��4�a3������p�[Ͱ���<=I�X���������5�3S� %é�fl�|���6��7��+����Vs��[8��e�^�p�r���⾅ߺ��M�������������,Oס���/�{��y����K&Lﺳ9;5ޜAF�=�z�c�F�����x�\�x��������g�.^h6�����%�b�b��9�-*�����]��� B�g3���[��!���a&��'63@ݘ$����k�ONB�+ �AO���q��'>��oR�*�K2������jd��+\Y���Qk�k�`>�}G��a`��uS���N��EEB�.z��lC�,$;�Y����/0� I��_�����x4H�Vt����%U���
�I{�{�#�rF���R��\���欳�i�.ƶ]�<[�CL���*U��3�R!�sڒ��m��2b�i8}�.�	�e��}�~��e�w�Z`�Mg� F��� �cW����:t���H̭y�U�%i�y�]X��%�6�㜜���8�zg(��f�|��8��Ҁ�|\L�g��pBt>(Mx��^��B��u�AД�7�@��1&	�sfg��%�W(<�X�+�DyJ�~��o�Cr�(����}ꝏO�5�h՝l��B�8j��f��E�@�('͌M4�S�>��Q�3#�:;�9��!�n}��"�+���N�XkӀ�g�1��H��f�fr�Y���ͅ�����p��l�6�,{���/h�;�>|��@��*�E�@���:&���'oy�D��K�����7��3q�۽޿���{�􁃓/��9=�k��i�4�M;���ə�fs�O��SO>�l,�0�]�Cw|�,dࠠx���a0��\!�t���y.2�Y@����1�����Q7F�}2㦅������8d�`�������O4�S�t�m�S&����G��Ύ�c5,��-�L+C�Y��fC�7$�!{يA-=��{�$5��"�q�3���l#P�U���ĢkPpb�3��'HrO>�$Em�%Q�.��(�9y���`Dp����S��׍{�*����Fi5��{���]�ֱ�C�QS���qk��k��+�x���?G�W��[�������n\=4�q(D��2����p^u�y�LR���"��p�u�c�4��� ~*H��RE!��c�Z�L �y8�t�2+�\#��!@a����y@�AKg��:��ɓ'�,vg�Xn�3��p
TL8�Ņ.h�'piPn�������Od�:�1"|^;�܏�;V���s�)8�w=���v�%y3�C�bS����J�䓏7�j.\8�l7�f2�=���9Xu
�ۇ;�[Wc�N3ݛh��&�E0���C�]z�=�<<7v Ё4w95�M��h_�:=7���_lf�5������f{g��p�rs��������z_6W�D3?���~�I�B5A�K�=.��ah�:t��w�~��~�}۽Ӈ�t�}/��/�nv�ω��/n��.;Ҝ��h.V��]�a�5��,����xsa�|�ĩSͩ�nVVW����������@3�9G�q&�3�W8D���Pk�X�P��M(�m{zV��y�cz�^F�lg��R0۷�����[���߿�����L�=�Jj�l����E}ё�W��M��=W�>_.X���h���K��֪)ʱ��'��`9�f}��XGv�����2�A`�A&un:X�u=�J0`U����ͣ�=Ҝ:�ϟR������E*��Y���6`�����ɧ-g����9"�Q��4�iz�b���l	�D�+%����"C���q�h��p�L����z�,e��%�!e��l���'��!Z�L�*��g1Цd�!�R'U
$�d���6T��}�f��W��-qt���9���PK#"ǩ.E���\�5`��P&}�n`�� �c�'����"qV.D 	�6��c}ab�1����â��@�ub^'���H.E�@�W8���%q��.�ˀ�V�E��T�-�%��d�>��zy�A�_�C���f��u������6���hΝ��7���7� l�:4�=Na��7������F-��q���ش$�IJF�/�
��fs}��o�4��9�ʜ4�u3B��LL�9�vn�?��A���?�~Ōd�(s�u����|�$h#Ȅ y&u��D���������׼�[{����z_�B�|}�g�o|��_�3�������[�=0�\�oVPSق����!CF���,�4�/]h�|����l._��E�ۢ�? �	�����pP�]mO�X��E�k��c���Ln������->��PԢ50���P���� �����ѣ�m��������fq���6`��}З9�FC�e.t��Jv�X׾l����[�ڣ7ԙ)�Yq���㊲�k����Z���ǚ�Y糖W�|��,C�2>�%?��	�� �>Z^|3����̌jp�&�*��g\�Ԍ%gVv >OT4r��%ө�����5�@��g��a�3%2a�,xr�_'��ڱ�E�)��*>$��$?�?#����N�#g��i̝�|+X�PЧ����0;p��ۄD�2H�� �욺ї���2[9���K�@"0�OC{}�Y]Y�vL@�3̔y�O����Ns�6 6Ɲ}p��ް���qp|�M�ށ6�^drZ����蘃.\����#��9C�>���^}5�Q{.�4��|�y�7�ߜ=�D��Z��e���(y�"C��e@���Gm �M!7�3$��t��� �GaC��'�&�3Ǜ���nc��C�5���q�n� ��a��T�o��拾�%��w��٢b�%k�.`���ɧ�fg~�׼��^��g��=�c�7��_�ڷ�^������ҕ����]s�5�g'����f�w��0�ho��Cv����f�����SO6�|���e�֛�΀ӓ�Ч�'��	Y���=j��m��59
N]�Zi�kh��gj�����^U���!v�k񨟣D�6xH��/47�tSs뭷5/|�]���<��I8=�	R����D!%0Lm�U{���"S��$fq&�(���FEJV���Z�4�q|������1 ��Z ��Я�A+0"	��(�]�8ئ�\QN�?z���\��}�����fw��p��/�����Xzf����^��lܭ5���v
4)z��� ���&b R%�]�D&��Q��a&n��R���]�t��}���"�4�BF�^�$����}�iZ3�0��D�9��D)
$Y[�hA�.�/��ū/���2^�81�y˔� f^%3��ɁW�7�5��Lυ���R���c2�2���ĸw��u���2��De��>�x�����9b� ��q
�XtP�7x>b�O0#%w#Z����XZ:�g�.�#G�4��@�-����Ψ�A��@ּ�XA^ͥ�5-��[E��c
�� ����H���3$�m(~��|���ӏ7뛫M[Y��	������*F!��|X�LX��C1щ���; z6k\�<s�h�p�`��"a�~?5���	�elqV:dd���y��n�?�|�����7��XNJ�
�Z���孭͏��.|����?ك��_������/y�/���>��G�x���w4��7[Pn����h�'Xw� �'���W�P�N�3������+�����q)g������#ee0ʀ�h49�HF5R��P4��	IB�^�"�h�߁65H�B���[n�A�c[
�MH#n ��0�m�";7Ɋ������p��w{�0�:G������n��Ʒ��0B��*5�9��F-g�~s��e
¸����;}�,5����aK;%W��3�Ǎ̄���Hr�]L݂�?`R�j��mJ�����3@p���z� �m�[;t�(�����Ⱦad��9�uO��CB��	u5�����]x��D:��C�m{�k��~�p:hp\U�1��1�N $R<t	,fh��zoq}�����kP��ц�����F�"�bݞh�&u*��g��Q��6�$�����? k⻥��m�"�z����`j�kv�j�r"�cдJ�r�D�I�I������rs��y^;DM ���i]๖@�{WCD\°��3Y�� @�
�]ܫK/U��:z�H3<�֎)�C/���s�G����ѵ��R�O�c�p���UM����ڍ`8 �="�3l._��|�O��9}�������*�Zj�I8����G\ZʘT��rt_0��gq�6�1qP���C����8`��N"8�l_ܮ?]�/��³��4w����[�h67���)d�
����l�ŉ��꛿�[��ر��_�?ч��y6{|����_��͵�o;�����-N���fza���~��&"����~a�9�֪K���J���-��
KVґ�6*�[C�ц^�I#ep�2%	V�~v��0�+��)�X��hف��(Pqۭ�����bq�¸��dsc���[�TKS��)>'yN���������*����0����f���:o�
K�=���	���c;K�Ԯ�Q��F����3/����u�����8_rv�{-4@�~`�'�{iy_^C�&����W4���0���T�J6r�vJ��}���ʽg��X�w�n:=K��=���� �H�5��|�����q\���6�:���*����~b�R6yR�Τd�q�pLNҙ��}���9�������U�R{�	��s/���B�X�V�����"���=h�\Z�����J�Fx얰���b��X!��C6���� �Q�!�;շA��D8�.)���^����_�cN�F}���r��$�V^'�����Ψ���a355�����d�t�l����
��ZY�.�Jd}�Q/�4��L����: �ӋVТ-��F��*���߁.a]�`��珠y�óN������<�U�I��h)�DNo\���꣏>������}��>p`��~�O}f�'���|]g�����'Z��_������^o�;�s���;�� �!�W�$4�b�F�U'���_��%f��#	]�$[�VuOtm��s��T�}Ջ�+ŭ�K�]F
5,�*é����InZ���Bm��U?���w	r�M7AJ��$Ţ�f��~�t����1d3��z.3~㌂0 H !�,,���GM٫Y��	:[����P��)�2B4ä:���x��t^1��׈�0s~��aM���T��'c���g
��f�(��h�����"�]���9	��<���a�r�b�`��_��z0����a�v�X�����5�D��M����_�{���$�\��~��~آ���#\�3#8;�|-6�BT:�C��r�� ���=�3N��G���?�A�f��YE����cN��ܚ���R��	jҢ1�@�'��\�ca�sZ�8�q����[R}/)�KC������9NR�%��	U�w �bK�Ą84Q�˙������;��l�+yP���M�!�;�ʑ����������� 8"�,�4n(�%�ԍ�9�8.x-�=�p��|��{ss=p��i�_m��5�|%�`�T��'��G`DG\D�D�4�I��ɘU��]7��� yR0��>;�����5�4�kaa�9z�&*s��	�/2u�=XoGk1z��ͣ�=t���}��n�����r�����^t|��{�a��\���o|�������o=�OΜ=��驹��n��w��-��Ha�l4��q��Q�� �.ş��&�#������M=���M^�7lj,<plr,(X����>Y��*�\�"��q�H���b\1F�]�$�89���-�Ƽ�f��){�e�`wC3��ꋚ��f� �
�5�A����#ŵ��L�7����ls}��\()�l��$��#��Z��cʲl�|�Y2�Kd��C(.�)w�_�c�N�Ԍ-�J��^Z���jp HXN�N��aP�w�������;۷c����b�N+q*�?�}g� ���
��k�����m|��=@ůc��g��?��1홙��l���C��n[K;���>`�a�r����Q�BIt<Ϗ�!G�n����d�L�s�F\� �P���N岉 \��H��G��3�7A?�����.�����wk)�d:��a��`�$Bc��A:���zO�j���w���~�ʭ�������@)/\8�sR�A��{�<��u�]͝'_�{����j>�O�5j�_x/P'�vA�*��7��أS�K��JIHrAfó%�	J)$�*���pP�WQ��Y���Q�@G����(�2���5����
�**�D�DB��aBT�� ������B�\��(z�1�k�9u���S��'�&6n�������^��S�w�}���9��)|�\}�3��W���5c�y��S�p��ʗ-.do �G�b#��N�bUә!�Y�/XИ��Qض� 	�aa�O�\#H�߅,���6{U	=YS�-_q��l���'Y4������NM��
P6�G��z�V�٘Ե`0+�ޅ�$@��� G�B�j��<7ծ��Jk�W�6!:Y9t��	*b6:a� I?&�g@��X��N���0t��ݐg�89�-K�0��֦�+;W�'������������Ȕe(�U����[2����0����9_���d�1!0�58#�q|��<8�g��� ��.�Ӂ��F]�Q$|W
�[�WC�>o;s9'1��8r�㒃ﯹ
9P�{��<��hM�&[�'s�Yf���;hW0;#��R�Չs�g Y�0�8���Q��gg�G��3AT�`F%��T�B+��#�$4�o0�нv�3g�Z�_�����©�/����|�@@��Γw�\|�A:t�5H��М8�}���~hs,�vs(Μ~�I�JnR��蕃�&�ϢD�ܯ*�Jx&K��P��GI-.CU�P��^R�$��M$2BpPƛ"��,?t#��9QS�ʛ��&�j�HFm�B@���N�h�n�3g�l�|�T����8��÷�~����z�;����Y�u������ao�-W��|y�3��'nmn��f.��m���E]p��ɭ�C�]��r`�3gg<��l���ke ;#Y�B�!����6<�L�2�Ap�[^��HA�Ɲi�xD�ز����%8F�Ԋ	[²ָ-j�B��5l(E�8r����T��io� 3�ݫ�~�A�WYCƃҼ1G\2�tG�{ �'j�䫲�*�"Ǥ�U�YȊ��Y��aP�H�J08ϑ�>>�����N���TZ�
n2�#���|��A[�#;h�I���Od�t4V���[��p`ոU;w��AL��0���3�Y�R˗r�,q�V��F���ENS����Nq��U���ȵg�BZ̹��R}����;oΙ��/f5�8�M��¡4Ϊ����Rb�k�{a��.�8>��t j@�����1v5R� JY$�K��a�P�'�+���1A/P�DMY��
*]�S������\S{&�cՋ�M7�0	�1A��|	</(�=���&�B���A
ˑ*��=H�._�L��Uj*D�#�0��*��)6V��R��e����h�y�_BP��M43�3<?�?QR�����	����R(j��I���9t,`��h�I��kC���n�\���橧�����C������/?j[�|�y];����_���~���ڗml�T� 䍛=ͩCgΞ)YI�΁�@�7�9    IDAT� a!j��#]��w��7_#����[��Tg᚜k�6H�\�Q������.�O�hUe��o��S=N-Vp� ��]+g/C��)����Z�2���vMR�vKh��*QF�L�N֎Z�f(Fg�U�{���_]�����������(S���U��h�G6���ʬ1�I"#20�0:�V�V���AP�'S]TuJiz�N)��R�,u�)� �Q_`�%a�T��1�ې�,�$)S����g������I�GP�a�5�m�W �g���Q|�[ug���ze�x�P+!OF��©b���(�X�f~:gղ]����b��%�������������}��"i�,~�7<;f�7��a'�p��pF@��� 4��"��1ja������J�{����"B���u��Ã!Qs��8�:�"�ɽ�886
��u{���ͣ6�Q(�����̖�%^l�:@�tX����61�������6L���1��N�j�$�K���A�5־x�3������§`K#�v�*OF$C�s��z�*H�B%!Kx~
�d��r�St��]����م"ۭ��]�<��V�/���/5���u�499����/��ß~����:�����_��_��/����S�X]]�{}cs�-S����*�p�*�0P����H��X� @`�x��	Gp�`�_�t��$��*9����qQ{vk�aC;eAMZ\̌�-t��{jAʀ��F�EP=:���H�Y����GA���iib㘥�* :�4�UB��|L]ʋ�%��bU�1�sQ-�Y[E;�!��A�BD�Z�T�~)��v�&'���:M��dؗ^8E�+�c��8��D�sIB��lm���+�TI��2:��|�l�筬��P*IO�hP�Oe�"k�wL}o�+D9��h�]���葃Vk&�P��%A���6C�8%��L��=q`��=;ȴ���&�c=�2x�G��wD��b-4:
*O��z�Q5�rUf��{RYS #����z�]��t���Ņ���P��ʶ��jYUg�P=C�5#�dc�7�d�w#�d0D�N�@�LT���4%�5á�\(p���:��o���"�)�E۬ߣ�� �r]�Ip��h?�?/�o�:b#QY�D��@ʉ�;%s,;潖��:��fbj���Y �X5����33�va�*��+�Os���/��͊��5hV�V�'�8�������=q˭���W~��7|�礝�u��z׻���?���?������mp�bX˩c�pX
��3Pgt��j���H*��{0�9�M�)�N��>���� �`�8 (,p|��ԩ�9�5%�S�:��H<���],p��h�P-Q��	8�n+���T"��]J��n���Y�bk�g)W����C�2�X1�U�z��Qv��;'��Z�6��^�(ʮ[J_4 �f���`Bx�DʘAΚ.���Isd�	i�Ʒ�6��A�!r�Cd�.�8(�Yd%5��NA�:4DY�k�0c���>@��ʁ�9<Ѣ���cz��ڦ���б�jq�5�ga#G0�DJ���-�[}�j�4���S�# Cӥ���:��D:�N�I�Zgp��nd����80"!�d���a{9F e�#���!@�:�I2��u*!�Z{}�B) Z���C �Q����^<�I��&(�l׏�^�:������=Q)�!)�-��\'��sF���i��P&�(��@b�aa�T��Wu)�h�Dy��8_d�n��Ev0������U�H�
�E�/H Jz��F+�`��qG�K.;�D��I�C3�qB��u	��6����y�)������2�ю��
v}uf�>��0p�M�j�=t�(K������s6���>�:;?�o� �Ϩ�c����C��v˛o��������'r"�|���u����/_��_~�����q��p�8K<H8d�s� �����4F�0���e����V��'n=��v�22�r`ߪ�a�7�[�M7��v��a�@ST���nCNw�q'892�Y1�e��b%�A ���nn�^�$;���-5Z���q����&H�4��
��Tb@Ί̫t!��h��4d߅����������ɚt�	�E�nc�ͩ[ٲ%^�G#;��V&N���]r��?��D?k�j�-�{d�r��0|M���Vp+"֐�32#��e���10D�ڮ�CʒD�`k��z�k?7>Ch8�o�.�TjR��,��G���ef�+�5���,�ܹ�4d�d��e���� Aϧvph(��BQ��x8mhYb[f���� ١}�8�K��-��Na�V��i�x&���V�ٜ;������c�cO����z~(�����H������'�A(����Til��8�h)�ZS��n(Ω�*A�*_������q�d�@�2�佥�+�zM��E׎�� �m����ĳ��Tn�1q�ާ*{��~�N�T�"����5MDC$C�Xh
��{�g��?�,�:%0��Dc���� w��Μ>�?���_,��w#������\�x�H&���ϱ.�l���} <�T��w,]��\�p�z!.��N��:�����y��hpO�A��{p���<��`멻�z���x��_��'����ˉ��^��5�y��?��oz������`pȆ��p����QC��d��P�]����8b�#�v�C��l�m�P��D�|-�ډ��V�+q{Õf;皷1��HQٹ��fL`k�%�o竒Dqf�,Bߛ��b�3S.s�=��}��vѯ�Ib1�ћ�l�d�xz��ȿi;�:U�PXߟ1`�m��Zʾ���F�@��uJ��!o^��z&�!�p�z�[����ߕ3t×Xp�0��9{�z]��Ñ#�EP�!!++�s���q��o��~�2��[�78���0LX�F����~�O�1�����1Yj����*����D�͂�!H��t̘`����x^�_�Pu��BI&�!�EP�c�9r��}^�zߥK�<��r�áC������}�^�����%� �¦��2�%�
�*K���v<����A��Q9n�,�~�N��!���~׈g�f�kR�s��|4N<O�=����	fTԽr�N<����^���N�f0L��+����K�}�3G@����	�= ]7=�>|�5{�ˁ M�lOz�˫+���Z��4IrX?+�����%&g����d�U��#����OP���'�b���	�h�\�~�ɘ�6�vH� q�/}�K�O/^�x�Çcvf���?�ܯ^;�������gΝ��?��G��ʕ�Cb4;Ԧ��e-��S��u6��m�O���p�^G���5��� @0&� S3a��=��}F5�ꌧ.����n&O�
�h[��lἵ�E��3��Vy�[�N]�����l ��n��M��o2�Z6 �"��o��%3f���Ѷdvs��md �=_!;�|v<u�T�V`���\���|H��%828u��g_�|���m1���ҁ`3C����u�HWk<�ѣGi�p?�� k�m�`��J����O�>͑�~V6�p�8L������9���s�w�7�pCs�ر���~�p�[�V�Vi(3"P���9s���9 8o@�8�[o�����̙3��o�.�3 �������p���!�P�_��s�9������#����{�<��܁��}�(�=8T�����ȁ!�י��2p����3r�+G��z�E �46#7�����"G�fy���ꈅNy����v��v$:?��ү�y��sR�������q[n9RܠR�p�!ͬ5"�]��&�V�xf��c�c8t\	d�Dlط>h�?��q��͡C��g�6�>�(%���2�g��5'O����p�����ӧ��z�k?�&��X���;N6'n9�`���fvvLAC@r�*�~ ��V����K�䋛�e����ə?����������C�k��U�=��7���������zD���7}n���Qz�����F�D,vPg1��f���`��uov��1�nJ�Ejp��D���1���B�4��NV4T��r���� ^��l�g?k��]^�:Qi��TU�2d�u�6ty'f���C�xȡ��� ���e���=�a'T��7�QT�+���}=�
�;SW{�&73��Cӝ���T�|�	�t����C�\���|ގ+���M���ϗ5B/���`|�1�횶Q#h���>\״�}�k�>�	�y�i�����̑�����y:i	�O*i5�a�ik���V��������������;���}[3cK��ɠ^�߅���̼�>��@#{ZD9���{�r���:B����Zsu�yr��/���J�zB�7<a�NV��y�����ϗ�R��h(=���L3٣���W��&yo��@��9�?���#'JUZ{�gqe�}L�dp�2�:/`�)�!6P��ޤ��,��}�+�l��46z�����!e����'��]1hKՠ��j�u��<Dp`xN�7�a��r�7}lfv��?�������z^�y�B�ox�ţ����>��,��Uv�iA��Wn��I�7N�D$������V�+��3j�SP��ZŲ��2����nj"�� ����[�`(p#� bYfhʯ���Zv��es��v?�j�֐�����T�������Z���w�$�YK�|K]��ھ����f�]�{5�H�><�zx�6���,�0FS����f}c}-��R�l������k��j�Z;����E�r�����L���C�������а��=�t�Ng�9��ʨ3��zu��'mb^��g?�#D#u.���B����7Y^aօV>�	;�A��r|�S`P��I:�t=�4E|C�oD�8Le�8{:�%���:�z�k��Yuj��cb�eW����j)�|kA�ڟ�P<�3�%ڈ�F'�&��vD�_���m��C	��|t���UA1b{q`8�J�֘|��r	>\֋�9��u�I��u�>�qI�@�����?�Ј1˞���P'�Q�
�g<֕	��w�B` 4��	�wǵT[� �_=v����ff~�����������v菝z�<��{V�C��z�:D"
@��\Dv��b�ix�-j�K�N
�C���%>��E��	�M�Еa�f!l���z�U�<6N��$���o�k��i��2���<�½�s��Ƅ!;�d\���B�@��H��K�[ٍ&�eG�윾>r=������q����zn�:bLq�iE�g�3t�0�	�a���Xv�v��cȡG��v=��=`X��O�kCǰ�L��A��}�uv@E�Q�ہ5m��.�gÜ�9�5�%|�Κ�nGr��8.�"���@���y��y�C��7�+�W�T���eޠC��`�ܜ]��U� b Hn��q�qn8���U��d7�%�	D$�p�z_�u���[Ӽ�]�N%'�.��� ��E�x����Z/�i3��V����Ď��5�Vک�P���_�5�;r���)�_�X�ߋC/μ�b("��������vT"��)�a�D{�
�Yg�b^�F#әr�y��k���U�&gf��
}�Z<������ǁX�R0��xJ�������Y�f��j�&�gi׸� �s���\=v�M�ufv��������g��U�N=�����Օ�#�Su�&c(�=F�Ѹ�A�ŀ#�,�V74�5v��zhxC),�0��[��jձ��1�,=U�P]m���S�nȬ�u��8���%���oUC��)"LP�'��L<C���iGRϧ�]жIU�I��(���<u���8P�AO���j�ϴ4_��G���zϠ��ei��㝍�*g��tu�Fm�Ӝ"S��:��n���z ������.�o������I���&5��sg�옰�FP�����8/�U�!2�o�"�TD�g����p<s�8g��L�s��P&��Z8��3E�s�RIz����q]:j��>���%2�Q����$�{��u����@���1t/4<�"/Ԇ�peFҦ0����]7��}Y���1X�L���b��������ϧ��,�\��j���i��x����Vl�<��Y��=~��%8���0���O�~ᱻ�s�QF�v�a>ge�8�=��V�`�v��(^~N8:����{­� r QL�����tꏄ �r8�`�c�Zٰ�pl�1]����B��e�Τ,���ʕ[��n	`�˸wl_<�z�7~bzz������������u��~��'������bmu�I�ˡ+���#L�d���9��N��$��7�Ա��KYʑ#���&���������G��j7���B��Ay����ECP2�u>�5�v-�.�Q7�e'���%���G��
=�3�b�:�K)	D `G�~eg��u�BY�f.;����Gͫ:��k���J88��ƈ�}�����n�<k�KMk�!����,^�'�����x}����]7�{�E�O����yx&;��a���p,����h��2�\NP��5�>�frC���=��y��iV�b���f���^�dB�W�ʡ�F�����%�[�|�N�������@�\���º}=n\
������
�~Ȏ'��lj��^�<fģ5C�1��ã>���Ķ�n�t���`�/e�yӆ�6���H[�A��{��'��r���]�T��t�cW��j�-����%$wF_�^s�hFr9�m�3s��w�g?%�ف��d���mD� �{�c��w�<��:�$��T ��Џ���G�>855�S��ğ�繻�k�u�~����SO����������a=(9b��� ,2	lV35he����eig�N���!A�(�"ḫ��(��l�FR��p�j'��iv�!%�a*�4S�4�A�6�C2:.&��9e(Ԁ!�]\+!�����wg]���O���{ҕ�4�=9X)+����<ŗel!p�.Ƙ��AAѶ����\�����2�j=x��a�2K|�5bd�h}qߪ��j�CK�֙z�-�	�����J�5t�k�Y3���oz�A���EkWv�m�>qd�r�Ȯ`��ޤ8C�X�!��Q��p8td֖yŝ�35R�kYT��;�L��9�'�<��a�:�0ʒ���sq ��f��Jl��AL�L'�&���Ɓ7d�g�����0\9��(Ͻ�Q���=�vgu� Vk6���x�d���]�m:�Qr�qD�"��'޲+/����,�}��Y��bh���8�(q�V9?�Q���6N�=֌Q�N3(`m�q�$hޔZi�#Y��)�.�8[��D00��#L������A�ʩMp6�Хt��h����5�8�����;>��O��������u���=���3��}�>�_^���v�+���)��i�VVզ@����2Se���C�	��	�|�ɪ~G �@�X�H�FFR]S� �CS������i��M�����t����4Ռ.�JT2D��u�u�7�8�l��d�*�"B\e����7�(�>ʱ�:����|Z��jＯU�֨�3&��*�#��4N�#�=-�������00�Ԣ3�Sá3C�F{L�C�d�0��M�5���<~�07��"$�?���}���q-x��n����G �5&:�tF��6V>�p9���"v�x�4��r肺�1_���Y8'���4;�}E��uk�*�Pj6������Uw��o�A��{��7���L�'�����%�i�ƝL�m�#���0�����U��{�mYm�'g�>��k<Z"��e�m0«8�p8uo�:8w��د��r]Yĭ�~����#��}�蓩IPݏ�<�K�ޮN�z?F@����v-�Lj���Q֤�P7�|���\c?���6��n�����'q�t�E�n8�f,PV��M��9B	��B�pz�k����c�*Al�    IDAT,>211�?�O�빻�k�u���-�~Ϲ�K���|��[[[[4LSZ�b�n��ʲT�(]�4[1դ����>Ke�R�b{��N3��N*B��Vd�r���4�]�@�!K�/���2%���\�~��d�יU�Ǣv7�Dio��96��U�*�n��ʆ��r���:��RN�מ�5uC�^�hT
Z���$v��~��J���t��g/U(��;�#sC&�<���
�����u8gݸve�r�8����DS��������3]���.9t3���C�wḨ�㼜U೸K��8^=���Lq- ���j�^��e
:u��J�vw ء��`��<+C��ǖJ����w����؄�x���#h���^�	�^#�v��]oա����mn0N�.�V����@p�����=��g٬�ڋe���sv裮m�c��%�����ͮ�@hL��!����=`��שsk��Be�Р~-A-�R1�&�����Z�yr�`��XP8��q�¦r��4[,Q���A��Ju#0��5d��/^ǔ x������������c������G��k������֡�����.]���?���_�����ȋ-ڜ��D��n֖��֠������S�Q��	�"	Ԫ��[I��>.g����U�<A��H�mk$N�Z7�E�����>���'�����>�	-b��F�;�Ԥl\z���d��Mec���t���\�����������[B�}��<5�,�)J�������{�{Y�#���Au�$�w�&fG�`9���~��p�����Ǒ5ۡùR�C[=�p�0١�V��=�Z�Z�U����f��4ezzʂ�༑;��9��r$j8\���t6��ER�C�=5Ɒ� ��#�Q���`ؿ�¬�4s��f����|LC�T/�nk�:Lc�l,}������])%�-���lw;��A)�^a!��гs���q�w���{Nw;�]{q����� =#p��+t���y��k�8�a
h;�KmC~��u�'>jvQv�\-W�4�'5����S.���('����'���?6.r+��g#[gy���5<WC��3�n81h��(��ȡ�9�k6gg�N�����O�z�sw��>�u�п�k��ryy�{>��O�����`g8]�[�K�ݬ�.��2C�!t����9a�����=�X�Z�Ɔ��tmLlx8t�[�3�N��[S���p\��2!���ۣ�O�Zr[�-��U0�B8r���A���Cμ��1qܰ�C������b�����i��P�8:C��&��ѹڙf���!ކvT�',�R���Ӿ�(�(�b}j2��6ft�:�4i�ݎ�D5���v;t�$˭���r蛛��ɍ���e�ְ�����C71/�6�՘���F��ύu�@$��w��!�.���+W0rX��_�8w��0��q5к�D:�(S��o���/��`V=�*�3M��Օeqg�ƚ�}�e���,�W�snwE��=Q�ے]:��k�� �k:;벦��}�@��?
��v��^E�l��hݶ�br�{��^L˵���9�/�� ���~V:m\/7�gr�t�ۨ`6
z_-�{�]�$5�`	��BLf2|���p�ak9��	 *��ó�>��iS�@-��i����+2�AYp��� G��8Y:Df�Ǿ.��4��9=5�x��{�ٳ�?���^��߾���}�y�/���ϱu+�D<(lL�VA�[R�:n.66��2D����U�S=^���\���G��(K*U�T}W����V�`��D�1�T�)6%/޴�:�Yh�����W��E���PW�\�ŝ�ץ�Ⱥٹ�7;��&�z�x58��a�������($ue�l�'tZ	Wq��=��fuס�󚪆�4�T�ǀ����"8�v�1����Ͷ.͐���,���:���TÊ�z��l�9E��D��q�����?~�z�΍�� �����Bۥ;t��1���E$�d�:8t!_c#:��2������^������x/�Ü�73�}������_mw�y��T��	�7E�bj�W�v*o�μ>���q{�%ya��]�Lj9,}O��G�f���$�b����7�5>Ra��I����AG����vC��ݭ��3fW���u�ԋ���S)��^d�`N�6�a��s�n���K�0O�m�8Λ��"����?@��ա�i��Sx;��B�5��	�B�ތU�N�9��5r����'�ǟ��zo]Z:�SW�����^����;_���~�������ԑ�]d;t��$^���~Bȹj��$�,H,2��bq�Q����a�2q��=��!�'���&y��Oe`
�j
��#s��M
NQ�yy��o�T��#d1����*�̣�P����dǪ�<D2]X]�W��.�>��X�5�"x���++�a'+�-�ԉ@�{���}�X���k_�f,�ܝu��[�/i�*dd����3��%,�8��X�ꊂI� z�qwrwf�ݰ��ia����l�c��@����t��Q�_����
���ׄ4(��0%��CƬ���yL���QC�r��:��*�ǣ&���TH�������ƭ�z=�KF��K�+L!8Y�C_^VPh���$�s��b�^�p��$ч��f����:ƻ�h7���b��>���3�XN�5 ��f���/���ݢ���S2�e��
z��+@dR�=Ʈ�f0��Pk�QȴE��&��e�k*g�� �ڎ��=�0~'D;����ڙ-g�A�x��$�C�����!5V��}@/ZL�n8��%N�=��x>F8t�8�Pt�@i����4&*��Nw8p-^�;�i��M���]s>�(7�����^o�'.\8��ώ˾�Q�c����^_�x�cO<q���&:n�G��h��a��!�A�D�Up�w��
[X�l!cR�!4|F$(;;�v�-�� �,c �R��BR��`&��Ib��x\P����Jr쥇������[��F�Ʃ:�vo�9g�+E�(R�Sr�'Mf�z-��v޵� �,D�'�[á{���Q�:�\�5�"�O���<�!��"hp��`_"�����p�fgJ=�lLnԔggI��5���0 �h���%�%���Hj��,��� p.p\v�� 6���C�5��	W�w����P�{8<�_��*���b��H�ނ��np*��`�&ѥ1$y�����t�8K���}6^�q�q�Z����С��1������'�8���!Cǃ�qDmB�q�0��0�߃��'�V��Z�'�,�/iBw_�Jcܕ�a m2���R�c Q���*�zrY�5�\Bl�h���3�i����K�h$r�P���wOC/�Nޒ�Sw��̼��d~ڿ�;l�ժ�}����t�
`T��|'I���P�Sd�x���Q"���֣�3�]'x/ed�*���hS���ڡ+aԵh�4F�hW`�Km��e��䨥n|�kzK5T��K�����C��������}����`Z�\�8?̒	�� .�u��! �>t��ݲ&���"3ౄ@��C��������R�8�{�<�bBgZF��C��ݪ䫥k3��=�eV%�Rq�٣?������������7�3������x�+vb����������S!�M�ɨ�H��jc��{43ڥ�u�w� �b��{��h
�&�$�m��ȓ��DnA���d�`6Վ'<"C�N�z�͊gr�Xhg��j�H�s�3���@�f$�ʠb0 \����=d^%g9,�\�`-�_�	.�D���ۙbzU 6�H��G�~��8������� ͣW�=��e q�T���@���3`�9����˼V�Nr`Q*\��}�} [>�<dHS��
Oe7��!([���Ee�vO�{�=�}��eiA����i���td&j��V��n�2�Y{K]�е���
@��m+���u�pާ�L�� �Y�K�G5�o��t���'���ǉ'�o2:F;��WL��M�v��ɊL곶<�|a�M-�|{�$�&Lf[�*�ĳp��3'��W��f�i��r���C?y��W�[oX�x���)�ܹ��dhS�`�P�F+[8uz=H�x?��٩�<�80B�k�a��.�/�#�& =Ùt,��������Fq�IӜ�����jv��d>+��n0C`�ш�"H���MɛV��ӣ�wO����cm9`�M�C���,I:jɸ�Io׺4n	�"á�9�?��u�I����4���)��An��S�2��FfZ!�5�� (�����?D��ʘɷ@�mr�ЗW����ҸZ_x�*����D�)@�"T�>#�4k˫t�oG���o �B�%���6_��F~�6A�׸���)kl������u v�X���*h�`�C�NrK��^1�]C����KKʆ��B1Oh �/�E6@&��� ���D�y������ǹ@�$ׅ������￢�uӳ���^�>Lk"�#?��++���,�E �a��p��P�L�\DU�z�)[Zsx�"ޒ�u]�'"��o\=�=|��i���]#M�6[9@r�B��7�����C�aܲ�}�������� =�b,�B��������Tt��w�;�D{��6mw��m��Ϥ�\o��d�?In���?�=�LVK��4q˦9h���;�;���^x[>����9�z���Y��O�v8�����흝IGZޤ�U��X1��A�{r��|�䚹�8����`�O�� �,w829Sioc1���#�O�PHn�')
���'�c�o��YT���/^�}Z���L��HK=�4t��c����x9�/A�~ݧ���ʻ�%�v-/���w}���$�X)���	;:�@` 3 �<N�Ņ�R,՛3r
L��}�I���g�EBto��!|%���YY
�6����v�h���3���ㄒ�@�Y�݊g��.�3����@��q�H5M}�X/p��g!n$���Yf�h§=[��N!����$��1@EC(,jG��@X������N���N�����'	}[>���'�%A�����d��O��mr��|�1�+����
�'�J�{�-}���k���\�ߣ��C9ZBE�T�83|b�叉)u
��s��P�c7��d@[�hF�ZF���p��	-q x�����[�&�E��G��	�w&�^{�}�{sM|�b�ҡ������ɞ�gڊ�p5�\<�ӽ�m�(�u�}�o�m*>�RBM(Z�U*�1ӎ�iY�@���r��:�������]��|���8$�v'����o�����~ߓ��[[[�;�;�j}�����>�]���n{�����66m�~(�>oF�\8hl.�|�ԫ��h�q��F}{�Y��Is��Ǘ�W��Y6����B�ȤH���4����A��}��$�y���\1��>�t�0�Ѯ=Q��rd��}-E�i��dD�-49�u�N�$�}��������w#2�"�d46,|���R^�Ds�s�a0J G*�1C窉>�����z�+��ƨ=&���2ζ��Y��c�)��;�����]�َˡ��GlYb\��/��^��� ���R�r �����֨�+��lW��2n0ȱ>QS���Tl�7{k��LMϩ����MJ��c.4��i����&�a���&����:�������9�7
x���,PR��w�8��&���8�$�E�C�18��̢s�w �0����F����<���v\���}l�k����QHVEuЛ\&�����A=̂R!�����Z�k-�n�)�_-D���*䝱�������"e[!�n���(�r��u{�� GN3�7�;ja �bU�C��sggڌq!b�g���]R������2k�J#p�=������2
�?����A�L^�ܸ=��*!�����[��o~Vo���v��7ml���&� �d�Sd��IR�����}�H���91� m�Qk;p�@������K4
8��R`x����;ԉ���Xd�СCEJ��E��'9��-G�VU���"�~����.9+dYt�$ęeG��[�ۿ��`x�@ql�v��]o7b �J�?�~�ؘ��e̥֭Z�
�����áW�ސc���V��_e,b�M��W�\U(�f�S��P��o�3�P��]�//_�sD���ʕvS��Ft��Ȅ7�Ͼ�L`XC�+���QLtJ���1�?�,[韫�z��\Jq���`����D�� s�|w}��b��J�]��-2���Ԩ��o 8�x�=���u��3�6Ŏ nE9�������{���z��Ǚ,r�7���!�w�gt�=�?��ث�0�rG�&�FɊ�#��߷�ȃ��,��2XC�@*��o�f�_�l��c�`+�0g��C-R�6��F�hĚTD�i8x�m��h�{]f�:Ȩ<n�{.��*/l�D}��/&)٦��G����x����Y��M��;M�dlDr�,lbv���x&p�x��Z"H��[="�|�¯	m&}�<4yVl_S�ͯ���{k{��<a�� RT9ZE�m��^�������F͹}Vn{�]������y���`a0���3���?��P�¿�!?$��l�ˇq��?w�la�"�siH��"AMs�"Zi�;�G�D����;v��8{�l�݉�\��I�52�v�
�'ֿ[���2l��l� ?C-��Ӌ�]��0�������m��P�ځ!g"��31��@g�ᣮX2�N.�U��X�he�ٵk�]�:~�2^"T6W'�x-�l4��/��cm!Ѓ��+��v��Ç���~��$������]0p؇"y�Jl|��=:����+�R�'��8��ǅS�3�ls��}�Ͼt����p��A A�A���v�f�GU��D<��\�ia�9|�ׅ���ap�GnM�����cGad��E�9��;{��%^XZ�6 ��$��M7�(R[t�`���._�����¹�s����*{HD�׈� ��|��zG�w��ҩ��A=}�4��R7,���@�'*oR��dFόD��f���/�C�?^P�Be7J.[Bٮ�K~A�����cזں+d��J�[�赂�k�nh�&$DC�\�k��#Pщʉ��4UeK�������+��m�R�Q\B5mM�p�?@����&Ӷ�V�`�S4i�9v�f@���Z�59�D<8�~��5>1�c�}ϻ�{�<�N��s�;;;�w���?�C�|�p����p{jk8d���I1�ȶ-��Eo��V�~�ф�F���A�\����������󁻿�2���\{��[���¿�[ʄ(nC��;±�R?���%%8g��p��l6<��c��8�v'�Ak�WM�\���{-<�� �p�:��n�?[�|�_B�2$*5���F(N��z�G)�o�z��OT�fu]m��[ ��n5��kF�L�}�:[:�D���"'����d�"ߺ�I4��EZ\�^���\�1�T�v�`/_���Cmdbnc?Ȱ�|@�a��n��ﶲ�s����Ɵ.-�;�&$K5h<�̊����7j�sa�Y?d6��b����~������atĭ~G��Y�Ǆ��X�`е�BGl^�k���|�
��;�^K	j�I,����H�h���aG� g��p<�C8���I�O-�̑�s���v�q�c١��ζ��|�t�	t������9����Ȇ��"��v��ƭi������pvn��Y������+w7����`ۈ$LH��(.]�C���-���Iu���ڵ����۳33o��_~߿������^��[��Z7���zt�c��k������hm}�M[�;c\0�ؠ�QY42���7��f}m��t�b�I�5�qEt4w
��=�0?��Dv�L*;`Â0�� a����?FCaG������yV�{u�������    IDAT��Yю(���d�3+6v�!7��3i��Xm0���]M@�
���q���h�	�Sy��J*C��$�PƧF�PHD�l���s������=�� ���%�7���;��2���.D�X7X�/�=v������P�����I(}}������r�y�����yg��o������^����sݹ`F�^p^Ȁ�,����D��46;��H��=�>7;U|?^��wF���j(�=!�,�8�!��F��%��mx�j�)�CP� E{T��=�r.\�0j�Zܿs�q=̅�Hr��.��5 �j�,v-�\׿�
�č}� 0:[�Zڙɡ���d���l3�|X��uۡGH�	*�j����yl's]���K��|��^���i!r�B �X�P 1࣫%_�%��{����5�@��߉��5���� �t0w�2<��ǟx��_�+<K�_�ds��Q�?�wr
�vb]���u�y����ف��7����g~�߼eaa���_�r�����Ρ��}�?x��·|˽�|uu���t���T�Rϰ6U ꘒbV���Ǚ���6t���u�����~�zDH��D `�i#/�v�@���ZXW�!3���q���Z_Zvrvt������s�����^���.�v�i�C-�v����{�U�	�:��K.�cRm�i^�a3��u�cwo�����88I5O-@�h�R�]�����.�u@\��Y�N��mvl�N׉+�!x�ٿ�X\�3�G��%#Y��yθar�3�SNJ蕯�u@��,.��E��B����#G���8:P����@����'��~�~�|`8�b`�"��y�r���Dd�Mr��� ��D�h{K�-]G�Rj[�B9����u��l��D7)�T��F�ުe*���ҜY�NH�2�]_���K{��^.9��ڨ��z��Y�_�bs��5R:�T(���ّ�il�E1
��&��]ܣ��u�X˧B�Μ9�J�Fk]����^�!8t;�� ol4�s�����T�il��x�������#���?��u8>u���>�<�\w�����ŋ�C������˯߈�҉h�_"�ؘ��6$�Щ�[�1I�N���,	u��l��ܑ,����T���#��HrXr b�;8U�v]E�dU��&����.G�2@�fs�]�������j��g�'�Ya����x%�cm���vC@�?y3R ���K�(���}���XzZ+�����@6Fd���\N���+����Ձ;s�3���g�q
22��}�\{���nׁ�� <?����Ip1Z��1�'$y+�ڶڥ�UN�W����PE%�$����n�� ��µ���CqS���U�hQ?_��W�"♋WE.1�a<���+B�zVp�R�װ��K��x#�����AA�dȇ|nՠh�-b�������d�Z5�L���#�Di�"vt�-�c������>�Ԯ���gPj�yEW�I�|P�m�����,��_��M辦��|o��C����ˁ���!N����S��$TKmx݁1R�w�ۥ!<��
���.��`���XI�S�A�J08��xӍ���o��w������^���]5��_w�}�{������׽�~`i���ױ�K�n�<g��~e��_�c���!"�6S�q����!B =�ԁ��$�P3��^�+���ظع��Г+�"{�-�}߆�
lV�!�]
:�T�����h��W�.����M���@Gy=Hs������|�N_Wι�x+�z�.�8�8�%��8	�m���	5�3j�2��\�>h;�U�!�]�:2 � pv.��"��-F{�ʱf}�;�[(�-ȪD���u�H�ڀ������D&��8?8M J�l���x#�=���Gx?�t�|h�w��Y���c�E �!�]�t �f�?#0���V��@�����C�O @����P��{'�}���U.���8v
�D�ړ���C���w�~Ȁ�5�<E\I�`++v:4�S ��Q n�P��Ё�����
q�e�2�5��n�|SIw.��B��ҫ�Ѽ7�Т��T�&�����uוt��lo�s�Yx�/Z�	ż��[��y�].�:˨�nج����	�`��|�.I�o�cCe!_oj�I��~��֜�#�	<
��9.�!�8v��]����fcc����{Ey�~�K�>����7���/-]�~ȳX��P�7�F^X�Ĭa��t��~~�56�l]���44̽��\��eK@�5j��!��t�2$4^hUS�!3�uza96��1�f�S#]�ֳ�Q�Vg����q]��9NO��N�%�4�F�-��c�)Q�tIa��pc�+�B�đ����)��vm�����%xSW�8�ʵD�s��a�� �3S
�b4}G�B��F�G�{U͂Ã�a��)}ྺ�<���"���*�%���A)�yuZ��J������XN�����~,�ں%Ǥ�ֆ�3ᓈ�f�n(x��I�|�<� C��jך�ά&�"{�E�R-M��B�<T��x%���N��y��y
>nEդ� 3dr��Mvr{��촻���گqP�T��i��?��(�h�1�K��,��Dv��η�xVD�;�҉Rzn��6�s@�$��̆���'~�{^���`�?��?�"���s�9�w������ȏ��ם_Z�^lD�b��E���Y����xhy�va/&]8-ߢ���Ǒc/������*�ޜh�ژ瑢-��#{�T��.)vy�m��m��5ס{�4`�x�C.灢Efj)�>��b��矉xяނ%}����дoN	Gv]Z��7)PɎ!.(��5���<t��r�~d��R�0�?��hMӢ�Sm�ֲ��i]�q�f&r�P��j�Ջ�g�`!T�&�I��|��г1���5�3'ðcUZ/��S����Gݻ�Ϣ@���uƴY���IL:�37*�]-��"e���W^�Rj��,^1��ܢw[̻�n?_acő^��9�lg�3j`��Y���"�u�<��@�������1�M��(̤`��(g�<:�m�F}W��ڗa�§8�2�	����L�~���_�����������[��OӔ>��=];���l>�w������-����={��?�Q-�^M����� �8��Fv&�dǟA�\,2�G�7�9#o/�6��۲�݈��jT�Tz5���^7R�H�
t��M0K�_j��G�M�����r�]�!�w�nn=�JjI�u��rݲ\Qa��Am�nW���N3�������m�$kZz5T׺t��_]��:m�!wV�>�ݵ��v�T3�jW�����-�5���s]=���bE�`�J #g�z��w!ʓ$���Dw�^�9�&�S�\���J�T���$�8���3D^1�
qs-�ى����� q�ih��|� y ��|����w��0�|w|�ZB��Ӳ%�U,�1����� w;q�kc����V�^�J�s0�q{�" �����~�ZF�4��r0Y�pY�eU��Q�Y��L8:�?F���ݿ�]E�d�Á�	a�8�hm�t�ǎ�e/{���������ܞ�'�}����>+��ٟ�ٙ�`�����5gΞ��g.)Fz��a�?|i�3҉ǆ/�����н�eD���T����f#d'?�[�	��<�s��K�Z����m����=��Q5���X��c~X]��)r��J������p*d�2��p�,��m�p�k���Wۘp����I*��]�|G/��h�ǳ�����]}᛽��N��G~ߕ���*�w�2�ܹ0���]mu���6�B����MY��]��IhAEÓ)*(@�6G�9�
�T����>w�Zq�~f�"�98Ѭ��7�s���U)QK�E��Џ,��@����`��V9N)�؂�G�!j�I��	�9F��?*t/��יI}�����s��}֍��kq���ƭ�H�3�[w�ڏN�����$�3���馛?��^�����=���+?wv�������CO����׷o{�[�5�Ν}U��d2Y���mܻi��j��5�b,�Q��W���T��nm�j5�.��5x���9�yq� �����նgy��.��N�v��*�N�k���^k�o��ՠ���m�Z(E���x�˄�n 4�����2t�S_3������rZ�\�u���%���m�s��'�i�\u�^�e$�V?�*tk��v���kGǈ%����{#�սC�	�����W��/l�9��4�j.1��4
�}&Я<x�!��a{��ݯ�@�]��u��);�r2c�A��{�0��U<'ۂJ�ol#��5�^��kWw[��4\�ȷt���խ��^W���92�>�������{�����o��S������[������5gΞ}��f��
ܴ�)i��?׎���C/}��M�7V�뵇�ƹ2��`�����0I(`2��9(C��),�I8���U��>'fd�:�a�	����9���e\f;6
�X���u����A@���R+P���ihi�Vg�l+ñ�����Gg�ޮNb�� ��ю��Z�a��Q�ˡ�����l$|.]'�v�]'�3k?�V�8ØIĪm�j���z��:��22��;���+,�w��чN���@�X��Z�k��^���~[9����K0�Y�^ϒ]��ݵ���]4�v��np��E���������[e��9�hw��<�r#���{�޹ ��� �{JLh-�,��*!�L,��{��J��R�ì�����o~�_i=��<���q���=�`y>ۯxf��ﾟ�YXX��=�y��/���4T�B2��)���ăPL�+ư����2�mLۡ�=f�z�yTA�n����*�*>��5�Z�n�a�p2��#�c1
��Z��F�}�(��έ���wU�jL>O:��� )�E��>R�i�����v�m��We�8T��u�ݕ\2�XK�Ā���EAL�J��m��g�{ɻ��E;Kq�{��]���䯪\�HF;��vu\�(gQ2�0�<�d�S��rFEh�*�ƺ'G�{ܢ��l�k5?�����Nj�g���^�jf�/��/6��^�Q�F�6�[�/nR�r:g� ���A݀�ں�3־hۊ��rP��� \v�����M\�z�z�,>x��������G?���v�s��5��s��g�����m���w��]���3g�|���No{{���Q�2��" ���:�ˣ���������V����+*;�|=~��8��v���g�`��|c5�v�v��,��8tF��ػ�ȟ�������[<���x�j9C����Q���3q��6�7�(C�vh�[Fb�Qo�����n#:j]��>�lt��7팾�@������5�i��U��rU�@�r��� `���rVwO���{�&��y�uy�����|���J���
��]��s��;�Rvx���jA�7ب�K����;������ G��Z�W���C����d��ގml%+#�����S7�[��y��� ��777������L��'?�g�<�g�L��9t�з�'n{�����O����7����Y�$X=�NS�$p�q�p���HR��9���+��&S�,�.��H0�G�'�t��֩\.c-9F�R��ҳ
4jY�"i:.豭O瑝������味�zb���Q��X���z.b��)������䍅��u+85�ȉ�|��
�FA�us�^�m��A���@�<���Q����3����*��J�������{�Fow�ߋ�Y���+���Z�mY�h%����]��N�$S=����1�Y0����(�S�q�
)��gƵV��TXw�����������׮*�ղ~��wg�\����W!r�Lb魝8�w Q�W�`�^�.���{:u��wPKل.��^?q*W�]��ε��ns�_�@ܟ��:�S���q�>�a��|zz��1�������6M���O=�L�3}�u���ﾱ�n�m����X�p����S�~����8��I�Z4_�Jjr�p���8=]���g�����v�ml�p�n�Ni����F䘊��=�9�)�ܳN����H�`��F{Q6�4(�2҇�nG�� ��C�<��q�a0��zV|�P8 X�ExG�[=�:%Ǜ+i5Ӓ�nU-�)�9y�����uf#:���ෳ��<u��7z�-nw���Z�ޠ�#�Tq��n7nͨ>U�'2gI��S��M5�К�{���BuўQ�"��[�9<�����˽�v�`�{���s�J{D��Q�@ރ~.9��+[�]�������B'��Y�2���i�;'���IG�Sף��Z��vO/�z��s��J��ẜ�����WI��*��8޻x��:0Fߙ.r���ۍVU��<+���ĵ����r(�3ܲ�-d�g���Y:u����N�����������s����������/��'_���yr��5����/]�T*�������Q�9����J����p|��놳�%�!8Q//r��?��_xj�0Avzj:! ����@��#cegQ�m9�̽0�|����|���<��ğt��3�#�ex�7i^A{��v���!{�x�@m�*�hC���
z�s��cǵ�S�"��ؠ2�������{e�������Ɂ�{Z�+�b�%u�Y��ʐ��.��3�.
�[Nk���	�F�0ͳ�����H����C(k
��>�+�L{ �6�u�
�ŧ�e8���<�h�]�IK-0���G]qu����;�K�k�7���9wNaԚ�k����~w�9��V~�y��u�=+Q�R�琮iԥ�\�44�+�<�s�>�z��Iٴ�|�3��>�׼;,)ad賳s��鈓���366��SS[���}��^{���3r��o}�����{����Lk���<�SO=ٜ~�t3�p(�7=M��	O��1}	}d��m�\۠é�����z�­�"'�1S	L��5s��t��d�)��m3�У061Q(�L�	�.iC�zk�lx3��ް�"�I-t�kK;ٛ���	]���^�xF-t%�R �ua�iK$��@*t��j$јE��a��8�N�SK�L���Z*Z� h�YaI�u�[����85�(!����n�8���k[b.���J��$F�T�{����S����Z�Y��uI�+4!Tr��ZN0α���������P��� �p���NޤU��J����Im0S `��؟�1*k��g�M�mO�:��L��7U��CMTA�T�h�h�J�ՉY��Z���t��[�����4M���!-��� ���	�؋VAt)��$PPë�W���1��o��}������ex+�X�:���{�ߞ��|%D�\=gX%?3���./�C8FO� k���dG�h�9l\V��>���P��;P.DM�־6sKhEO&ɸU%��:7珲F���#��������-z���>2.9Q#�����0:5p���ꫯ_p����%������/��U��3��?�Ԁ���쪴���p4zq��l�:�z���#�9����������w�%�@��� e��n*HDh!�H*�"k��z,kIoi*���3����;�)^��'�T)�VF̮���;��%D�o��Џ��e��+�G�7����?RH��Θ���Eީ#�/\����FK� W ˑ�$ ^TG�*8y�*���Z_j��Y0�q��gVfh;(V׾��]�qٻ˹c��9��&�$y��,OA  tC���8l���<���AQCM���j#I-уL�C�n�g�A�	�����(�k|T�\�bI�6�<���8B�"�:ph�R�k����r'�1���f�u��b}��5KEO.; ��K&'�K�z�Md$�!��u��Q��<��.@1,�5�kk��/M����_��~������#G���/���cǎ53;N��e�Ԁ~��Ͽz6X|���h�H�N�:�N��h�    IDAT>����Ⱥ^�X�m���,m�>�N����V�g-.�V�O���M$�a�ߚ d������.�1��:	��m!3��A�}��۞F��û������x`EX\� �L(�`�����l�x��&�'�+[��t+�3ܛ=�Cao��vD���	�H'�[���U� -"�Q���2����֚��8�kcA� ��pG�$~g%�R'@�b�\oC�@�5�O�-0+o�QK�B?XJ�=�R2��:���IXa-��!�I���m͡����6��2H��vɖ��ѨU)ω�$��+9�9d�;A�zf����m��z��T�x�L{�����.�.���l�Z>[ߠ�����̱�$_���(�o����K/KG�\��92���ڻw�����w��.t�X�����.�ꙋ��ó���t���O��FxT��gϞt��Ҿ}{YKz��f�ƉGҩS'�'I\�ek��0��)'��x������iYa���<m��kR�)���(+W	�c��\���ŕ,�C
sPlL����t:����өN#�K�J�G�d!���v�����6�m���~~�g��&�Z�Z�uS���F��_[�s̽9ʜ�T�E��=�Qƶ�p���)vH�GhWhn����� `Q=�BI�y��V�7��I�yMT��T�]�EW6ˀ� ���ea �9�h�9z%��DJvl)�P�Bc��{��q�[�������U����
V%H��Q �ɂ )�j��Wp4ɷr�4�I��P���3��hn�p66z�c�����@(]�W�+z,�	FQ�c�l���4�ڑ��I�PH�y�H�=��2j�ķ��pEH�*Xg�a�e��%'5��TO�:PB2�N�t��Q628oq����`0|�'>��w?V��r�75�_x�e�\�?7�ͯ��{(f1Z[O����8���,��h��3J����\@1u��o�Ll����=���){�C KǶ�R���f�uI��B����� ���$7��X���K�_����L`�C:�:�y�Ӊ^����`(`��5�� ���6k�5B�"D�B�4����^�tjP��w�p��D�����t�x��ƶ��$�H��/N9{���{|^�&�QܨM4�)A�s.HQ�g@���<Y3WTD� ��"�R��KH��4T�r���_���T����_n�։�_ϊ� �L�����8���^�,:�U�y)��ꭒИ��eC�)�WЧ5�1�`=�_z�Z���~�BG1� ���j��vݯ
`e[�9�-.�� �(3D|D�*?�GG��<���t0R�)��@j@t���<��fI��%:�L�t�a�uh�E2
��J�'�Q�,�?��9�B�WYl1W*(�ѽ*g(�қ��(b�K�(���;����tL���m(�U}����*Y��������{%s���'i����l�I�I�^z)��	�N�x4mmm�p������������z�c7���U�Ɏ��+7\|�3�X���O�u2�^@�9��>tbH�r�NW\hG9�Gg`Ԇ�Y6l�j!����g���ʤ"\����UK0�"����Σ���q2T~$�$ȑ��.ހB�T��D?��EY��Us��G�R)}����,J9G۸��������p[�?4%x��u���a�r�k%
�<!?Q��A�OF(��V%(Q�䚔���m�"^���^�eE���S��5@���TwM�؂��� ��t�bN&-�g�ph��g(G��	��/!z�M�3@�3��=)]PJ�g��Ã΁�%�]TkK�WtD��.kJ�\���BN�������)� �NJ�c @�����6pҚ���Ӕ&^f_�Ea�3���ý�e��4����b��ã5YRf�e����4ˉ�!Y�&t� h��g�D��G��(ͨç&��j�)�:��҂�U�d�}�3E.��+��P*����]�G��$J���S������&NI#,�u��e��۷�������8mom�r@@����Q��ɓ��Z����I�{o��=������W��~�z$�]��M�W\�����O�:���Nm=k<���z�>5P!72z��&ӿ'c�8LT����`�%F��W�֔�Q�:��{�(�.�j�n�W�6I�cr��B {�t������FL59�o���� ����Oʓ���� ���+<`4�[�9���s�x�����3шs�����9�Ū��{Uh̷>6X��aP��U����V��މ�}�^����֩�+�@V����c����+@w2��4{����Tg����	4��Y���X!�����sajk��7@� �[6�Y�P�^�k�}u\�X�3z�,Axt*��[�����d�k�{���u�lh�ù��Zv�`�3$�F�ЊZ46s9+p�kA��c�Y������� ���������'��|A���Ǿ�GA�5����1"�!O��纴�,��W�����-2'�R,��43��4�,���T��G#�^YNҞ�{9s),��	��T�əx�.��t���o�}>�������}{��y��C}�.Ax��oj@����۷wm�9_�җ��'N�W[g�O��g�����'����X�p��iٛ���AZ��G�?G&D�t����L6u���,ǚ��^悆�7��0����+1/�7@:1vF�$��v��Mߣ�-�p5^V z7�x�0�ۈ� J<g�@�������z	�Z����pt}���
�Cf݇1��xN:�K��B@_�g�G��(BY�s i�NY�Wz+���]4���J�й"!�t ֹ³b�� a��<�wjЊ!%kb��^�yau�X���G*���J%9�&�� c�w�����j2��Y�;���Ӓ�{C&���G'P�#[s�(-k��N�����\*ﵱ� r����R�<X����H��� ]-t����('�m/7��!6�QjR��>u��3=��q>04XeS����U���7����	�	�7���}>H�N:���@A�0�a`$�)g)�=�߇��|<�ٻw��?���׿��s���n|�_8��O�ƳO>����}�<}�����������1sgX� ƒ�#s�:D�u'Uk4O�
4bq�=��4�R��)�L'�!t +�gV�T��n��4��rE"0����U�B��u��g�>O��h���x,B<+�c=�w��5|�E/ �^W���5��|	
��;R@G�	��'�,G�.P���ke��I�@7@/�;��k�Q:���io�g������3�*+E�g��
{��s�� �`�Q�	)�������sm�C4�\�Ai�D���֪�vaL�qk�<���-�,X�"����`��t�0f��j}sR�%�.�&��d�E����zb�`T��CrJ�Gx���<o�~O��3������gX���9����=�ٻw�766>����/��E/�������oj=N����Ŭ�=�����~��~��tRN ��Q) ��G?w0�2�c�	�(P���$q�y	I��@�<hak��J�S�/Ć����0n^ʵ�Db�yl��*m�NP�X���@�Y(�e���3������8�Sh��VIP�ց-�Фg�u�[�B5�k�et�GNK���n��:��/ZN�so�Ryq:v2����J�������)�ȇq���{K�-���hPdk�b&�~v���l��F�*"H#�sIر@9�K)K��q��2қ.�z`�˄Q�d��I�Q�$��<�T�r�x����g��)y8�{v
�7ܥ�PO7��j�!Q���_�dQ�}���{q�zNq�~/���~�?��_]__��S����{߾������??��Iv�s�_���^0��������_����9o��r N��p�9,Cgbvhiɗ���;�����˭] ^��B �#�y&?��DE UZ�Q��|.����]]��?r�>XA(�\s� G=i��?���>W�*�s��yS�q	�qF�m9�Z~G���͢,�_E?��
���(� �6e!���"}b�����ʬإ��}j�*u�c9�!�Уp���ʨ$(�5o������
�I��9����X�1�=���ץܿU���8����q}j��H��6�c֧B�,�,5��C�6F]?Ј���(Ċv��J �>�XO͉�{9�J�p1܋%�Z^��LWPgR���x�3g��<p���/���_<y��]��փ���'O��������nx��)�^���'_}�=����.Y��˝6��
֚���VM;�&E�Z�)�U�)d�� �EZh�F$Ț�-��t:�tɸ]�Z)�Zz���ޒ�9ԄDW��8V�j���5t��'�������|�|eh��漓&/�4׫&�E�e��G�9@�Y%��xb�^-��Ԡ.�����X(-Sbw����VUZx����r*��E��%����5��X��+��]ֶ�����%o�y?2Ƅ1 F\1S"*1.��e�7�[� m|W��etY��GZ]�<�\�L{\*��Q�jyY���Oons��ZI0֤P�j���?%�*��g��26W )��;��V􌵵�օ^t��#G>��W����~�g6�;��&���;g ��o���;op�G�{�����?�.��eC�4���O�vp
'�!#�2$���v�d�Y�!�'�DK���rXfu�y�$i,(Hf�&X��b�zצ�;TIU��e���w��Z>���[ ��e�퀾�����oA��][�	e-�/j�Q�'^�tMZӲ��c��Q�NES����Eٶ* ti���L�f��D�@���5�z %�!�T����	��:v�|�4kIW�,&�ej4g��m"��hx�f5��i}�N�G�jʲ5��%lJ��5Y��dnG�;�֞�Wc�yv�+��EI��B�z/���t�!Q6ʓ�T��s\o�{[i�e<�����޹���4��h
�*G.{b�2�iGJ^J����(i�u&�%� ��k�����wsweK3�M=c�*YLV��d�U�~@ђ�Q�J�N�^�ZJ|����aFpG5�:�)�dH����`��.����>��O��/��t�{�9�?��?��ԩ��~������FkNDB�H��4�JG�"��`0��7��R  �MN<��c��>/[�)������T#�e�" +���<��[�[.��o��(d#.�Xy�Ah5\��<Jg���ڸ��{�?���ZԔ�ƨT;�zb-�"�cm���
�����@kFd��,�x@����1<6O��K�H�T�P���喥mz�1��e�8Z�E��������f	Eכ�� ���)e��'a�	S� eewR� FB�5�!�1��M2�
� �II�nxqMt�P�hd��(���{�N
�(���n���S����&����GXW���[S��:����Ö��'�B����|eS�i�	4��6LJϬ�24�A�����0���i+����������8ZߢPQ�<T�i�x������<V�_��D�	�̸Ξ�0�4L�Hk�G/���O8��������׫�v� ��������=���ؿ����tK�	��V��a���)W��	���yt��,�e�L#�x_��F�FK��O�@I�H�{�n�ee�;v�;1�����r�u�F��n�\�֕�R����Y-���E9�e.��| �g�۟J�׭5�a-/��;�,A�-d�E��T΂:�����O�����у��&���7��*@�l�B��!bR�e�#�
 v�����d�k��%�ʻ&y<����a	�QW@�~��r1w�&�]�t��/������g�\*�e����D�vHi�fT>#�}->?���m^n��Z�����ͤ|�2G��{.��c�$h���N����=�i�voA��������h߾����S���w��sЏ������g}��?����w���TYPr� ��=&�9�+�j�W�%�yY��"n_�v��r.�?ٴJ �3����:N�F1B���b�Ү`�	��HAر,�YE�M��5��_�,OfWl&��R�f·�Xc��N���f��� ]3ѱ�P����m���l�f���p��"��DEx��{�j�vZ��JX��K������Qן�<�y5�b���O]�b/�l+�l{on����B��r�W�Q z0׳�#��ͲP_�K �r}��x�J��^��sTG�Iγ�>�8���A���I����}_r��"{Q���p:=�.���.���xE��CKEt%����7�~��������������*�ۿ�S��w��g~��?���߫� qwȩk��"��6سv��Q��rW,�t��`� �K�]s�GkMECE�Ŷ���Y'���xc��u��;\��K�^���Ș�U^e����S�� ��k.DacM�T���L0�$�ቭ9 4���ڗs�yy2�Dƺ�P�`=�֍ZL,���hm5�����:��Q�m¸�N����J��r������������ry~Lmt�B&x�<d�s9@uᑛ!�1���U��*[��]��6w�����isٺ)�X��n�t�z��|���q-ٯ|}V�)����4:�$+�p#*�ۀ��T�W�3��8��C��{!�2��W<��8������Z�!��E�D�.��u�ر�����G~��=��k��@����'����i��Dk�Qw;�u�x�e\s��o)�3+���f���[�kY�O�g�톖������5%�m���9�/�R�<j�4��s��s/�S�-�ƌ�s!���EpF�9�v��q����u�fٺ�h���=pa($11O�t�h���}(=����<�%�jc�7��ym�n�yh*fM�����q.�ޛܣT��%�p�Fk�z��x;et~r[ �|���_M6��f~��,y���d�s�K����5�)�>(��R���q�ֆ�\y��s�y�}��~���8��K�@��߿�̙ٕ?�}���|-��D-�
$��d����LZsF]V���Km_r&/˔B��S)P�6�(�#X�Q]�,�#aԁ$���zۣ#@,���3��Y��U¡wyKRQӓ���-��ǭ��,��O	`�"?����=�eY�g
�f�����@�x?�ߠX�2Ьq�=e/9�+X�Y�n�cM�*��2�-�j�wl�[�#_��:�e����v`��/f��Ҡ�ը)X9��̍V\W�*��
aZ�B�J����\C	�D:�|�����:����>N4��;�Ω�C�����:�����Nֹ>CY�Ç�y���u�y?�ۿ����m�w�s��B߻���>�s�������tl(�� �pXߢ�Ǥ����ܵ��z�q�D�ǆEĖ�o�J�:�-�����^F �.VV��	Ɲ�|��m���.$���v�]�<v��;H	dW ]{�����[5�-�l�tY���+���֪UXFq�d��Rf�ii�w���]е�(���d����֧� �N֡m�� =*�exϪ�+��E�������e{��D��賖�L�i7=̭�� �@_N�o�OV�(6�B �Wᝠ{~?��#�]�5�N��~L'z$+\�Ї��C�|�U�q�����[�����m���u:%ŝ�����c?p���	q,ZX;Bf�2�����qcE��:�1��@�L�E'�U�o�]Xg҆E,�(�n���m����8��{ۜj�
ժ���5E�]Ȋ{�2q�ѱ��y�3�5�ϧ��n�n\U��xĥ�zm�]��
|�:Cc�́�%�]����)=V���kJ0.��6@��X�@��[mE�8^�?]��]�N��s�\)�p՞.��à�=��������ݪ�jW9v�D��vtez�	}����S26}?z�s���G��_��_��.{��ל����*���]�A\[r>���/Q�    IDAT[U&A�6J�9}��	aƲ%��zC��A���LcI�A햬ZC� mև��d�����b��$q��A6��R��h��]H<O do��m��7��g�uɟ��Z�$J}tK,yޑ�b"fZ��WA��'�%����V�����oy�{)ī�[�߱�zX��+4��{��8b�&�<k���*]*�)'�"�G����܅�ē�U��beV�4WZ����^�pByͪ��y�j�q���e����L5����`�� N��K��a�Yi2@���C�b���9@I˯�Л�s�Su����H3r�?��g?�����' }	������Y,��$��$����H�qk^X�p�jc���C��^�%��������e2,\�������ַ�܅P�&s��b�e2K�� DmXF�8uՄ����NéWv���f9���=B�;0h��m}/����Ѫ�5c�晽\��bv~��x�Ϭ���_Y�5����o촖__����]�
S�.���n���%\���O(��ϼ� x�s��
����y=������/��Q!\�f]�����K�l��d��z�Qt�)��fN��7���K�C�c_���o�-���6�W[AGP�{Nb�h :ٓ\.����p�����_=r�_��_���u��v�.�Ю�e�().�}W����7<�����M���]Uh͇FwyF��|i=�r��V[���Aa�(�cd�etmԥ�\�*��+VӪ��{�U��j�c�mB�����*&�]�7���1;r��D��,� (eJ��J��/�&�k�ܣ�^ ��k��/���y9ٛ�Ŵ�㈥�B]y��5)?�3�=�@��he��P�����D�[�8U8�r�ȶ��`7���2U��x���e��o��䉆�G�C����z=�;�Y9���Z��{}�u�4�s������Ӊ�r rx�<,���8�$IX��qً]+]ʥ#��DG���?������G��������s)�w�γz� �����?�<���l-�i7L�Vf �s'� D*MEІ�(�N�9p�7D-]W��u�M�H���x�ν`	3����L��E�WJY�-e���M�e�X��� �T����PTv�ʾ/�h�u��/b��U���o]��ܖz�F�r�{k�`>�eS�Kh�1�
D ��D���쀎�6X4�4ω���RS���E�*�Ř8e��-�ӈ�k�ﳆ$�Sx�ҥ��=h�h��cv���^\��Pm:۪��9��~������,?�#QR���s	�Ѐ[�u�5�����������
�GѳX�B�U�}��|�n/�-���Yf8���J>1@�EX��4x�/�rW��>�! }48���?��G�>���������1��F��ᑏϭ�kk����?�At�A��5i�?����c'1p=�x�-�G��ܥY2��:�YM@��T�� %����x�Y%��XT�CkͰbe�x�l���_I�˼����rхi' ���*�� EQ	ie풳A`q�!����!�n��(��Z�����,l]a�e(��-W��rtuVM�e$Jѩ=�E�����I�P�I�L4q4l%�~���4V���w��Ԧ �)0u��|�Ј���|�FfeJ��K�C�{1»�㽆�!�+��������CWh��Z�L�,�t�ᳶ�o��rA	T�
.kZ�ҕ�.�j�nf�^h�~��h�}^BR�E*���\��+m,��*u^��� �KOPŁ����Z����ǵ"E�z�w�K�g�1�Pw��]G =H��EZ���5���ѧ>����~��v�#��s�?�lln.��?��O�����_ﱌ[訩�cU}�5&��p�f}��o��}h����!�:FlMy4�b +��Dq��$� � �j�Z��.`U~�ó�\V��W�ٺ��k7g�G�!�z�5���" *�R0��e�P�Zh��=y��H�㽍�#"�[(j]�r�{��"PY�`�
W�	"����@h�<1b�v�$�&��k����� �R������K�����M=���XQVU�h������@.<X-�PԲY��M�"U���Voɛ�ə" �\�X�˟�q?_� ��{�de��P�`8�Is�s��n�����=�{Į�Csf��^V�~��>�b�-�9� 0�g6E;|uQB��+T�drC�a�d@��Gt0K^�²����E��X��k_��/��W~����c◳����c�>�q��K����MǏ�����_i�䊷�4"��Y��1��f-',�/�*p���=b6��E�jf&>�iA�2�����
����Q���0���YȈ̲���Ѽ�A-����+6i�'�H�nQ8��>d���Z�5D��e��´)}�%15�h���w����x�S<,f�'�@kA'����\Q��*�s�4����?��L���T�Lxl�.B3S��I�_�1�0!���U>��[�f��8B�/E2)�8���Jt+��PY�C��[�aA���h]�M�����T8�a�j�fX�@	vG�r����������a����\Q*8�\%r�χ�g���sƖ��ʣ�c踟�!@�IP��bh:5����Pi[�� �h��4:�gQ,��蒈��}�W���{�^����z�}�#�����t�9��v��x<x�;��#�?���oD�;m�����v�������%��f��Έ��e��e|j�Nhqֺ}b�T����t� +OM6����"�A(�l��U�'����X ���$�FXB�_�d�m3)s�~f�`�� ~�7���$hD��xM�Y�:+4�����E �B��@Y੅d�"^�y�7��Y"�gK������C4I�	?PFBNn�#.,ˠ�]���/�A-�T�S@��W��a��_BА�g"s7�F#l����$�>�R�ݭ*�FT����Yu4r���|3�AF˦L��Q�m<o����.��dc�g])��y_X��4�r �h������
1>�R��+���3G@/H.kR��_Z��]�Q�V@7Ê���%����Z�;������>����#k�����QM�7��}�_��K/���>����O�b������x��oz�M�O�����	��Qyh���t�y!��:ز�i-���X�X��b�-τv\�q�@l����, '����,FY�@.� SZF\�����j�� k�-Ɋߥ2���T��~����G<T�@iOa��=0���`� ��,�lQ�X)lT��J��=SP ࣀ^(�2~���~�k���6Թ� dBۀAÿ���%+��ŗW�[�Iq�J-��k��̡��jg�D)m�d�W� BH��A��g�+B	�}�gEuFڦ�&@O�������x)�fh9F�t�)+�Ɔu���&no�$錍I!oa�:��ܝ�dE@N@-�t�=Q}��G�7�8���p��r�2>���2D� ��b��+-tyF���
�yZ_���_�]z�%���~�3�f/}�9�Ţ��~p��z��������mK0��.���N.��F�{W]��Ẹrd�յZ��ukX�&3�0�s3�I��p�Q�mQb����$�����;�҃�]����'�ɓ���"5%ؔ�	�����p��(�3�� 
B���ާ7�k0/�JdT�b�u�]9R�PC'
�\��NY��,�ͦ���[� w��p`xE��BOֲ�6��+��l���Vd��ʫ\��rs���kK;�����L?�����,�SV��i�� ��鿔-��A@�d�V�Zg��5�'s�U3�q�`�
9.Y���$7�X�\o0��B��{��k]��M+\���.l��k%�gh�<3��سI����ͰZ
���N#0�}&�O�.�v :=�����N�[[}�[��[>x��.�����O���޲��v�`��K���u��M�N�f�5&^�3b=)�v�,��5�Q�RnsψD��Y{��(8��=.��]�h��L�x�����hYﲨ{�����:�T�|b.6�\�|]kgp�Zb�In�Bn0n�L��	f��ڤUmR�!���%��'�G���⧆�t����wګ+�a?B%��D��L.�u���� U��sL�A1�DB%�>�Jp�����V}n �0Ht[dJ�ѥZh@�����Cax]��D�� $�DΈ`O����	��Z���Zv����8�l��e��k��sE�r�gcC�9쵲&''������֖�ǆ�$���MI��U#���a����� ��͸+]���#N]H��<���}�/����?�7~�'~�ϻP�n^�E��������G������'On��b����H��0�7��2q�	Х���Z�ŗ�>3���V��G:
K��,�V��2�3��ZW�n�����KK�i����y��L[)���  Ȋ����M�f����!�J�N-\��K����2=�O�lV���$d#
��na�����\��弍�3̒e�pP��븩��|�+ժ��W�ɕt�f�Wi���
�V��`���:Dn	b����H�~��r���]���6x��!2�+�����ȵl��*�HN,Tm����$2�A�a�P1�}��P*f�Er|� n���X�	�5����0~�p30tÐ�)���v\g�p���*b�톗��� ��2��-:)��u]h����g7Kkkk����/�ɫ�u�o��{��Wgxgy�N��,_�;�E@?u�$:�1�C�	K�ؤƺ8�j���b5���ؔ��s@�g��iD�`uʝJ�(="&@.�y��1�m��6ϲ���P���c��ot�$*�3�B��P<��hJ���h'�Y� ��Q��E8x��Ie�	y���l�����X�j���(@',�X�z��GzԊ���lV��f��l�R�eJQ�U����Z&A�׋bj�B��y�L!l�g��-Js�71��\W�9JW���3K9SE+��^�������M�X]x+hc����rz2�B�D6Uz��c�h���O2��cҦ�+���#���/fp�H���(�"R@W����n$�e0jx���B�A�vOB��NUN/�ʉ�_�uɬWr�g��~ӌU2Խ`��rXs�@_�Ik��$�9g�+��˺İ-7�Q�|�6��˾�e?���^���{�����j��u�����?���Mth�%��l�YY@n�@���>2s�p/YR���Vb�p�y�Ԃ�z\XUЯJf�@# "�e���

��⚨��Ϩ����Tl����PT�Q�g�W�ʾD��TŅ�e���LU�Ӭ�W[x]L��nU8���ⶨ��"��_X;$�q˅s����Vt���������C4!"�gp�#��7���XW@~��\FcXO`���q��vޡJ��}'@�҅�2e@�$���ʱ1��yL �r���� �e� -^}��r THʖ�a86U��JD�_�ZA�-�Ԭl�M�-^��no�GH��~���l�B��-ky�{8�HW�Y�LD4p��[ނ*Xt���S�(MB��4��-���)��M[��1t��'"
ﰗ8��|��^������{��M_:۵?���@�ԧ>5��W9��w��Ɠ'7����$�򰄃���r�CG��(�v�ٳVnMwwcS,)$w��Vv���w�j�tUh�d�KY���
�,*�U�x�R3�!]���o�"�BgQ�V8&؈qb�bƲhq�+"��]�<P�E�f���$J�/֗ ���%k�5��
'����}`�A^�2*UH����%��it�� L���ř�y�c� <!XG��
d�+p�5U�+J,��\竳�)���\��Vo��!�R��<������v����� :[l�6�S�'8Ɇ�nz�=q�žozuĻ�Շ����c���Lܗ!E#͆��m�
���~�P'� � ��8�ey�zh��%��s�wE en�Rv7��-u��ס��+]IY�P�ҵ�W��e����6$~��|`t��e�����o8q��[bc�x���\ā�#c��.wa��O�( <i3� ����T��
!f��Ʌ��1����o|�fG�c��~�	SѩT��g�� �Ƶ#�W�"c�0!�i�"܂�.Xi�Ǚ� =ľ�^c^�Z��tԴb\��|}�Eb^P�j|!
R0׭�(8z�J��ĨV���hy��t�F��|{��ͽ/�\t��
���q	�ɥP���PR�$Ty7ꔕ��eK����{(�eݬ���Ž ����-tT���P��,z	�xՔK��A�r�l��T�*W�\�	�u=�˴V�k�g`P���'h�	U��%���L&C�I�UT�caH}�P� ���f��̴���~����c���h�j,ӗ�g�����=��E�3:�P/���#<���/�����E/��[o}����8��3��qD��~���_;�#��ַ}��xS�F�I?1������h��M���=J���5����ŵQ�@a�W�f�W͖5�V�l4M���F��jeD"֗;fmkA~���1�u��y�, ��;X�j�0c�>���p)/3yp����'X",+N���]g�����Hqx8��p�5&q��	�ӵT9��z���>E/mAA9\�+�8%�S5x���p�J~JK�X�O��DRV5w�������5t��jHb��_��$b��0����@��<k���;��RTh�0d��d���:�5�]in�M�c��l�
 :��v"��iS��0�*�B�M�F����ܸO��ݖw��/Ǽ���D���YL�����K���[�i'QHG��\D.�X*���i4<~#@���#��r��J�p� }>�R�/_���������;�r����/?� ���v�7wt��%�ig��@����L�-`�i��v&�\��f�r�m�3,^��,�<0�%��r>��8hcs���WT`� s�BR�TC6�^��'0F}�+i�nvHa2 �������rC#�2ĿWE����*�E,�T~dX͆E���_�*�B�����1_u#*뢠��GB�B���ͤ$V8!p�ګuFp�{�h�Ii֦ ��n����2Ù�� ϙ�^���H�ixr�:׺d掾���giR��]���V>�dF�W��Q�TX�Џ):�����"Bt��`(���
n�wA�����D�yMi��Bsn���Q��i��'�T!�+d�kb�X����`�X�/�T�j,c�h�=]Z� ��ӽ���Ϧi8��u���~�K_��o{��~,�<�{�Jͳy���C.�C�.>r�M7���G��f*Ms�:�F��Ͳfk5��	��]��0�N�M���K���e�3�1C��l1b�I<�@�OE�p֫38�w���t��9Y��a=�	ul�iI
������Al��R�[������,?~�]ݚH�	3���H���~[$������ec�J<N�E�%D�,��k47�J8j����Q��c������9K�W%Bc��l^�d�,y/[:f.Q2ue5V�<b^�)Y(�����
�Ӊ��5k�1��8YW�*H�2�Q_&�n ��
@<9�עE��o�w-��j�F1Z�f�A3�}>��V�<V�ʠ��u��5��a.{F���V��q��^q�*Z�K��K��L�U� ��@
��^��6W=�{�+��� @��1�N�ń�'թRJ�2��]U6��n޾z�������]c��%�*t�
Хl��i��W\w�/}�\�|��v�sБ��c�n��|�zj,K��P�У+�l,â1d���̥�띷5�T"�����`�c����,�F�8��fͶ�KC-װ���� ���u*�Z��ɭ{$"�4�+X��f������I�"|�9!D:)���a@�1H�I{X��� aHׁ	�D�!�X��~���4	�Gw�3���a=qg0}u<F��Uq���9��    IDAT�Bb��v�	.�\�b�L�Ĥ�w�,���'C�4�9��3���H�)�p\�A�7PR��%���/��y�lJn�U&gI+�����Z/b���S@'h) ��G��.v=���)��^C�"��0��)'b!��BD�Y-�\Ҡip�f�DQ�����JkP��]�l���s�F�ʋ6Q)�r� �V�La���,ƶ
:��`R�}���F�V:<`�%Һ�D.�g�7�Ni��zi��:�e�����^��X�-���W��N�ےi����
�E!w�{�����V%����W\���e���������j�w��s�Q���7� 7��� �:�ɩ��1QH��qN0z��v�&��]s��a�FL�sj�#`�5�20�I���|�\��8~G����\�b%�}�_c�1i��(��M�Q��[(AY��n���4�+ʉ>ń��Z��dF�"uH@���[�ǈ�]��z�ۿ�Z{
/B�� �e�驮BO��0���:�����+�DJ����`���kP]��:���wZV����f��'��@,>U�x|�H���{�B�9
殴���%a���p��t�#�^�'~���4���5�V�E�2զ@�H��''sy�&E���}.�ę��(,|�k�'HʪYۙ!��q�����T���H��>�8VW�bj�S��N�S7]�-F���Wu|:-&g�bv:�&����J��$�ӌ]Y�`�/D�9�c��z���6o��]���f��#�h�
����xŷ��_���������w	>.?�S��ҡ�o��M���,qQK]p-W%ͽRh�w����˼�l˔��
��`��`�ŢVH�y�1 E���%y��v|���pܧM=��� �%3f�� ���f�� ���hE�q��qPMu���"�����z3�	�[չ�l��,@�ʄ>�bԳ2D�ERÞ��wI�{<�-S�+���F]�������t�u//�ҕ�Z�kA���ak�Zw�ڌ��7J@�i�l�髀�GF�KKw%ꮣ���(dy���a8Xi�����y�3t��g��B�����
��#��X���¼#)a~��PP�9_F��%A�\��� ��@L�0V�7�˼VJ{z���y/-l�����5"ʥ�{C�<��v�]�L�z���/��邒Ȅ�H�@���x+���4?�N>�����L��8Ҕ�dRʔ��U�З{�}ĸ۬x�Z�n��BN���TL�����/����O��կ>�rw��s
����haK��kVz�jQ(-s�4��u@��߼^�,Ӭ7J��z�9?��?/�ٳW~��y��I �����ڈ�7�(�.4��d�_0�{�[hC��I��6���4q#j5��Ld��e���\�p%�V�~sɆ�LŚӬ`v[��p8b~����G�����{B\M��*6�.���̅��`dP��'a��D,DL�~g��a���>73�k�q�c֨)��]�d��h`���M�X"��t,[�`wK��'MŻ��ʼ@܈Ic�!�-k�;b������gVx�B�$���D�><4�g����x�|��`�-���s�0@k#�eM��'FoӒ6�8t�Wx��;4�TI��� s���s���H�~{J��m�K4��a0{%�e���;r�:K�9��%�H��ip��"���N$LSo�h:����l����Ї�����!�c@ף�; z��;�x��z��D@��{�����^���'��=���.���ǝS�N��o�M'O�2�{�e,���Bw��i/t0��"?��)���i�[K�������L���im�ƬAD?�Q)���)��Dܝ�#K�
��
!K
$�?H3v7�ZY����*�Z��"?Vw�Y�_S7.��D%�q��xs�GZ�� �$��
���z�����7Z�6�>չY��O�Tpv��F��g�oXGN~����e��W(�C|߄;�ܯ��Z��k��R��R^�@��!��x�����Y!����!�Ax��|O�������I� :R�Р�,8ƜU(	y�DA�%k��,n��J�E�Li�JK@QE<:m3�s˔��\)T]۵p8����5T9N�4����,�x�t�5#L�E���~��P�HP8��2��	�)�}��H{F�ԟ�L~��i��H��4XP,}�Ql���#L�%�/�.Wb[f�t��#�K:��;��=�_�7��(˽�O_z��{�������3�������Q��]vvw�x�O�zJi��o��w�<)�G����v
���V�[@��jQ�pvm�B�<�o�����q��4L�޺f�[9��`�qִ
��CB���W/�����>�BY�IЄU.$N��$�ng+5|��qB�!�Z="2u|\�x�&d�Y8�w j �G(#���&*53TI躴	BSd��ka��s�*�Y�O���*KX��_d�{M�s���n�M��h�u[�q���i	���=X����yw4.�r��	��v�dH$�1�0J�E�Ȅ��:���F��\	8e��߾�~Y}��kɜ<x�N�5/
�'��g��@�+_m���W�ݫ��{�
= ��4�_��Z��gi0?��� Y����L��i����¦�x1d�o�*��Uk���$��>��a�x�Ƀ�r��#=������߼��׾�]����]�uj�w��sЏ;��Ӟ�v�;�w�������%�#G��36x�F7��J��r@�mb@�I���ix��4L�� �����M�Dm��d��3Q�+�K=�	���
���뫀��y)f�g"S�ba-;��O�� *-�\�$�,I7?L"s�c�P�l�R<S�Bcx�v���B\,QArK�W�cC4�3�e߃�X�-�б,b��7�I УJ���k�O��ʐ�M��`A�M˕��t@f(f�v[���K�U�X<'=Cx�~��cKg��EM� ]��h�zƤt���Wd��D2'-ڜ�F(�2I����R�o
_�4��|I�/���<����K3����������t�u��S��`1Nk��4�m�S��mZ�I���ԟ��`N�q�h.��%:�k�`Χ;�f��ϑ �f�ûQ ��r f�!�|4�����=��������O�6`�z�9����v[�Moy�͓�����3�9+�k a���]��M�h�©�M�R��J��?+^F.�A�������4<|U��q�P�sᗉ�$��_ex�^��#�v��m�-d����Ez�Xe�L\� m�֕�<��`�G9-��!��5� ���� �W-�`,�+�,-+�r�h�~/�<f�� ђ܊5B 5�1�J��JIᎍ�]&��<���BO=D7��*6�5�~��^	Р��@D��p�2� ���
<Ux��bE��k�7C��*TABO�.BY�_�{�C���~P&
Z,���R:ߞ��1��oC��aZ΁�G%��i�L�p��N?|G�o?�zӓ\�F<��*/��6�RV$dB)�Ѯr����<����uz�j"	�
�SX��$� �#
�o�)M���y��^s��o��W��g���x}߅v�w��s���+o^,��9sfm>��#.G�c/waHw�.'(��ǌ�,J���;���0D���k�ߗf��ᡫ�dx8��[�����{=�-�E3-@,,JJ�wZ[sZ���m6W�#��PAG�/(#�ɦT�3�`Ff.�䔵��;G7'��z] ���xJ��D�㰊�C�2iY>S�3X��j�fX��6شLSQ�C���ar/�BCi�2<"��E��@-d�[StmmJ�m/,�@*rDa@cy\��Ѳ8�o������"�[ֿ���G�E�� ��C �#~�����:����c��s8�(C �~����(��<?�C�n����
��I[�i:e�K�p���-���Oi�h�����ǿ��[��d3��Ě�{��N}��N�:�NP٦򙮩��g�|�'����?��`ا�N �__}ճ_��?��?���Ζ���sЏ>����Y��}�D�$�86�$����Wg��U�嬢H��6��E`�ͦ�'���4�O������4J��F�1��à��YFVm�3����̳#�%�����1�2��h�	�r}uD��2��VRKw5�{�1����7�z�p�
�.\��XQQ]tܑhy���--�k��6���aL��*���gG�8+�U.��i+-��r�w��O��O)�5x��9\͕�M<��L����Ie�+��=�sm�[%S]��ΐ��V��1��'e?�r�"�d\}�:�E?b��&z�~�;����#��}�K�3����8�4��bW)����w�����0KHF$�Щڈ,���1�?��N�վ�����p�UW���~�_����a�}�;R��<����f��sY�Zx���p˸p�g>wA$Q�i'%Q�"���Y(��6����+�tp0M�r@�杽�vz�E��%`$w[wx ,���/),�.��������v�[fx7��;Y�[#� *�d-�PyG	X+@�AA@�fy&���^�wa�.[��25V�|��{V*>��1�u';�r�{j�,<Q��� ����=-�G�x�kK��e���[��,qv�H�h�3�K�_���~�3�����i�Ϧޙ{�`v�,{�ŧ��jNֲ8��l:la�,�5p�G0�k)oos�	�mD�D؁�	u�I��_~�e������|�ëw���b�]�v��O��,��t�� ��%X�х���]�5� �ق�H�
�:P�Da����C$�5��Lb�f@/���g'vg�wN��3�w����X�z������}��Kw�bm#�4�L�>g�sc!]Ji���o}���{E�� q�����HF����V}�])��i��6r�FB[:\k��_�c��~�]/<W1AQ�2�3�G}~�^V�!�V�N�|L��*�NO$@���$����}�I�3����tZ������D
e��U��0(T�H%�#�R*丹6=��ޤ�!|v�,�d>�.���O}�S_����_^w�u�H�w�g���t\�/#@_,�͓ɤ�"Ü�V���h��~�� �!���V�O�{@g�9������Ч�Ci���h���G���;a��%�
zx��j��ڕ�����}��Fdi���F��n�����'�ͥ=2� ����y���� =*��۠��2�9��Y���*>��vP�و��,Q��<�=�Z�]�$�2�%�|��a9�O��՟+�ZH���<rZ,G �^��Z�π3��� �6�5���i��Ϧ���Щ�g�Tdg8�4�K�E���a�Zgލ�ޖ8gim:��^!H��:r�,��q����K.y�G?��|�_<y�|V��Dޜ�v�� ��r�B���f���q�6;ZX�.��ĕ$��I��%��b@ߐ��)ա��줸�5�`�w�݄�-�e-���er9���,ږ��P�mn�d��NBmE�`���}lHU:�sjrB-��6$���|޵�n}��4���FH��.Z%�U.�Ӯ��ݙ�x��2������Hr��L�<7�t�/����L����z�`@��1	C��yJk�i�I��,�9�~J��S�K����))	Y׳�_� ]x{&	�C�N�t��f��S=#������ף֯��b���]z��މSJ] �6)hh]67tw���e2+��y�K	�N��y���,��i��4b@W=+�i�}].X�]׳�u`Hѕw(4����� :��������ٴq\��K ���H�㲄+��-�K�V�h�vW>+��˃�����n>{�v/�zsX��r=[r۔a�7]u�2��*�Z��^������?@�,8t�Ӟ��Z:9Oi}H�~"M���Щl�����yY�6j������YU��eu����N�)����Zm��O�iN��9��O��x2�O���/z����ƿz��_����j����x�|>7���[iԪ��3@'"a��p���<�^� tq���ߪy/�))np��e�+�:Ȫ�h��iw���|uW����r���N��ɵ��ca钴5[鰩�4��k�ʬ�.�RS[�����k�q��^}NW�YVR՜aTv��k�r�)bj]rXA�h]�kU�B�`c��(;�U�[u��/��:���Ĺa�<%u�A���I!Z��Z:���UJ��Ki�����ԧ�2��5�sT	Лm��9vQJk�A��d�[���x��n i��g��N'�ͦ���l����U���u�<�[>�k���c|����\���k��E� ���b%
<P�3@G�/m/NM�g�����Չc�=r�/aޝZ�1V?��1m �{�tz��wb��5�eZke͚x\l�ec�1Z]���܋���ܝ�9 ���VJv�ŉ�ն�;x�壬''���m�3�Ń�n��unQAQ�n
EC,�����]P,�lk�AUM:I�R馜tbJu�[�x�/~�����Ɖ��/V9{��| ��[Q]?mp��f�=�`@4M��*,y�I며=J���
���%��_�>���N�����Y�^g-�큔<�ҐZoO�[���������x�]�d7��Db�������O����b~�x<�K:m^Y�~6`�� tm^��À�m�n	�N�L��1���lt8M���&,ճ���La��V�eu�e�ﱮ�+�2�� -L����Y�/>=w���gs����x�{9f5�$�@�	��r��QE@��a�:���HZAt�ћ}��j��ҽff��w���| mK����P�t'�\�Y���ܲ|V��9�	�C�7�H2D?
�Z��,ODl�L�+��K���4�Q�^�E�=Z�1�3F�{O�p���)�,��I�,βg��&}�}1~�]���A�U�'��x�-tjZ��WI�:>P����N��0	й��s)Y�{i:���N��_������ =-7m����΀�i���{D��ȓ�̡�I�G��������ѧ,��it��i6:ĭ_9_`ǒ@�-=�ЅpTPP���/��g
�����;�7�W��d��질u��w,���=�S�I�{�������M1��J��"�'wA��󤺮s,�!2`�z��{����˔ҥkۥD"�gk�VlsU���obS���&`i�����c�2�N����������<����������ڷ��j�o�LqrI���a+i΀���L���gHi��fH���ҁ,z$+�< �f_NL�RM��C�6@�n�t����Y�So+�:��i��OOg۟���}З�@���S��!�����N?E���:�t�M%rQМ��yD��W����6���8ĭ�K3r��Mk��)���!PsAZM�]���M$:��˜�Q�w���L��&����Y���'6�2��fU �^/�GeF�狝��aE8
Rެ��^1�DI�%��h�p�GW)K+Pτ��0�#Z��5l��S��b������Z�bM�ĲJ���4��%C�����V��=��Z(�~G+_��L*z����;���9D��A��k��|'�NN�E�T�cU78�~*m�RZ�y0��)�%���C!h�l�5��~�w��`Y]W�d���@-����q`5����W@��i2��N�?��/^����7;%�ݸ����/ڭg<�)W�}>��4����f��A!���)pY�o.'�)���.�5tnl�/:%ŭ�: z�\�da�\��.�{�8�c�rG��e_X��z|�Our�V]��Ҽ���>�!.�|���%+Qseן�n�,uW�0NxB,��+`�X���hO��V����� -IO2/JP�Џ*�ܿC��sͯZ@f��k�0�z�?K]��hU�+��@����]��wI��Yӽ�V��@߅�Y�nb�){��Zơx����z���G~z�6�՞U׊���-��:�3�F����a�HAU8�=\���+�:�E��&b�TG�D����l;(A��	е#=�Ы�*`N��6����h��_�q�| ��~�"    IDATg,k�U�� :g�se��g8�o�����R����A��N�$@�j	�����t�lrz<�zл�
�9�g�=-�7M������o�^��Z��Ev�y���.�~��3�)�e�����,-��Ro�Ѵq�J>mm{����w�E@�oY^'�6�$���l� X�$��t����DC�K#��k\4V�2��XB�F%$ ��[XP��� �蚖��V�c^?��Z�|Ȉ|8	=G��yA�������p�	ݥqC�I.������E"�ǖe���+�������l��0�����j>c!I--y<���C�Lb��,���{J��ʀ�ˤ�g8�ր~Q�U���2"}�]��U�&��ji0�{�/[�^4lk��6�c=H��H�!�Xi<�4�9[���I=�<G���B���T[)cb�J���(��K��1B�P ̀վ���Ɖ9b,Lg� ^�C��K�k#9���z�rI�S�0w~F_ʳ�f �
�L+���b��ș�i�K�/ߝ~�����������$�bϛD����U��v��������eY@��f�k�nV:4&��t�;=�O>7�^����z`W@�l6=@:�(?-k  ����i�r�X��c�M_��+�Yt�Z� t�b�k����'����4�����M���UI�F����`�dħ
�dh�X��clK$�-kn���������_$�4�/��Z��I�U�c"w��%�Xy"�����&�/?	<G�ǢD��ay&�VlEXhkjRt����"��� ̱��[ZF-u�	pDk>
�Pn��`�2 �Q�*J��Ɯ{9O�D`,�:��Z\d�����"�Sw.��%y�&��EJ�a/G�,zq���[6�����^���⾘bLs4�m���\oc�)���Q	�~Hrv4���) �����Jt���*(��|�I�|���U'y@����z��G�a�Os���?W~έ�Y��A��Lo��O�&MU }ră:��u.J#��/.h1��܀��yS�8�6}���ӭo�������0M�Ӧ��<W��=�HV��<�1a��2����H�+"��'����$�QR�b1;5�O�����	@_������������y��l��3B������{l�X3J�br+3����0��z�����xH�[�s~:���ӳ��i��P�H�@�G�)�qO`v�"36�B7��-���&ա�<�?	��YG�Np�,$��H.C[/��5i�p���VD�	H��"���{���~����Q� >�C-c�V.$MA�`tqaW��Fd11��el���F����5~rC��k#q���?�~#�k/ֹ�$Y�躐�+em	���*�%nn���G O��P*�(%�'سK\&�,nVY�qg k*7p��We��X�}��U͎̟�ZT�t��.�X�oo�w���������(MP�+�ړ�k��S|)bG�ޜ�6��jx�&�V�+��X/5B��Tv����P!<T e�������w����}If�2���N{s�|��_J�^��t��_b���]-�u�pary��?ՐЉ֌��B7_6ׁ�ge_��	�l��~� t/g�:��bzR�uO zG�~�S�z�<�o��	�q�Z�E�<��kk�Zo���
�$�	(C��{����L�|�sӛ������.IS�Ι�H8����0n��S�,]��[�1��ږ��>���/$g(��^X*��)�ߘ>3 ���d �'\�-���f����|F���,�쒦�&�E�����< �y8t�q�ˊ�$�ѿ%Q��u�,a��5�!��$���GYOqz�V[��O�kH�!�|H� ���7j���7I�CA^�W���GC�L�{�7 N�xW&[ߒ�ċ+T@�@ÕK5+����m�����z�)!��e\�Aм��ٌ��QX+�y/�j��u3�b������ c�N��yG����B"ύ �<��Ad����A�Pv��w�y{z�ۮOw��7�| ��b�x�=)qL˓C˹,#�(�k���)/!�3�P�{(~nY���`CL ���4x��ޑ��r�Uo]��7l�Ǉj��D@V�ơ�ؕ�g*M�SU��=�� 
�e�/����`��k�;�uk���K�t�6*u�M�⇵�Z=߮c�Zxe���)@B�Ĥ��r�Rg�J �q�L�S��E�VC>��'a�QH�)h�{	��ThJ�Dzxq �Z�q|%֗�q$�����=fmNs)d/|͉~�>��*Ⲑ$7 4,tq��ל���'�*�	���%�Q���GA��& �6lxA򝂌��5o'>V?:r��˚c�����k�m K02>G+�[����ݬ������Ae�h��DA���
��屉��m�!���-2ıy&��~�fdP�hx�b���%.3;:X���3�~	�o��m�ۿ��Nt-����j^MM��N5K]x�yC����G�� ]CW걄un�eT!d��jlf����)���' }5�����[[[�ذh����t�����Iq���mtNRW0��U7�)��N�^{m���[�E]�&�q��TP�8
{ ����2�Z2�<R!k���E��B[a4�]�w9]a�	N ��V2Rd8|��.s��n���3a����d�?K]'=٩9Xp����!J�窛+��x�Dxj�,�%In�T��s�A/MfS��㽔�E�w�vh_ɒ �����A(q~ƀ����v6�{��f�5eY��]��Cf��gȈn|Q<�X���F\�x~P`�#`����ѵV�?�7���5,���`�ĔN�6�o�ZMG���<a|Z#�`T���jת5��(�eg�e�&�M���|���l�a����1��=EvĔd�����>��i%�t-��+(��z���;ӭ7�=�u��i>��))�*hqv��>W��E�5����#\�,�塡&�I���l���,<'˃�&8L�Gi��4�}���_�.9v��v�h�ޱ�Or@?sh6��2�9���Bo�r�+��Ft?�6	�L[��J/ @���t�E��D �C�fȟ�5Ě$S�����I�  *(rL~Xe#	o��iV Hy�,e{N͔���±$wq�B�/c�l>8s�����/[��і�HG��V�X�)-�z��(�����M�gǓ	��Jh8�~m����>Ӕp8D�r w��]��Y��2�1>��/�`��'�w�1��]u�HZ�K ��z�+�i�<ؙ�$�7��(Z�wuU�_CIYkn���t�ċX?+'����|<Z��<���ʀ�Y�
d�j�U��Fx�9S�ri�xʀ�-��u>�p0�+�
��R)4BM�߮���$O#L��s�����S.�ӯ g�^��C��{)�}��nLw�~� �u� @_�(�}���*09k@g��,,kT��#J2�9�<�}����g������:����W��N�>'�;Y��� �֬� ������ƛ�Q��20�#�������$����&���w2�o��.B5��2(6�<f�(n@�6T	�5�9��� �����]֨����Ƽ�L�q���,QF��[�n���w���sP���4moo��t�����%W�y{2N[�q"۠?r�2}�1=2�)�!�o���u��6^#��3 ov#��.S̯�`@���я/�=�f���g�����۞�/��k�{Yh�gt"���>H,Q�J�ZXc�/� "�9��5�N��Q���yDH�������Z�cU�&C���4��*�l�h&�f��}�]�nJw�q{��E���Bg�NY�ؑ:�Y%��T��Y�:C~+ =�Y)�q�@������?��ox���w�^ցw�}��a��omo�ϩ5��+�V�E�&��@#�C`��(��X�<K��w�y�y/xA��]?d�N���@/K� sL��7Y�2;ȋ�wq��ǚ��ݒ���Ţ�M�`#Ʈ��_� �Hf�CMAhe9��'{|,s
�Fb��Zdmu�{"#@��-R�S׬��t3��k�-��,�8q"mnn�5�^_Kkk�i}4J��$���J[�IZ[_O{8�y�̙t��i������}��������p���kkk����3|s�G�X%�5~�v;��O�eN��IW�'��b>��zU���uTr�fFh$��V�cc�+�m��D�".�T�BA�a^�Z�Zi��n��G��$����g�h�j�? �v�	����"�V�F��W� ꭻ�ﺋ ��t�wro��b¿ӟ?D�:�BS�e޽�FS*�m�:����/=8/	M�8A(F$)�ғ@<K�^z��O<��x�����W�w����r�"G�ĥ5�]S9ow��oѝjq���өx����{^:��?�.�蒴�M���,�PS��d�6���! b}N��4��vJ�Ȣ�3\��.߲j�s,���`����>h<F��$Ԃ�`*�m�V\W�hA�;Wd��s/..���'�l��JQ���iB.��]�$�(���J��w_�|�Q���hĂb��}iϞ},l�y��5?��m��H���O���e7<�%��:����ˍD��q�1]&+����r�M�Va���%K��%V�c������-�kf:`���(o��K�֫���n�6!r���ZSf��0u/K�͵`X��j_eh��;�&I�\q�\�3� �ҹy��#L�
��#"%�aNHʕ�+<1�jRrF�xq�ߝn��tG�SX	�F�䢇����@�<{��
@��X�.�!��ՠkxH�H:~����ߛ�����w�Av�s�B�E�|�b1�����Ƕ�I�i��Ե���]����q��	U�^�w�����>/���;]t���*\Qw^�Y�`��i�t��V	��2�wwɮb �]W��xk��nF,W�{���bI�8��5#;�=�k�E=�L�X�͓����N��{/3�gȝ.��'�M�p0�~J��X��d�?��x�N�:����8����0�<x0>|��G��")�
bU�X^/�ϰŪJR��ؕ˙�s�d��z���r*�����K����$S#Y���E�v:����[�����KJi�q\kJ*.b$zZ��v�\�����T�UZ�9�x�4nK��/��$�&#�*�&��yݨ9	����� ���Zӑ+�W�lYz�t3�i�6=cH��j��Q<���Ҕr0���aB"�p1O�s �9$�i�':	�{�^����� �f@s���S����]wޝn���t��d���.�<+ �W�7 ��e@oxp�}-���TU��<�3.������sT�.��t|0L����o9~��' �����g�u��й�f �\b閄��Obً��Ӥ8X�e6�l2�r�	�~ڳw_z�s��~�G�e��K�x[��iQ>,���m=b����� =jn�X����]Um�]_-�B�QQ��pL�le��V<�������Uv#�I̲E�4�[~/zRw�LC�t���$�'5��f�%�������W�vO���ӟ��t�5פ��,tR�Gki2�2h���Ϩ�(����|�~���{�I��?����'�u���2�?�IOJ��D�v�D��D ��\u�'z�o�&`�OU���Y.fim>M��4f�4X��d탣�M)hb����h �4����(�Ґw�7�G�RS]=e����<���4�NRk+���1�x��7%�Q���ZJ���1L�~?M9�`��Z�|����4�M��p��㭴o���V�mm[�)���i�g#�6���p�&�|Gi���-� 5O��<狴F����$(Yv�t�m�I��8��8!���������z�&�K�)����im6Kk�qZ;y"�'4FR)�i��)]���&��2.�i��@K�`>�N��I��8qPF��)�q�ۗf{����,5c�Ԏ��Y]䂽����ǀ,��8�~�4���Hk�>$ױ���<��^=���s���|eT5H�'��[�	�b�����e�zR��t|0�}z���	@��)�K.y�[g�ō[����D,���cK>S0%�Y�Z�[�=�7��P,��ٝ�\{�X��=�ҳ���/�$��M�`�Z6s�}D""UFW.KAG�Hgzn3�W;k����XZg�"��e�][qu�Հ�ɛx�*�3��T�Y�9�;�r$��R�$�˲��N��(��o�`E�h�_�Jz��qv����C�����:w��;�,�)��g�4����� Y��4��ҩӧ�=_�j:��7X���ӣ����_Ȯ{r�S��[}�.�lʱK�,�i�OiF?)Ypuâ�sIb!N�{�qMϤ���i4>����ԛl�H�OGj����p��D�*�Ii�yi��?�����X�i��JӴ����F�^Z�L��x�6(�k+-~8m}���ѯ~%m>�`�no���_�H{/xr:���yW\��<)��Gi����4]Y���G�Ԝ�f��fi�l�ֶM��������/��{w:���i@�DL��k������"�{�sR���l��t�����a�Hi�|Z�4I��4m���4<y:͎?�N�����wݑN|�i�y"�锽�iJ���?�wp]��&���"r��L��(����(��ޙ�ݝ٩�ڪ��c�5cY����mKr��t�u���{�m����s�s@H���囷��݋� $hQkJp�������}�|�;�AeG;7o�����	Y�`u�"p-z� e�f���qh�TEGA�PLV@[���.h"�fj��.��mB>wÏ>
��yă��BB.�@d��n؄ʮ؞ۣ���:��A�x�3�e���=w��5t1����.�ᒿG��\|�ZL�&j���[`�c��.�����l��Q�͉u����TE:�(ʫ���0116����
>�һ�|�+q� й�	��� ����c��Ѓe�ee�&QS*�?�x,�9g!�<1J0\E��Ű�_n�?����)�*�
a�/�!�t_�<ާ��{LiB�b���1�Kg���]�g���.�X�y�R�7�s	$bu�u%���h�@���ew������gP,x8HEE:;:�I�V_��uo�"�欜hY^c��'Z��f��j��t:�l6�hr 
y����������USy����3���>@'���S��< )XׄVHC�8����H�ðP�>d�K-��l|Ci��22�*U�����QӀ��͐kja)2lY��P���w]>nB��
�L
��dGGQ�r�4��	س��a��ˣ��+ ��Aik���
����F��Z�G+a+Q��, 

ttۄ��B��A����z6`�,$���PF*C�P�*!7��km��֎DG�W������p�&x��"�:�rY��D~h�yn��$g�2��\�Tȉ$���m�P��Y���VA���K�rd�,ܡ~�����TR�&)���֣r�To���K��3p<�\�á��h#è�mf�Ҫ�Lu���@����]L�/)Ap7w�Η� &��Dَ�_DP�*M1ɽ(e�G������-$����TC�m���6_b@�h0h(H�(��4圦����򅉉��}9����>�z�
�B:��Rj7��C li�V)Kdr�P��2�e���6�hT ���2�v���}�z9}���ci��|@���]�式K	g���.���)�C#
�75ո�硡!�>}���hjjBuu5���(fff؄���yk,�@�^bE!�w��T*=gI� )p8{f�����^WW'���}Yv�G?R�O��,����B����z��U<D|Zf�#���ӏa���P�a�hJ�� �m�?4������VQ�(:�d%�-h]�	�[�A��u��I�9��e����-T�q��y�q�wp��QdG�Q�[0l�m#�:�$#��H�Eu����F횵h�p5��p�H;T�U�J*b�L_@a�$ƞӇނ=:�Z�2j:�4�.e��Q��|��fTZ[��oB����w��R� K�`:6<���Z�    IDATDB��ffa����˯`����@�)°��R[�>��PX�p�w�4�#�f���GŚuP�Za��|��G��7����4����U[�p���؅�u�I2\M���p\�L8z�|�k���ޱ9�L:2��������-(�:LI���tЪR\�����nt��<���]����g/�"���<��"O)W�s����E@!j�%�(��% �5!�4�n<5^�<�}�����]«~�C�{���\�Pg!@/���b�y�V	��JaJ�.FF�en���τo��X��J������(��ly1@��%� �^~�,�'K�ʗ8��=�o�,��:&������� ����_u�k�R)�u���%PN$8z�(�-���Y;��<�B|�Kϥ|ffvN�K*yj_����c��
���QYY)�j$����A�Ώ4�$8$��3Q�.y�s�S܄�X�{�rv%I8��R�������/<�V�Z6$�E�(�}Nv=8��� ]	�ϖ���\x��БWttn߉��7�[��D� )
⮋x�ujg�����4�L�����|����
;RY��#�y���4X����p#*6]��YO'Ҕ�����U�?�$�G`LO"VHC5ЩK@���D���l��(8��*�

�8��J�M�`����;��E���˱P�Y��>�4��GKM#n!�&3
Y8{T���Bq�}�&\]����XU�bS+�n�+�� ;Z�X@��1���Qqf���|�����Ҏ�[�D���[������v�֐��l�cx�@�c��m�٦f��݌ƽ7�v��§uˋ"�T��#�sɛ�������'a`g	�@@]8�	��Y����F�$�}߿����ǀ����c���+e�����k .3��"�� =P���9�a!pп��,<�p�D"�]�_��W�2�:�������t�����r���<f�	�E��t:͠N=攑��,��n���g�w�ug���k���p��!.�l���`�^�6�ڪj�� #���17lXZ��xp�`a��_D��`Ng@�c�f��*4!eX�."����w}�>���F�� ���k��UΒ=��2C��&���ɵ!��N�b�Dnݨ�f�?�{�Zۑ��{�G�j���a�0��k�;�h��[�}X�*!�0P�$����J�5���l�AAS`U&��Z���{Ѱ}��f��ٶ��g0��cy�Q$.L ^��pL��EK�F0*��YH��O�6��yb**!��
��oĊ�ۑ�u�2h!��`���0��3H\8���g��da.e�Tϗ#�$2D(8q�K���t���P�{:o���C�\���o~���;i#�bKn�*��c�:du&	)�u,Tg3ЏǑ��8e��f/3�V�=�Q�e�����A�9kNXp�C/u���_dc���������g��&{�g�=?��ܛ<GN��RY/?�=��!����H��8�}}}��З��vt��]t���8L��FY��[�4�S��VN�ӆV�}g�\@/���?�~o���ޏ�6QC�� })�Z,B�0��;��/v��Pװ�5���,���Z�?�Ȇ���d��'''111�U�V����g���o��6p���u��k��7+\����#�/2p�7!�7��s�Ok�^+����==]�{>W��ƞ�
l�ԮJ
E�l���j��n=D9�g. 24�����g�B�YDR���.�K��q��
H�$� |N���/@ͥ��'a�����>?/�ȵwa�}ƆMp*�����IX'���?��~$sY(��*v��a]�1�D�0�^�o6Ͳa�`���U���✪�u�~��v �ƭ�b	��,���x�a�y�Y4�j�2�{6
�̂7��M��"	8��bv3gO#}~�i�"+ڱ�λ[�nC#g���S��~�9J���C����������W@�������FA�$�9������Ͳ�?ն�WT�b�5hٵM�v 	ţGq�?}�����
�T)�@���w}ۮ��j�(LE�6�uP�NC;~Ǿ�MD��PG�~��=�؈�ޛаg�6oFVӸ�@�΢�@�K��� ��w�:S��-]��ܽv���� }�}����z@���6 ��]�3�H&c���/�K��}��9��}�J?�#G�wtl���}�h�4]����.��.���K-k�!���qi���͖����������0��a��ź�}����u[��F�o���q��!��`
��ܨnN`Ku��Ǐ3��~��L���	l��ӥv�`J���(w��2�7�|����+�12<���F����PO˚2���V�����]ޮh����.��rG�t.��pH�d��T:��)�G�`���1���h�\�T녇YB���h��& ���"`�p�]L��"���&��M)"+����k�#��Yr1{�8&�x	�|щ3� �q|8zf<�Lu�6_�[6C���[ݹ0���~�l_���Pr3P)�W�����?����o0ZZ��3H���=�,f�}u���_E��I����~�-�c��d*[ Rc�8{����{{�i�k����Fш@���|8ã8�����a�S�P�,|��㟓|�lي��{���)Q-�Zf�¹��D��q�i���v�B���P�q�X5�|�ѣ8���Q52�f߅�S��lc#j�U۷#�fg�D�S˛�H����c8��o 20�:j�S�Y]C���=��9C�4hP���#Wi����)v�������Ej�s�ux�e z��W�����T�_�T�%���cc��)w�!�9tώ64�=�/���~���[���������m�ו�nζPdK}� ]�,�s��.����C�-g:YxR��U��U�_��_�b�{�9]��˼���~�2�ץ�͕��_,
���vMY1��֔�8p���M3�M����c��8q}}}\C'@�J��;s5u��(�B��E����O���=��AKKV�X���i>�ӑ#��z�*lٲ��<��f�ӗ��#\I#��"�Ή�C<U����,�C�1�ȯ0�³���$���O+?�{@�^$�Q����#�]���?B=3�x1���R#�6�@�O���]�]��o���/��3��{�U�g��XP��"0�[P��&4l�ս�p1����fP�ԛo`��_C>?����� �"���r-����Xo�B���^}	���QC3�V�p���x�h��f�j��/k���d��0�w��h�]	��̀����da?����."#C�qM�~9�E!��ށ�]{Ѳc����8��) )����C~�����vTm�FO/��f�1���0N}��@�c�t=d�o����ތ�믃�f5��}**��3������-D�GPG#|��j �ۇ��{Q�er��"g������'4�X�X�_^�l��?	��  ��B�q�F�X�0�'������8AwPS]5�����,�_~��gG.�}�He��K���u=�>�q4�qdڌX����(k�]�K�8�H�Of�}� ��Z���63�9zebk֬�Wx�k�a�^����/�/�i��}n�ە��b��v\ĩ��u�ֲ-��E��g0/M��0<<�;�gJ����z[!��/�`Q�O꤈�:	����`�L����3�S�NA�k����k�b�u��y����M*�(p�@��9@W�)����rkTuz��#�c/<�tɃ)�8]������ï��M�P��R6�b�I���@�C2O}�RZ��H��)4�؍�U� ������C?Eř~$�Yh��4d��Pz�aݿ���t����*�Dy
Q��*��k���S(z��$�`�.H��X�G�����<��3o��©S�2�f�%c0֮B���H~b;�x-�h��BS�H��P(���JV�W�`���b}�4
o�����o��?��C^v�6؍h�wj�߉�((d��i�jǟx��:V� m��@QS����w���`j��
���f��݃�k`���@N&̀�qi�,r'O��_�5"�㨥���0���#�o/���A��[��ɬ
_as;���@/�*%@������% ]�mY��o��/dZ���;� �2�u@���D���]���{���2t׵QW[sjŊ��]�{�W�����?�#��?��O�����1m�^˶˶%tr�
�8�
U��eszh���,U	��e����P�`�W�Y��x+Vt�f\�y�A =� :�D�����r�ˉ��6<|�]�#,�=^	@_�u��T'�ob��vN�}��9Κ)S&p�/�u���hnn����x.mn�dbn�S"~3X���i���1�}�]�ao�o@}]-&'&��[�n��"������uC�8�Pa�����U�	�l�:�~',ə��}�_|�d�Z(�6�4������PQ?b�Qߚ�<�}'q�/�mh����0��V��?��nE����p����Z�)��%��d�]sV��k�G��YYge=����n�G���8���5gϠ�:�CZ� �ڎ�w���k���F��gq��1u� *�"d���(ģ�Y�u�l��~����8$M"*<U�YȰ �W�T&ϑ�:@�s1����x�)x�����讅Վ��ݸ����ڻ`��c�2Lꔰ\D�ς2��)�U�a��,TH0���?tǿ�5ć��ِ5($��f+�k� ���e�/@"y�frȏ��ԣC��B�#�FB�)�z7�F�~�9UG*l_���,�c�Z/>�g@j�ŉ���"�� �|O��-go��y�<R8�������f�m����dgg�S��|����/�������u����?��{
�eI�M�����-}�y�>��\.��|@/�niP��D��п��X�?�K-��A������]�ݸWȗ�1��4��Mz_� zz��j�J�??��5Q�/��2���9;�uL�8e��lz^�\�רO:QF 6F�y�,�������r�ZKs3��N�����p��73���g2�ܶV]]���Z�(���7�o�e�TK�N��\	j�b�u�6�H���8������A�*CvL��̀кs'V��3����,J�L8{n���p^��4"E�DQ����z�����Nh�yb?�)��%��<���*�İ��;�s�Ӱ[��$������Z ���-�!�D�����IT�s�"6��\#��݀�];Q������xc/���A�v�� ���z�
�Z���B���V�@����:hqH�(<5
qv�Ѩ[ε1��{��8�Xf�����#��*�^�7�����.��2��0:9�T�dk�M|b(��g ���;|G��u$F�໐U	y�|L��RM�d*	=.1�/`;�3i����~�(���n �X�Ɲ�ݷ�[6#�j(@���P�Xh�ΆA�b�����G�(���,�����R�w��IJ�N^b3��S�t,<�>�q�vi����]]�O����'����r^�J?棔��O>�d����{
���E�(��m�������1Ë�|h+R����%����/�B
g���zu���w� j1����=�[��-�#Cρ����]��x%������<dg�@��p�:�,�С#����ڵ�1>>!\�
��S�G�l�܏;ƽ�B���AZ�����d��h�6e>����	]]]ܻN:Q����"�=�,�m��YVءζ-����� ������Z�B�zr����'���v���`'�\$�(%3��I�z�}�I��2��8��5䚞^���"���1Ʌk�054���0�ț>g�5Q}�ĶmG�[!WW��� �a�G0��Sh0�Pࢨk8_]�������PP�L5
��:�"*�""cC8�����@?w�,aV������k���C�M@z'{�>����"&U��GAA�q��a&�@M%�*Tu����U]Ыk!ǫ���!�1h�gq�a�g?B��iċY�hڵ-7��ڈbm���,3�fPG8����O�"�z�����U�T
��8�o"12���42LIFVVP K]*�Rئ�8I�.ɠW2\�G��+�7@c@߅�͛�UU���#P�8$1Ś��<��2 �D��r�y�^}ʽ�>�R���y@����ܥҞ�a4��q�������h��З����/��\}����ey�q����X&̢�8��7\�%��d��n�2�d�A|�B*��/�Ú�l+W��zgggW�-�����庄7�2�������~���"O)?����J����T��*�C� ��������}b�۳��^__� L�ڑ#G0::�����3e
l/
�x��X�۴�/w������������^�fR�6������߲��F��霌h��m�`(
�<mL�.�L�z����%P��{&�p�(�~c�>�6��C�Z<ؒ��v/G^Sa���L�U�n����2����n�Ʈ=��]��0tR�A>vC�>�3�>��B�r�Pm��m��,�>�)X����!2Y��@Բ��)"6>�����_�38���"[[��mhڽ͛���οwg^|S���Dj�L�ې}���tUt�N.q6��)�o�@9�m�����s��џ�?���O�0�p<3�8�n�]w}^K'
���,�iZ#R�q_�Ǻ�xh��T�q�?����=���@�e�w@���*�T���
�	9�^H�K�;ntɁF}��ę{�0�i���'���ⶵ�n����C��d P��tQ�����{�� :������=Vb��U�-2��,�R
���{j�\��J�T�l|�epf�G��4����XA��͏��[����X�����u��\>�:�H_<F��]ʖJY��RV����^
(�b�s����ޕ�p�����+�W�S,��r��KS�W���G���^l�ߥ^/s1�ej�ر�]]ݜ-� ����]�(r�Ç���1�x����t�RNh,#^'����N�O�cR�N���n�f�12<�f�V���PvN�>�c��D��� ���R��M<�S�D�,]!���W���cn��4����{䗜���6*\���sN�VE}�Dg2�8욦:b��%�I�ݨ�#*���� �<�9�G�c�'1���h'[Yx(D4L�5��s�Fǁ;Y��S�Ȧ2;ǳ�Y�c"9q���9ү���ID]yEF��
�uעe�>�\s-<)����~�M��Fqd�Y@L�	�ಃ^ 2�}��S��v�Bݰ�WoC��54��~�c��GX��D�"�:3�Zo��w}^[72�JdTa�K�82��8�3t2��K(����7K���{��� �Fˁ��OA��j�|�e���q�ҧ��������Q �zS=�}�Q�� }
zy��h��J�`��z����{zh�f���� X˒������Q��b|�<�W/�|F��{	�I�>�o�y���=��������~��N_zǸ��(Q�����ߨ_�/�l��\!�����B@DXO/s~���d���ʕ+���DgW�<@]x������苽�ǀ~�0��	�)��V�S�������O�Az6�t'�ǐ�:���}��!���b߾���s�P�<:����$��XM�i:g��4.���l�{�	�i���ڝ(}�]�,��ٰ�8��Ѕ���V�q۾R�.hwtZ������G,=e����č��*�Gē`y2��*O㱨��(�Ȭ�B	*-�i��FQ��:4��}�UP�Ӿ`�>r�=��/��.�V]9MF��m����;��L    IDAT�Ԧ�a�1x��t:IB�̣�5QI��~�̾�
z� ]���� �]���nD�'��� �A6-ȃ}z�E��:��⮃��f��E��
C����O�N���D%&����Oa㭷q6�ָ?�'4O�E�&��ǔC�7�������F*^�Y�)db7|�my	�٘M.s�$��,:���ÿƱ�~ɑA49dfk��X��"M����"�Ւ:���H1�*�48IR1kȒ���=hؽ��Q$�݉'�y��H�s���>��Y蔡��r_�"�	@�*���rvu�^�0�"&5�K��7O����2���v����1�u������nq�����K��W���}�bQw]���ezx�J����<@�D�|,�-�����Z�] :eib_��Y���?l@_���k�^���_��(���].�~��I��kP��}�8q���uttblt�\�?�h,��
���c|�3t�w�}���e��$1���=�Yf�(�>t��PM���cxh��y�W��;=���&Y��z�J��	�(&�6l;��,��^��.F���+�Or�p-$�3������_a��)Dߒ��T%�E��`z.�p�D�.�Y"AFni�dVG;�?y u6 A��S�8��c}�yt�*[��5 �V���|
w��F��[(д9�[m�B�c"v~S?�1�o�whI_�~�lu%�k6��Ѽml?�=�T�����ȝ;�铧�Evt���P��L�dK+�,��`!�ʘQ��X��&l��V��G�~��ӓ�,�!9ι@˾�~�.�k7 U]��e�ܵ}�������l4J�j��A����Q���p� �˨B3=�!E�*�p*�p�	���N�w����b�<02�h>�(��
���h2Y��ڋ�MW�@����a/|�eϳ�K��j��:Q��C��� ;�����39>�b��½�R�3�� �<��&�Ω���Ll-оO�~����Q]׾���?��/�������{׽/_,�a���\��{�Un�2'p(�йQ�2}a�p1�χ)��Ul,Cz������RW@��c@�.�_��h�Ů��6�ŞC�3j��+�,N�<�3)�G�O����NV]S�F$�b?y�Ξ=�k����*Jk3#����5t2�	���B��vp��Q�={�w��U�::��8��Fe�i�r`��߲�5��N�H�6*�)H����ÿd@o�D�9�C֗_�k6V����ɳ9��:5}�҅I���|M+2f*��6]��oD�����	���z�)tP[�G�j.TE���O�瓟��A�H ���3t�5D�XI#����;���4"����"�Py�'аw�l���9�%F;b8,ೳ���R(LN�pa�t
�L
��4"c�pΝ������a)@N�qN�aŶ��ݿ������|�a��#9;�S�R����6�n�~$n���3�G =���R˚� B�5b7\�ϋZ�
$ZT�EO�Wt�H	@?���C�CjxEE����!���oi�K>��<b�<�8Zi�4��x��9f"�����߹���1�uyr&� 30�k�^Z�,hka�"j��:�.���f9O��Ų��ٛ�$�C�(ߺ ��GB}K�+�P_��ʕݏȲ�W�%���П�y������^�q�-��rI����B����e ����J��t>�W�+A���M٬�����R�Mi1-�����r?��(lժ*ܛJ�N�;կ�����ۅ�+{04t�{v	LO�<��4=)�	�)s�~u�E�4��-��i&:����	e��#�6#
�i�C�d����l����}�i���JM�s�h[�Jc��J��9{`B{@��{8A���
�����$�/0��ShV%���� �A��w����*�S���"�N�@����?v��3,�"����㔮cݧ>��w �&���<�(ZM1r��\Lj۱v��)(m+��U"O�����]plj�>;���8���"26�2�):�h

-���f��܉䪍p-����9x��V���wE�4��|����0�ƛ�:z���O�:���G�U��B�ݷg��q��g��
���4���	�ƫ���
~G'
�$�h��ٲ�m�Z�jф��f�A�E����(d炃��4�cq��_Ct�$�TY�q��m�܊��� �^O���tV��T
�#G��߂6<�
�*�Eq艝�Ѱs��t�	�!�
��R�� ��)n�Ɔ�s���\�T���~1h	/�TA����pYLDӡp���0� �����իW>,���<�Џ�/iʟ?2�;��cǴ������S�L���R*����\�]���Ƚ��Q�B@_M.����g%�������MH�Y�܋��?L@���.R+����bV~S07h�w=L]�b#�RX���]�:��R����+�05�y�f��
t��ƶѾǙ�^A���o��E�t\>�iZ��3Ml#j�}�
D�������}
���3gY	��Ԉ�kV#��35�jݹ{��)QG���E�K}�s��y��\T�,�#�8�{�9T�٩����iEB��s�g��f8�*�F�l�����z^|ӿ~�U�%o��=	�{�a��7M�{�9?�0j.L!^�C#���
���-�P{�g!�uD��
�<�k��$�E0���8{U4�MRpA��mmDϿ�C��shj�j��BWLg0|�0�ښи���B�g	y��u\Ċp>���>��'GҜ�W̡��G��X��;���}(�y\x����8wuA	6�jp��víHn���5�������
ݶ����)���24�C���-��U��V�:�l��C8��� >ևF��- K��i��������֭��BE��e铍d2p���@ld���'�ܶ��}׍hع5��r׹u� ���b�n��Jg���Ҁ^��� *_��g�%Z�����~-kdx0P�&]� ]ܗ\6�n� �}-͍�^�~�/%I�۟���^jo�0���t�������j蜡��±5����P��ˋ!��4T��t}�<���X/�h>ND~2zzW�ʽ�[ z���"��wK�ˇ���%@�Թ.|-�\�s���������8w�<.��kj�����%�{||�Ej�u�����lz33��uMda�Bf3!���NtT�K7����;]��^{��o���esH��p�y�U��={�<^x�9��o۶�)z�9)	Mb��<y>4W�I�L�dTK'����rO��}�Q���Txp$����]����um�bIxDm:6d+��yX�����R�E��_d\��8-��س�o�	�l���o��SOA��Gb6ʹ0���	�m]���H��
zK3�:mrxF�t�fFꭷ�>�h&������"�{:����_��Z	ĒPr�F0~��������ס��JU���/�1�N�>���C���c����B�| i5���Q�c�{w��� N��P�PI�6��hJg/*�\��U��55@�HB�Ux�Y���c������zh�6!ѻ�����
���o�bc�h�񸮂�A��u�߅���׬��K��6�-�Hd2��őD|h�{ة�pVבmlFd�hؽ�=π.��=aBfa�Xi��\��m^�{u�w�QK�z�Z�����0�-�BhJ�.`�̤k����Ѕh�w]��6��y����?��=w9{Ǖz�G� �������}�|�j�NqP� ��/�W��2P��D:��;g"e=�eWz9����"���eQ\wO�%=<���/�K�a���rn��X�� o�c|�s @A#Yf�����	��o[6o�ig���Njs�7ղ����Ͻ���f+�0tX���M-I���Y B�L�X,�:��5���:OW�6�S'N����'��fE� Mv{啗�a�\��z��m��u"8���Ͽ#�,���@G��h����4��a=�+�>�$�l��,���|������7��#|\�>��<��ga��҇�xz
�7K��2&�:n��w������)�{�5�_x��)���|�%*ߴU�BEo7���n&�|�νw��N���gm�3�����[����
Fc#ܢstC����7߄�I���
͝�h�|5"͍�*b�HO�ә��s8�싘x�5�yED	��aB�Q��h޻��WC���=u����(��6��c�)O����bZVa���r�jԬ]���;��i̎� 50�|� ��	���;:Q��j�n��l�n��yo�+��0����A���w~�}�i|j1�,�T���*��z�(���s���g`6b ��}�~�Ӵ��[�,���&Ƃ��6J\R��}l��k�_�'�񤂹u8?����O)3YNp^�A>|~ɻ]���0C����6<e�����R��>\�Akkˋ��ĵ�,��?���5��=�J?�#���{{�~�q�{��l���q���B�MڸB@�r������ԝ?�`8�r��V����s�N���0����b�{x����r��%@��.�]����49lqv�"�ͳ�	��H�j�d�r��7"�/�ܹIΤIGj��.������0��v+jk��U�V��y"�\o-e����@�Lch͐ب�����/��z{��q�LNN�yd��Φ��ى���4�������9V�;m��)�6mE�㘊w��fR�F���Cz�	�Ý��UR����-��Z�5(+$��CL�`�f`^8#E��4DŃd�*[CZ10�F���X���kt8�2'O��_�ѱ��!3φ��p�H�F��5�Q�-�$4-�E�Y��tR��Q��ݻ�{�06ne��ԩ>���Oa����9�Q���P+��k���w߁�����t!#�A,�)g$cJ�@���i�B��42�>����ԛ�����hЎ���"�"�t'�[��x64�`F�f�[0=9�5_Y�B]#"���?�CT�b�?����6;�5Rm���Rud�ZQu�'�ܶ��5��4��|�W�ļ#Gxz�o �ź�TD�ls���P��з��s�=�%Ū\������T�����r��Y����f�Kz��4�7��ް�$�f�gz(��-+�Z�ݱ������}o�r��+�؏"����{ҙL�q���I1P�taĐ�R��>p^@���?D@' ����)[
n9����EK~�KqY��2V�ǀ>�������KL?��^'Ψ�>=Ι1�����X<Y6���d��r�z��i�ܹ��e(�&KL���c��[����'\��ln�~�l�V�[6V�h�́[�N�>�t:������!�3��cvU�G�﹩��N��P�SZ���;�0��f!���?��SO��z�)� ���lD4u�x�+�AY� ���A.*7ΑPg/�\�f�
��q+�n�;N9���9���/��0~�Z��>�o�c����Ɂ��yP�sB���*#� �X��[n�ʛn�]�?o"{������TsP<~J6�KfA�Հ
��uy���Cg��Z/H��A���}]�@>Y_U�XE(�}��y�IT�L#�/���P���x;�ѧ�)�%N4�&�7��}#�Ħ-hڹ��nGTѐ;ه���b#�h`Q Ms3�onE�4}bk�"O�|$����[��@:z���ućF��4)CC��꾽�ۻ��T���<��Z0��Lpg̡}�b��lCC�Ҝ�M��+�C�+�r������2����1��)���).��Q���ԅ2�)�'���U,�}����{���:�|��ߟZ�|�������G�u��I����2�+4���}�zA��de^*C�G�p�$v�Pi�K{�UwwS��D�{�{0W�a�.q3-�uq�Y�/v�[]AYi�ۻ��Jz��G1��x/>=�%n����jp���8Lm��=b��7�Na����&9r���4�L�T�:u
�Ξ���5��<�5��3Ń:D�@���ӿgR�s�V-��I�r��ٺU��B�����>��L�[��0�(,�~!�\YS��e�⪄�2��	�:�h�����H#�8�˟c���ѩj�������ڦ�u��|Q��eA� E���Ú���xz�x%��fTn����#�e=�˃���|�]�{�uL�{�粐N��н<��"�%�}�2zEH�K�	�c(���ظ�{��i�6�m���?����ΩcP'��J��}�e�Emch.��:���$7��'Ѣ*!g�(��"z�5h�{j�َ�*T�k�&&_{	g�y։�P��`�
 ���&�p�_'��œ�<}9��($��WU���;��;�1HE�Sx�[߃12�z2��l�fK+�n��;v"�n-2���|%r ���d�;���&bc�h���8<=�T�Ⱦ�hؽ՛7���O��z	
xBG=�T��uSnCA\@�S�#Uп�mkԎFF��s��PԨyy�ݺ�$��=.&�-��K����K�O�������7mM 9�⨫�l�)�*�����M7��C������%ZI~�_d�-��x���M_�<��l6w��DL� ���
O,�y���9�N.B@_���9����D4zCU�&
+�,���dKٕ �_n
P�yk�]���(���L��h�viq�J��Z
�i)u�_
�]����h����)S�.<{q�K5�����(������e[<Z�l�f�8��I�F��Tj�b������̙3سg�����'�6v�5'K�y���܇n[x�wy�$:���}�?���Ν?�,`۶O���DՋ���!����7<ؔCE	�b	�C?G���Yd�Μű_>��'�@��"a�0L�Ćm�HMӬ\��.* kf)�5RU���kP�y3j��Zg;��J̸&$���<$�&�GN��[�a��a��Gs)�zy0"�ϴE�L�M�R�u��(&��;�Q���|7"�=�jj�sehdW[,g�~�-L���?=�E��#���I�K�M��	0(��T�92��LBkkCb�:��t3��n��H�*��>�@���$
�C�~�=�{�̞:��A�z�i�;��ϝD��� 5��G٨f�M7�f�FD���(����A�����<:�ׁ�"olF�mw�~�v$׮����q>���T��'��_� ��8*,]��X��ݟ@ˮm�ߴv,��/�*�nui|*���%ː���� ���۽��/~	�C|��$A�d�#ę��"4GGpp}�}NIDW^�
}I���,"�� cHp�&�*�Ͳ�m�>���2I�Эw����)?������/�Wn�������޽���ޓ����*�
ӒA�؀����"���,�`��6�U/��V~螇��|����r�j�v��#��o�z�Y����1J��M� b�U(Q�eUR�{s0v� 0�$.�=�♲ܶ<�� ?_A@_�s�=2�������y���{�`c�z|�{R�sݍ>;QV���X4y,*)؅�Vb�[}]L��^u�ȩ_�|�o��V��ՉaA���D��ǥ͇�F4>�<�j�Dh,j5�k���4��C&����'PYU�7���K^ü�)���N�Ikbu|e���'�� �r'�lDs9�����#����Ϡ�۹F�i���Ŝw��)���N�ѿurU��F�=�H��"���}�xy]�I �%!�u*g�<.�@����>x��P33����9*�
���hT���n����NT�\3�D���M�smD
9��c�!=2kt��p&&!��x��ϯ��A���V_��zg��n�V��[U%��	�)�s}Ty@̲���(��Fj`��(c�p'�����B1��*1䓧��L"��rw��ԭ^��H$�D e�(����_=��*��Uv�VnW� ��:$ׯG�c
*Mף�/>�(e�G������<�B�,~Iɮʰ+���A��UHt��4t<��C�U�U�y��S    IDAT��O�N'�f@g�y��� ;�?�p�>�Ay���T9Q��i�y!�h9�,�y
[�.�Wp6/ }��B���9�W���[M[kim�ŝ������������op�I9@o��x��3��<�c@/����tN�X��T��?�`_^�#�𚇏��t�H��կ`ժլX�)[�윍�Y+)6j
J%h�	��RR��Z��
�|AF������@8�#3��DK���g��Tb	���n����y��zx'��R|D�TXT���������y���}��+�������q��Ju�Z[�8S��sx��w�T&�b����N뎨=R����?#o$"�����u�:19��;v�����@gfR��34�� 6lXϭjtL��%��܉.��7�b2Tr!�
���+P�u@S�T�F��7-x��p��W��Ư�I2�����%���5]̑v](�n���4�����k� �a=��z��8����0A��A�e(�%GCR���f0{�.P/��ð&�C*�Sk�,�w<��]h�p�6_��n<��`�8��"Q.����g':ݷ!�Ȝ<��#�0�?;��_,£��t)TZ"�����Er�*��-p*���e��;������'�XP-r>��x��P?��ǐ��b@�5������Ԣa�$6^��y߅MɁ�C�T(y΅i̜89�F�w�}��nE��ڡ5�B��B��{.$��A.�f��C�[H�42+"P�ֹ�J(Ր�+QTei���C#���V��nĮ$��s�-�b#����A���_�P�0:=��E�"S�������T�S�2�}`@�E9Hڟ� �:�G�đDq-�M�������?�eF&!���0[	)���J�r��|���Ώ+�$�A<�9|-��\��ގ/����K�8��d�m��
:�OE,����y�C�e�r�O�1�!\F�/
K�/�7J�R��m��\"w�+M\�񤶺r��k��9�VA�4������r,=�*�K>>8�a�
QY��e��>t�u�����È�p��Dbs`M��Z�4�|��A��SM���=���D��������Q��9�ؼy	P���%�k��IUi��bH:[|��J�ޕ��p�k�Fц93���,���6cj�sx�h�ѱd{kِH�N���]ӡ�Թ�j:/-�~�4�[&1m����Vxԧ��1~6/��O�&��\����P�u(�$�dj<	߈�V���(,��F ��:@�{�q��E�4C]� s�YxY����g!Ȁg������[�o�����u��,P��ӷ͵���L�I�?	�L�����4��K��&`1v��I�')0�-�iB)�O|���*L��O���|�@�+2���Q�}�d�\rE�����14!��xdt��:��C:>
2��"Y�+�5�QP½����jσ�������Cb/�L �p�J� =�O^ �K��s&1K�*��H����91�B T�!���!@oi�فw���y/=����˄�+��+�^��Z�`��禮�B�]H��6Sf*S��^I@/�pA��I,t�̩����g<ƒ6������Ǡ<���s��}�a���d,
?>A�ӡ\� ~Ȇ�{ cs�B��p|8�>�7�zq���ayK��K7��/��KU�2#t>΢D�Ǻ4�NA�����
n�k�`q\V�ŞɤyH���.2q��<����~�&�Ӷ�͠�e(O`s8'��>�4����sL�ӿir9���im��=��t^7��uǫ�J��T�P�$&��,����W����A���K�//���"J�Ms�Y<<��E�
t�0J�G��J�sM�T߂>�*�b.9��%���O��M��mS{Z�ڱ(����AH� U��Ѵ0A�l����f�S�����.��TgC����J�7M/#��k���
�q��g�9��:tO��9:Y�H�G���:R���T=�vh���sI�O0Waw8rz�H'�˜)�.."$6�m�0a+\�����!	�qH��O�mr)6�9�����|��HaA�)�Qp@�>
���l��4n7�g_��)C�����z��1�Si'��9��Z��/���Ϳ��Ιn��ez��gq���g����`Ϣs���{p���\����N�M�[�,K�1����`:	�LI0`C�8������ܔ�)�!�ӱq�6�*�լ�#�H:���.�?���͜�t�u�?�#�$�ٳ�׻ֻ޵V�'��7_��������Yq��F�G�&�	���:
����]�D�p����_7
?��1 �n���T�9�/�_��_��sנ�@])T?LSU�lH��Ѝr���бy���>�۬>�li�G��W#��o�k���Y�.���2;��:�^}T� H�9�$�ME�4�L(mz"5�y�z8q�w�����,`�.q�.���xFz� Й�D��za����u_F�\��&P��.��<m�� �[Z�l�R��NkP#��Ԯ@ ]>|�&f�g��d5I�`I���D�f��j�Y�'��6%e{��y�����)�뚩W~g��L~D@POm/�i)'�� $�p��EМ&J�/�����G'�����Kj�ݛ�^YQ�.����%��U�Τ�e�\�9(#�C�=jYKMD��0�T�P~�k�I�M���O�F$L�	�"�
rs|Dj����؄�}�� ���I����&��K����$M$�A�ː3S�q��s�(����4-�!����1����\"Gמ�g١�F)�Hd�4��F��Ì�'��	�%M#��iN�G�sĖ��㴫�D�"������{��H�t���N���2��K��+�:��=ۺ�iSW[겖ͫt~׵d��`����k^���2�n���۲gn���� =����d���_35iy�S���[Y�ksɥ�O�dT?~ӟc�5h$j��N)"�J"t�YST.�R5�^/�n)q��uH��)VD�^ٺ�����N%~����4��4���[��U)�M�mu=�н�3������|.;�D�Q+��,d;<xX:ŭX�=�I E�M�05561ENk�wD�uOkȐd<�O�HQ�}��φ�`�Ǵ47�XH�>]���#*�Wnr�L�E�!ݿ86V �>��k�r��4��V�E}��
j^C���YG����y�T���K��K�؊_�����	�t��1! �3,0�̫�ZNQ��y\b两Φ�7�}��gǂz��x�K���E�!׀�6,�x�=]7�;��F��Q	^F��B��TF����-U�ؔ�&�:E@�N��U���bZ���:T�cN��)���xt�i�v�l�ș	�BV�'���d潌����9�%^J��F~�Fr�w�%�;CN]��QĢB�dv{5�+`;���?�}�J�3/�_�	z� ��� ��>�=Bg�M�j��w�"2�R��ٍ65�U�����7^����n�ᆉg�羧�D@粵���&�C���Z��`Ƚ,��s��-�Z�����Z�R�Q+Ώ~�cX{�Z47�����%o^)w�vmu��Ir���$k���5�t��qڲ5C��jR�~��d�-�0B����.�*��'�6�]�%lF��
�m������4��6�p��O�H��FFFXG� �r����I(GT<�G��ff�<͍�M��T[�����qAGG��sVD����O
��, ��l�D�Dթ�iN#)�m��̷T:���
2\F���K��c�7]E<�� m�� ���m�r.�(	Zȱ�uCK�d�x;���]�3"Q33 J�3H{���!(�W�Wy:E��?h�zV���K�l�A!P�(��x��g�R�W#Q{��hLj$�@�(U_�z���F��9�ì5�%Pa��x\�O)���I	2(�s#����gzV2+�7���IaI<I��`HȬNTA�ֶ�:�m��D�����ڍ�}�F�}j�qW|�.���%{��kI.�tzmt.���a΂2tc:̐�B����,	8y�JD�Y��w~�w�)��7�t�M�s��gn��H@�T��Э�Ǣ�����k��L�\�&�����d4��ȟ}�ϰv�:�P$F]�D��Py���3������"��ǯ��l��� v��S���j�~?�6�ǍC�8�lf���O����T�wF@g�g`�6~{�s�YƙW������8U!FW���}�J%�T����	diM�g���jݨhMUN�N�;�N�\8���i-�ff�Y��g0�S�}����_�t	S�����pgJ���I9u�n9M��Pu�h���Sk��� ,#���Δ�6ס�C�gu;9$:�52�Rd�X��&�|bW[���<�8Qq�!��6���h���hJ:�	���4��#Va��f�{B�Mg�q�V�!5x�4���PH�̀�����I�X��-�)9(r_�Y�C0΋Ȋ������b`����w,h%6�@����q�Lеjڂ�ce�%���Y�Hy����[��E�D�Ss.b'���@P�����	��HG�"�h����䀵��Y�ƀ..�!��v�c7ހ�{vk��	��@��b@g祺�,���C���j?��P�i[��5��ǀ�e������}��k���t��?���g�羧�`@��:t�e$��,B7�e^h�����{�^��3wYێ~ǀ�`>>�q޺�����/Qs��h�*��EcN	ײ�s���$�i�,�E��9�Ο�:��}�m���i�dG�=��?�23�	+~FpwA��6W�8������c�yۦ��]݈^�
��陗�e�X�?��љE K�a	LL�F���ű�q�['Ц^�,z����0�S����.nPC�/��M8:>�hdMX�Z�,D@ʥkL�z�_eOO��F��v@�	pz���[#E�rL� W��%ڜ(n�ɑ娝��H�M%l��8`�O��T0*�� �����䜽��ef���hti��"��}+��3e�)���
��������һ�r�+۽#��9!2Ԇt	TF/�3�(�2�Q����q�A�"���� �G_~�S�bx輞�%�N���	��:��ʊ��E�N��	3y��M�5�+�A5�8������%�s����������קN�D�"��C�D�3`syz�����=�丑0��t����*w8�k�ܴ�3�XAT���ZʝD�wQ�������g��泀>G'd�����G&���Mg�k�t�Nc��A>]�n��nc�n���k@��?|#֭[���t}1�� XƉ�(YDBvʢ50����'a�:1%]CG���l���s�9>�3nfրhȄU9���mP�5�xWٞhyf�%�_g��=��K��k����8�D&��j�.�8E��h���8Ϫj�,��D�����'S���'ı�pŢ�̹a���A���HɄL�w�~H�d�`9�%���%}�5�uqtɠH�m���U(	�#�{��'H�G~�H�Vr��	�)t>�;�3��������?��HY(�b(]&iH	��I`F���Joy�2Gߑ|?��mQ�R�D�t�a�:`�Eq���}�=6�]Dc�y�)I�逸*]�)J(W-@g`Nt=C�iX!�,
�F�TVF?��cGD�.n�D�퇔��>�;W�E��l����L	�bjK�&JZ�8�4��y]��w��~?�=�C'��}&��t�<������m�U"�z�©=I��y��~��o?�?-��d���a��ɩ�W�ny�n�+����kA�j�]���mMNf��~�7�����N^B�S��D��DG�喚��-g�Z_v+-�ZN�xۍ��D�ꎟA�e2���V���8�#N ]�ޙ�?��k.��X��2�b*�����2IG�ӝ��Vi$�m;�r3˷���5) ����Yg9Y��ڑ@ �T<�">��d���G��s$�$�p7;���}���T��m�t�J-ˬkcM�),�)��]�,0s��Q���(�G9����4{�Z�s��QMRڋ(�-�u��K��  ��H���0�ov�eB*i�G|/�?�n���ڏ�t%�C���Dݭ	n|bQ=9V��>�ũ�G�"#������>����rl�q���PE;Y�{�v���~T��Q�z��e��柎M�:B�$ΫP������������k���A�1J,�Lt�t��;a?D
�����u@שQ���5'���X��ط{n�ȟbߞ��NKs4yG��4��Z��hW�޺�͡�������Ŏc܍T>��������7�CKK˓�~����l���-���̟���Ȁ�����t�݅S�ѹ:7���hb����j�T�"�����R=���·T�����zTwv�|j*Ց��v�R�,:��}���^�Run�[�*�s=��LΟ��,�8b��uE$$.mS��}�,���u���r��H��vv�~*�^^�a���w���j@'�+���z�.�17+rj�?���w�j�֋���킂��!j �2@K�(J�����IbgRv$�p�S[�(ϧ�����v)��&C/��4መK���M(Y�K"eID�S�@Yqv(8ʤ���2�µ'<�m�~5{/�W�Q���F����GG��HtΏ��	'	Ԕ���Ǌ����rBM���砿�k�(X�i}��[�'����d�#�G��,
��4|M�h�7_��vX���T>FU<W=ōd���9B�[:,R���Z^�y����48}��ﱾ�̐�8�L��g@����)�n�+#��w���؟� :q�����R�b�	�{� �~���r��t�3��ގx���������z׵���R8�su/���H"��Z�����A$�Q�US�6�m�A�${�.@��/�C;������oD�:z	����D�7b�@� �S�e��X]�?�{й�V��v�=v��c@��� �Y-����d��F�1��;��wl�����Ki�L����������42�m�EB���>@��r�ђ(���e���:��g����+A��� �ߦ�����^���;7�O��H@���pJ��0�|*KS%3�����=iv��3������4�n'jXՠ���=x�.��ѱ�1�V�isP��%�\y��
Ո[/�o�a���u%�l����b:v)��4�Ys����ў��mJh�VbsT���K������T���0��s)9V�j��w���*(ӠJ���"q?/���E�vK�qT̓��s{GL��w(V��C�{i��0�ԑ ������ٹ`gK���y��8��~��R1 �4�]3���r����	l΄I�f��3{*@g����%8��+ѽл��4�%�������|�u����D~�M7�����|���a�8%�΅�.к���u��k�}���g�Q�y���x-�Ks��-X����p޺h����'ce�PĮ��D�f� Hͬ�ؖHŋ(g%l���z�,� A�v�A��P���Tq�Faʮ�X������q-���蝢���9Ci��(i�Nzqi�X-����Zg������ȁ��.n̫�p�Z�mLD����fA�h����!qӑ�H��єs�q��9��r/���"zP�+�(B��ה����@@�#n2\
�|tt�-�jf�_�gFs�c���D=�%B�-	̹����C���1f$a_�\��9t���KGy0���CD#��A��p�N�QBn��m��y�kN�[�JL��w�Q�ֿԭ몳�2�vu\/ݯ������هX/ �<f�(��HVn���m*w�aښ��R�;��V	A���(]�����4�ݲ��u`���5�:p��'�M�;IJgK���I�^�ify�FS�$�u�&NB:�@�RF*bՅj&L�Y�ڡmN@a� �Et��Z�.C�@�cR#!m�ej"�-�<5a��z{>�u��l*�|���?��#^    IDAT3��|&���ߞ�=��#�(�qjj�5{�bP��_Sl \�U�֚�:�?����^<t�/���,[�-m�2�RkN%��+�F�X`$��j(j ���P��DA9�(�E%/YJ��S��m��h�(�&TZ�d�,�sI����<����W֪�.ӛĖK�~U��ۿY�f��zT�ĩ�eU��vͻV�;�p��0L��:����vf�y���'�����;LN9]���ߙi�@$q��z%])�.��u�� 0�j��+��v6̒��|7@w,����ȑJ�����TC��պ.�C+�+~����1�	�j���Ӣ�Y�4�+�-'�B��\n�1��.�ʽc��k��Պ�w}ɛ(�:�����`���g"`i�AN%��U|l�Z�6�� 1��@���u+ʕΧ�B�J�w6~���!�F/�z�3�Q
�0-�nr~����M�X���
�b�����>O�K,���6�Z�.�-A�3b�F>�'03�i�Ѝ���b�N]!�W0�?n�^�rw�t.�<����qGu
Ϝ$z&����������Xf��}��i��������6�Ы�zT��z��z �A˟9��8�:]�A�m��r����=�}�Qhn���\:��[�Τ�.1v�Q��oԲ*-9���_j�X��6�hbj�,���^���NY�!�!�.E�x�yk��T�PY���H�"�"��u��o@\�T��[K�VE;'c4�9G���K�^��m�V��'KJ�P-�c�q?w�]��>O��(0�>�������u��*��l�F�V;L5���#+���qJ�d;tVY��6+;2%�0H�T��*ۉv@w׼,�$*�=�������ֵ�f[�����m��k7��p�*�cZ8��%`U}�v6R�6+��<��X������@R"_G��
x�%��Ds����=�O���-�3H[w:s���]}�)!4�Ez��,��^�_��'G� �C>"��8�)٨��35�")�dpV�h�[�~R�Z�#�{�d�W��,����%*{�D�/b��	#6��{����u�kΧw�ŝ��Ŀ]�j��a�859�nz=cI7ܦ]�Ƴ:�����B*�\��VE�u���K�'���Ӎr����)�" �	|,*e�օjmb0����H-�3���8�Zhѯ8:���ذ�ͭ��X��uMPl�j���P5���/�9�@�2��Y,�r�����g�D�U��)����9��[�8_4a���;k�'Q���uN}x���"B����#��Y]ڣb\ٵs^V�����Q�ʸK�*k�&�N���K�����#��xF�_l�8�R3�)6�J��!���.�u$����d�Ҝ&�݊����ʔ�IZJ�ȱ�]���]�DɠG����3z�ڰ���u튔}V�mRC��W	�e�ʦ������N�V�I�W~R��t���� B^�qI��=jf���Ψ/3빨����^璋�:���̍�4�� �(9tuXY8��nր�'�˹���.S�il��e���Ǣ4P� ������-���%8t�F��n��,���і���C�us-�3=��i�ts�g	�Nsz������ �G�iAԴ��n ����YTm��$�e9	��^�#r�nR�b��E��R�2�f0@�m��Q�-�S^�XVsD-)��f) ����%�x��&�x�~$�ǽ�8�r�qm~=;��J^{�8V_��*j�D\3{�E���a�g7����ԡ�}�)�S�����3�hӢNZP��g���t�߈��*���ʻ�����#M���	h�[5��6��4B����ut�d+��QuA�V0���6(�kÖ�Ap�L�WE���A�_���`oט;���q͝��)�%�.:^��ʝj���v[G�Z+:�?���^Ĉ1��'��k�%˪�{lA����ISr�=��aXl�D��8-3�YL�<�5?���'��'@��/�p�ъ�{�ӼYu~�<Wg%��q�4����X���Ի?D__���'�}�1��y6B��"@���ɉɎ(Q�= kS)�[�j��c�-�u#�:��{��Qx]���Sy��6D͋��^tZ����h��e���%HGUG���Ešo �|\��i������dS�%���g�"�z9�ڣi�:ޓF�UgŬ�D�1�+}g�� ��j��U�ql���e��Š�|+>�ٍ,fq5��<�9�槷Gf?-�� �5��X�ǯ�^�_Ɔ,�l=��N^��=CQ0(T!�%#[w3�
��)*D�2N�_]�A˿e��%����8U�pS� ��1�V��XP�vh�'�#�F�~�ֳE�yǜӰ�(2�N#~��6�f�W% ���޾c�b��@��&R��$c��Z��bH��%� &(8���pq��=sƨ$P��W[Ê$�z����?�,34~S'7#�G�R�i�����99�
���I����>� ���tW������3P�t�A�9����?;<��u6�~�g�[,[u���0����DgY�8��1%@��]P��ު��8J>uz&@w�#�r�A�B���\��bLӘEjK/�
P\Cm��z�FЬ�7\���S륶Y�4����:�6�pv���E�ꯙs�@{!]v~O3��p\�5��%�5���j�u���k#�8�V�č^���صU+l�<u&U5�p�/�8#���pU������	�m�
�$h�?.,&'HB�x7t3G��p�gE�*4#Sж+ۍtz��r�V�.uNä|HH�X�ɺ���������Q�I��9{['ڴE����V�����q�0'��i�����G�+i��{�9�-�li	R�pF�+�@#O�ng`��']��ST�j�ϩ���)�<B�v�^����B{�ncR�KD��oǏo��n��q�
���җ�S��fk�3:�Ρ���1y�q��!�@�;�k{-�:_@+U�N�i����q����\S���U�MM��!�Z'=C��B���������?E�]gU�s�� V���?	��Cc�c��n^�{S;�ݭ��K��f�&��9D�s���X�~�Q�B�(BoeQwK{�X�Z�kY��?��_��$�A��bT�8�<�uo�f��~���>�����vr_|NZsϿ�Ȍ^j��&��[+��.�Ŕ�'���zw'7��c�ex�YU�|""�ã�u��<��!vLlo�Ap�^�A��1]�v�m":��Ѫw��1�`U�ޫ/]�K�����u4@����G�@��Uܓ�8���:,�-#΂��n�U�'�/�>��@��o�F���Z�������{Q�p��Oױ\���� ;I1�Lp>����uR��4�5���s�^��Vˑh�h�5�.&�s�q\���������c}��t~x��h,l�t��&���!π��Zt*IЅ���S��;G��u��z��e9%ok�ר�WX��h��ڠ�m���������������=�^{m�i��3�q=�����f7�~���ѱ��!��̦Z	u'ޕ�?���c��O���s�V�o�}R=1���Si:픤jp���w���Y6S��Ua
P�i-9F+GѳNBCmE��H~�h4�<p���F8-2���[�����T3 ����2��S'LC�jQkKY�F�s+T!��"��8ۨ8qvd��Y9ʍ3=h�R�Op"�� y]4�WS�����{�L�^�d�x�Ը.���v�q7����U��sz��]N�qS�W]Ob��V�������J��;_�ԗ�"W����R\վ�z�1�\u1I'��ڏ��(�*D.��VXTq_	����S�eo6��'�4��}��W���l�	9%�|'vN���\]'����|ܦ�'��<wO�;Ho���e2l*�E�UO2��ş�zH��XV���謁x�hj�*[C	��8fF���3�{QV5�!�˻����x��Ũ/S�����vR�{Y��8��u��;��h{�Juz�{��}����46f���9�s.��0>8:2�E!O5q4Q����h��b8�/�ٹ�y�Zo��xg�=7H�+�Cw"tɉҌk_-�6��6�f�Ͱj}'��)�B/zq������kQa�}�8�}j�P�-2�+ԫ;�JX'/�^z
>�(���Ec!� L��e�*E�6���S�쵱�5�Hw�"
9My��d�(1S�f��)�2i��|���IZ�9��M�,�1#KEL}�%V�2R<(cM47�MS�.�K�A�s���#��G���G䤰P���^E�9�`'������3���%�8_�q�n�)ȕ�4���[�S�
�>���!b�Y��.�����?��4�<�D���m�MNV����� �1���1?�V@�8�M�^P�񳉷uT�1�-�U23�̡,uU1%��+%U�����E�����e�o�#kU��U����@���'���y:`n�_]@�(�7W���B���|r�)���� F�W1.�s�݌��(�v�^��
ug��!�d�(�>/<���W�9�"��vI{j3�A��)�٣V-wE�It��c�Azq���Z^�PjD�x���)�L\!��������gr9�;�O��F�)B�����6/��w҄��j�-y����lj#�3�j�B3@gQ\CR�6�.H�*��/��t�S��Y}3����&?�z9��TJ@0�L�G_o3�,Y@��>��G1tlG�G)L!�
�
2� �w�4��R!�)��4�_��׬bZot|���ֽ�� �7����h����*#(㜥p���8g�b4�
���Û�b���<9*�#������e2�\>k׬�9������٤0>6��Ol�Ïnö�Ge{��5"���<}Ͼ�\z�Ft��)�q��J�����PFCcSر� ~�ӻ0<1�J� д;�&2�~YE@�?����1���Ϩ��}�TW�BTXS����N����,%B���{��h�IN�яN&�ޜV���љ1%��:�3V��Q�&i3�^�PrE�B�@�D�ҔF��~G�'J*�\��M�W	����/>o�aE���+��l�xi���ǽN���L����Q�������T��ŀ^��q����{�k���'cM�[�/Y�� zl͉�8ڇl�RƤcl7��᫔�|m��i��e�Z���,����ݧ=x)eͧ���(��
/8ɀ.��!6��J�N�$8O̹v
XB��W�F'ywK��vֺ�S)�-��٬�А����$��IWA:Q�2���F�����|�O?]��;𾗾T�$����]���sxZ���c��st9��r�� �QB��y���kӡ@	�%�N*�>�r��e=/^���St�9vr^��Qϑ@�}���9�U��c�����-���mm��159���	�b��I�=|����[����74�괠�!z:��9k�q�R,[�� {lh���7��+�3P��N^%�0
2D�B=�Mx�K�v�|�\0��]�{Ke�9|�w��cO�����0]�e@�`Ѽ~�]�l\�eK硿��|24�۟��CG�䮃xl�A��C��.�!*�!��/�5W��[ДM#G`Z$P&p̠�����)<�e/�x��pdx�5 \��\����Sa�DK5�+�Zm�?m�����)dnoj�TU$�>12JW�]���i|D�)�m?k?k ���@��NK���c��4F�*g(��k��5�qA�L�����%
��%h�`��Q���k�q�8G_�	$*���s2�@nX��@n������kcG���Ve��0P��ݥ�g'���W<�.>��k@�6�]ό�����\g̞��8R�X��^�H?9e�:������S"��?dg��a��S��I�R�nf�_���V��<M��R=b>i��j�j�o9Z}@wS�q��J1��yX�����&XC,:!������:�;?��?��S3����{���z,����5��\.� =�B��]OKl�,�d��.'�^O 1[x���WQJ9g��7-d@G��l�-<Si�Й&N =�Ϊ����>�P����K3h̄�p�b\u�%����A�x3�%���<</���O�܋�݊�ߵCc%��r)�p��-Y�Y1�}��jI7��D]�p`p�?����w1xrF���D>RV�H��y(�!�{ڰ���x׵Wa��.*f��s�\.���&�>8��مo��B�HB�/|��x��^������fLN�`xx�\
�m���`j&����o�>��:���	x�;��J��mW��f��156�U�� H�O��������ű�IT��@�^d5�E3���c���"��� W:��9)�����jz�I�Ȁ,e�D_r� B��=x���喿d�<r
D�ͭ�iAF�8`�Z0�����i�1��C$���5Ki����t	ڈV�z`+����e�X���)�$W�s������j���Vp���Yř�[1�N�C_�s|oU$f��:FH�htj硑��#�j?��+�R�Wy�����r
K3�|�\-=�:=
��0���vf�Mri��Zp׫��\���_�����s����]�ƫ4�ѐ�"��WD&8	����Pc���=��� z��d�ԵB�}U�lUK��SM�t׉}/9�:�NI�)�eujM���!%ƦơC���wv������?�;��]s�5��������	������xo��rw�Ԋ���*�SȻ��}��m��$B@�j�m֓ʔ%�q'6[�@֣Q8�a?�������^��_���V�
����u�>��L�U˱�s��ؔ184��}�n<�y/��'��"�P.Nb㺕��g�ŗ�G_g�����}���go�����JE�2D���>�����^��_u�u�"t�0~b�}�(N�X�h����hhi������q�]�a��X�ׇk^��xͫ_�|s������n�Ï>�֖֯[�׾��0���w�w��6mނT8����j��m�g��޷��}�NdӍLca�T.�ɒ���2Ƌ!J�� �C:S8��Ue�m+%���ݷl��ɲ@ό0�;׵о�$�(�9h4���c �!E���y��:��T��x�4A��;��!�R~� ��-��L눩rEe�G�t�rr��@*>��%f.;[�J"��ŻqA��[.���F�� �����sp��X{��$�\r��!��Ɔ�2G�Pc%�ܬ�����~��n�_tmܛ6�1�VMu`r��� ��Ը	.;b-�5ۯjނ{/�	��D�1�b�F�ƍ��y�3���}�����꒲�8�#) �@O���tIk%�$9gI!�C�
�N�b��Q8��U3n��}���.n��.kM���m����?��A0~���~��kG�Ө9�_�˜�)�|`tl����w��Aj&��6��j5��N�t�~*a���Щ�r���\�홀�Jw<t�tP!/����TPb�W�<���m���u�.D.���	�u�C���M(����a͹+q��b�4�'w���wl��'01>Ù�\:�,��Sx�K/��~1�-�B�O�\�Fk[�O�ǟ§��6>1�t�iR�G��d�2$"(!(����
o{�0���<��;��_���>9�ŋ�mo}����T&�O�׿�]��'wbaO/^�����K��T&�{؄;~� �=�l&s�?}/���d�>�����p�}�D!�ڷ_�����(��?+���o!�nм5���N�l��f*�r,#l�0	u���䵫:��r�!@iv�(ҋ�o/G���9V܏�Lyt�)�����C���P@��I��
J�Ӽ�
���x��P�&J��eRf�3�����
��B^�ujH���:
1����5��_���u\�/��Y0�|́�¡m�K�c�v�'ѭ{,v��FX�Z ������ndħ�;�"�5�,�4�I��s��Q�9AC�-ɥ����8�C��$cR�t�]���Bs�n��]P��Al�2̹t��V����w��"taR� N�{pb���o��g=�\�Eћh5���8U�N̖�q�6��,nU���M    IDAT���ah�x.�UK�s�t%]7و��֖�O��_�o.���+d�֯��o^�~�E�����t^W��F�.�����z�V
��ٜ^e�P��CoCظ@r��ND�ǭ^Z������*�5�%�#3Xf@�?�%�:��>�^�w�|T�<�����;p�=��ॳ�����_�:r>�	�����}f"�l����~W��ř�a��0�r�,��T�������7q��$�L�C�\r���eFe0�Ż��\��ף1����r��+?��#'h��sݛpᅫ��׎�2��/�|�[hjh����`�U�d
yoٺ�yx�2�.��_|�=X�h>�G�qσ;�߃�zm-y���W�w��J��E��܎[o�
�Fd�$ Lcf��RXA9Jc����d ��Z���M�P	K����E>��$
� �O�F03�
�y�cA_*�F�������� ��S�19>����!��(J&���	��46�p�����4B?�1$�g%��~���^�"�´����p�O�w>�U��ߘ�N�g�5ѳm��s�MOmX���LM����>�ѝ��B��{�+qDnt�yD��Gqn4o����	f)�ю�a�;v��O�����Ѵ�"6P���XL�+a��a1�qr�z��I���Iˡ��
E�Ȩ�M�
mʃt��1��5��KBt�ˌ���Ԇ1.�[�Ng���l�u�u(w7j���%9tܖ�n��礬�({�ބt�]q��#���������3���Ottt���9z2+� zm� ���-Ux� ����z�A�܅r�z*ߎ�BQ����.Y!iXF狧8��>B�Q�R��|d`Ţ^|��w��,h��/�{w�s��?����Q
�]�(����aq��J~��oz��p�W����+�Cc�	��=�]��nރ���me}=zXP��,�t�L�ަo�K��k^�l���Gp��~��ً�#S��lÛ_�b<���X�d��������[�#S!R�F�r��B���MEḩ�x~.\�oxݕ���ľ����/ގG6���#h)d��}	�y�oat����w���X�b��ff�/�{�?��%�Y@�k@�Q���g�?��aQR!�>�f��"�K��t���b��s�^AX�F�!���n�;w���3~�]wchh�RI���d����vd�A g�/�Q��FX,#�/p��B_���R���rg�<V֧�e�x��g���+�I���DTuV�)SQ���=�@��V��T2Y�l��j��І�B�ڇ���~nԿ�N��S�$�ń�v���e��@����0UQ�@"�Q�Q�=��\�s���p67�@>b,�_�c�:9�}�����V�T9������)�/����Krۍ]g|4���IwK8i"d5�	��.��k��"tr7Bw+��l-�΂9ifۚ�u���{]-�3��S��.��r�"�#Z�Ri��S���)���4��O~�/����g�,��C�:�	�~`tl4���$v�ڃw#tw�����B��F駢��[5/�֯D�W�Z�&ɡs񖖣�D�־Ƭ����ڋ"xa�{��]��^��P��`pp���Q�M�06����8v�;����QD!�T"d��.�.ـ�._��\��{��k_��/�e�_���ct&`@��?�L �.��]��iij
�)`�@#���u����m�觿�7�s'�6��]��x����l��u+PhL�?��S�|ˏp`���4�N�e��t6�Y��˚1������lI?�ܱw��a���>91� J���o~���׼ S�FG�1=3���,��r.b���C���_<��I�t#�H�Ԉ-�#�	�qȦ��T@Gw.Y���~�OLbϞ��ࠔR�:��e����ų7^����e{v�ơ�ԧ���S���e�e3�
ȵ�#CLR(NLß�FT�Yh�yY�2�?@� ~��`�9�u�:�"�҂�D�y��OM.=Ԛ�Uq4y��f-1:�b�D��F^�Yӿc<p���H�QN(_�s�L��KJBA��t�Z��8��+�c���	�U��4b�]��1Įu��D�%ޒ6dA�P0n~#���w��w��qe���5��>)�s��1���M|D;���֗��̦�c@g�{��8Nk׸�@�Gg6��b�����!b�Z{o���+�0�%�Հ���QD�ȻG�yss�����������7#@��#5�n`�R+n��_���r��@oA�<_s�����JY�G��%��c�<*����� ����r�Y\y�Ex�e�����@%�\.�|��l6����p	۟<�|?�����t�`�9����
o��*��۶n�=wއ;|/6�^����/�xp�^|����CSHgZ�idH�$�T��������;�/ë_z	���ރ��v~r��
��Z��KV�%W\�Qz���m?�ͷ܁�CӘ.��T��K.܀�_�<\v�|t�XMO��wo��~�86���4��9,]� �}�%x�o=�R������	�w������-(�<l�y���î�tNi���H�)�!u}��ITB�1���V,\��֯ǒe�q��Q<��/�أ�!��rS��/�J���������~�ݗ��151�#�G�ٚ�G@`�� �Ѐ�\�:�\w��P'G�ʢfO�+ş� ���+�M���N6�\�.ѹ� �(#��4$
?�މj�2�Y�������#�J�]��p/�Ũ�ƅҕ��NPr��Kv[貽T$�(N�3�k`�����^{0��T�O� ��3�Сjw��1VvW�W�٨�M�tB��g]�s-֗���j.�Ą�~�Y��;YIi|EԽ�#tn߬ת�f �k� tW�nB7sT�MQ�]�U�C��]@��hx��\�tsw_�=��k#��<��rgʝ�;�0���_~�{���馛�����+�<���0�~ttl �����ڼ��?7�;�N$�����]�'%�:�rg�]"t^���1JS}��w��۔�˫�<)6CpiV�q_�uk����`����exgG����'J������C�ڭ���'��43�g�_��~�b<���
����_�C��p��/ī�~V�7~�G�؋O��á��2M�h������u�h�X��o��2���"����{��݉�v�`b����&���q�e����A��[�s7���;�kp���;���j�"\x�9ذn1��p������4��m?~>�G��c�Uظ~V�\�%p�7?��[C�`��^\��\����������������}�t�K70xF~��"{9r�B��\k#zz{�a�F�\�CG���Cc˦��y
\�p����GWO/.��4��:��}^:����u%)!�� ntb��c@&�*w�ȧ�N"��H>Λ�X0�9j~A� ��҃�r=�D�ll-g�(Q)C���Ǘ�f�@�8\�⤳�U�˷܈1����DGӸ\ILK	��ӫ���4�׾�U�H-��99`J�[P�[>89�8Pu^�Z>�����U�%.���P��V�'�e���X_K̢�T��]�XF]�d�t���{5�SiO�&�%���rw"t��dЉK��WG��sc�U'D�s���ǌ������E�n����
��Sm}��r^��q��
��ǧ����LLL�U����^��?*���c��A���>�Z�������Syݢ%�� ��s�ޣ��S@�<�FSL�k�n�ί�
Y,/�/��hkͣ����=hnkBssm�,�׃e��c��yhj(`dx
���c���1||�x�+pх�����'���㱇7#��X�~#����з�3Q����߹�o�ˍjX�B���d"��Vƒ��}Ë���^ɕZ?��C��{���M01SFOW+^���x�`ú�ܤ�k�ށ/��c�C9$�+�����=]��hDsC�z�ʫ�����yT�CO�ŭ߽w��(�;z��ً֖�Z78xG�BƋ�і��k���,Y<���������O�z�o�P[^ʧsYq�<���q���\@SK3.ظk׬����|b�mނ�!4
hooCcC�ӓ�{��9�E[s+FO��Ο݁���
�2d����-��#�cص�)�P�ZTA�:ؑq��3��,����V���T��݄�������)����M��P��S�� ��@��
+��@]�N�RL��w�Uױ�ݥ�c8��p��`�)���0�U5P(��L�^�_�����D�z\c��%]Ӓ��0��5�܂���t�3��S F����֢'�*��$�-��\o�uđiE��ʈ�u�Z��C��th�^�������Q��Sٚ����q�4c!�D�|N V��&���n��wh1��3ܭe��Zg����#��`�H�B[k˧���?z�����5�{����w�}Vn\P�!�=���*g^K�K�ތ�i�giGt2�noL���Y�:�B#���PCu�Aj�J�^�J��B��,���zkTP�rX�j	.}�z\��+��ف�	�m:�����pp�S��z/�/��b������q�f|�z{�8�o�����89YƖ�����]w?��,Ӫ(����+!�t抸�-/�;��
���G��� n��a�M1�߅�\�<\���X�z	�t��[��/���i���y�L�(��Hq��G1��7\֯?��m({i������[(䚸�\6�G��X"
��L���E,[܍���a�ʅ��ķo�?��#xd���6D�s_yNoD���6�o̡ДCcs6n\���C�سk7�ش��la!M�� ֬=���������݋r�̢��`xd�3�(4��ۇ5k�CWoJ��_�{N�<��!=d�/H�0�@��3�O��>��q>]FV�]Q����.����9S��Ϥ�\�<D�k	w������ͦ�y�yL2����+��z���k\�u�i�㎀��OL8�s'�V�G�D]Š�W8�M��B_�Վy&j���GL��硑��k�r��*hn�����t��=ZD���؁$��m�?����۽s�;�O�L��`_�C�]���^����[������N��W�>'i�j~�}�N��L9|�!8�#��5W����C��_n6�}����IhV��onM���'�پ��F\�����EdOKK����'o:+��U }dtt�աת����q/���c:��z`]+�;�y���H7�(.@����AMcx�}W�#�=^����%2�^�#�����_������~���I�l%�B��U�����,^�� [�<�o�Gسw'�����t%�D\2ETl�ʩhA��3S���4�Je�����_�	RQ^"Z��&L�P��Q\��W��o{-
���I<��v���_��#�0o��{o���������z����n�^xť8o�Z�}l�v<��#����x痧��Ղ?}�;�q�jt�v �����[�����b���h�b��w�oތ��w�ˤ�ؐƹ�,��o�C,[� �O��+߼wܻO�<��׊�BbAb`�~���{���.Ɔ�p���l�ؼ�>� �܅0���+d��Չ��>,\�,DgG�����SOa��xj���ed2�y�͟���>�� �Ã-�چ�
+�d�����ilBKG��%�G�j�yrc�4��z;)cc#L�Ed�� ���C�+ �m����;mm5GO�#e}��k��=� �|%9��+��>e�4*�T�J)M#%v�����t��	��gW�g�F:L���#"��s&,����_����)9�{FǢN����Ӡ�I�����6��.�O�<P8��W�"O�"�C��P���0�N�2 ���R
p4���E(qsM��~�z���r����k1*9Q����^��Ym1M��%u�� ���F����B�����K���<S#)���"nd�G�#�$u�	���J�/D���HݫL����U���I=0s���߈e�:t��չuqD-Rw1C:;�0)�CN��ܥ|�R�R��7&�����ɿ���|b۶��M7��C��[�^�m���qs#gsv�-2��ljA�T�y�%�Ô�׌�q^��Kq�)�e��Z@W4C���nq�(@C>����x��kqޚhjl���<�}{a��(����,�Y>׽�j�`|���7��~pv>���5���@� �,]s�	t�w����y��G&g�c� n�ν�яE&�$�x�C���2ҕ"��i�򷟏k^�b�Z����}G�կ� G�GOO��;/�ҥ����=5�[o�>z���%W���?+V,��CG�ˇ�0� f3���UW]��K�o����I����Oz^x���g_��+bxd�����'wc�8��y]8o�2\v�Ehmk�������&ټG�O!L5"d�{b�eZ\�i�|c�͍�?���>���C894�B:�z�MN������hmi��E��h�tttb��qG���C8�� ��c�hniEk{
�l` �S��(�>�;:X�0M�K��^.���^6��D�Ie���7�FP	oi2�j0�J)w������Ǵ�E�b����՚;�cP�c�ECN`&��LMέ븩uȣ�K=�M����.��J���c�C��t5Rr+.	��T8ѧt>f%�!1m g1�#Dq���b���E�Ǥ��=��̈�v��"���*3
946fP.�p�"�ezľE���@Cc�Bã����K#�� �ϲ�53=%��S�6�#T��M�Tf&+�e��#��a||�����N�C991���^^C��Hgr��b$ϋ�F#a��q�g�����P�3���ܓ���Ma��?���^�.[�Qمt� }*ٚ���U��&mN��v�-ys��I�G��<C��ej��%n�\���"WymE��ӟ�ߟ F&������	֞��������fG��=�~�|�z=ţy].����#�B'�(�0t����'����T�M�G�Z��Z[�8w���{^����qv��v<���ރ���t�c��Ex�E碹�'F'��;7�gw?���������@��Ӿ�a}`���ל��.\��y](�:x��~~����w�i��t�J`RD%�3����p��6�/��ݭ�����܆��I��4��K������'p�w��}>��CG�܍kqՋ���_rr��8��a��̛��p��,��B!�ѱ)�����O��Ν;�+_�4��5����a��(�����0/���+s�����xr���ľC�(��-./�e���82��-�G�1�?����ΰ1�eshki��E�P����cG0|r��I��(z��>��,ƒ���i]�L��Ǳe�f�.��$����z�X�6>9���K��������&�|4vu! cC�JT����I:?�5O�%�	 Q/������������;���k$Kѵ	��|�(�]��zB�}O�sQ��<<!��im��鵥���C��ǽ��fq�X����(N��J��ij�L�2�h����p.b�R�|������yI�(
�;uN��]�R��#��s��),�߉�B~����G�=���`���~��e��yj7\������@GW<���q�|Ų|�S�8~�����B��,���z�#G�q9$1D���CWWFN���mm-�=z�ccX�|5;�����b)@� �)� TS:ֵ2���|���!� K)[W���"?!H�s$�U�e0q�v�#@���-�%c�����~@��K���Z�`&D�"t�,wI��{�U�B>���������_���������Fz藯aQ\��������u��_�G��HSc�B��6"S���zꋌ�q���@7�'�s����z�ex�ek�n� ��!�b�[�R�����P��Χq��>��o`�����PhhV� �L�tn�R
��_����r�\��L�]����%��w%?D�L�dS�    IDAT�S�2@	�bW��$��Fa�����+{�\�01Z�/�M����v���l�w���8zba:��l
W]y^��+�rE7�,�����
�I{h�g�\���	<��>|�?ƾ�(�h�f�+^�W��r�{N;�F���u��C�΁��Q���|�>6�C^(2��$`i�<E�e�H��EhioŅ_��81=�|��==�����.Ө���p�� ¡�#�?zV�B#������Ճ۷c��P.���YW�jeL��,^��k�)r�H���cG�p�� N��s�NyMI]SiԐ'��k&Pa5��8U���)���>�$z�	�N��x����X��}���f '�E�.�2��Mz���L�S#]�-�=�e$0Q�Tc�JK3%:�R�U���R,w�����V�d�40��J�R	WH~\���'����YR�Ǳ62��^~Y"cv�(��V��њ��������[����:���a�����m�C6�����hi/��;��FsS3���OlBSs��z1:Z£�o���	|���b��$���c�����g]���9y�=����бQ��g?ǽ�����U6�G�4�f0S����{�>�Z[�|�jf��؅GzS� �6��xrv��N1SD�dN��d��$� C�6z����J�v0u���˝��ک�k4���hJא�����A����!�����6Y:���=�3¬��Q��u����ǁW��Tʹl�_��������*�t�Mg}.�"���?92�9tt��.�n`>'P�#���nw�g�S�CP�n9t�/-���GKy8C)�Cc�2YnbB����q�b����w���GC.�B>��ڈΔp���FF�ԡ�����qt4@�Fn?+�Qz�������(�)<w�:<�y`��D�
�:�/��8zbH7!

�P�Ñ�ӝԭ�R�9\z�z�\ڃ��m�j�d�����(�lߏǶ��S���%/�|�<��zV�@Gg#G��" 8`f|{��`��!<�m7&�e�r�\���p��˱jE7:�Q�g�ɦ�K�����C�x��'��ݨ��J���VJ�r�aTʈ��(Xh����.y>rM�(�� �@�k��6\�@f�'qt�0��܉�ǎb|�"�4Z[[�zokm�a1D�U*L�R�W2�D��A���G���s]]���ю����u`brãc*:�?ӥ�D�J��Զt��+��H�09Җ<6w��7J5�}DL�J}1��b
_)Y�+�J@2�S$+�-L]�h���FŀJ����ꠘ8:s�.��D+/����&���HN��q��64���VJ���5G/B��!��U(_Z��I��z�%S�5u���@Y�!��e,�߅�~���e�زi'�u�w��҂+#W�v�*N�u�tuu���w�������@�l{r?6mz��x�;���}��a�۰r�J�[������Fgg<�|�������|͚5X��|,\� e��M���!�T����01S}pםwcl�ȃ�x�M�#�*Mx"6G�LĽM��7o��ιduƈ�a&�y7y�j�T�N�A�+!�p��*G*�p�ʭ[��&H�7?�9G��`n�Ύ�3u���Nps��,Pr0�J)b�����k��JU*E/���׿��O\~��a��I�\����74B?5��Cq�J-�^������� �ˀ�n�L��Q�6�`լ
�4/�.�3�I��B�J�B&DwG�wcղE�hm@����2,V���b������w�FK|�{��!k�V�)f�B�K��c�~��Q~-���1<�iƧh�H*!��ڷ��瘺ԩRԪ6("����݆����l�"d�,&����� ���	�[Q
C�&sŕ�9�xQ�:��ԒGKs#�*g�J8>8��''0<YB��q9��<�{��!�����ڌ����J~��"�bb&�_I#�mf���,��������B%@��+�فe眃��N����H�F��Ϯ�v4�s�{)d#�&�m�������ѓ�w��`�|,Z����n�yhjn�~<� ��X.q���� 7��'�@#�n��ē;��c�0:9�����֗�dsc)��\'O�����$~�kg@#�lG�1��`�xX��B�[���H	Ϩ�l 5�<F�f"("�L����xDa+AGr�X\I3�P�Nw�3v����g[ɼ(���|7�=20��9q�/�&Y5-�҉n�*r`��;�~Q�dZ�<�RҰE穀{!pΜ*�8Q�����������-�p�O��hy����1�Y�
K/��-���;������?���y��`��!�ڽ��/��R,]�MM�8|� S꭭m�f3���:�`��/�Iꑰj�*fNOM"�l�x:�]O�CW?;����G���4�(�L��R��tL��� �T��ZR�=�%a�R2~6],,oB��N$��[@���W��i��ߏ*�k���7k7����t�����x��P*+�)���L����)�P���O�����W`.��o����?<2<�(w@�>1@����C���-p ��ZAܙnY=�;��\��^xD���`�:��TM�/���h�l*��"
�K���L}��W�ˀ�b\Vē�����9��(�C�h@�����t1��+�?=B��BC�C>#�u����x����fᥨ:�"�F����3�@tu4�B6�Fr08�����X�b�ьr�� �n����{����$��oxP��5(�|� Q>+�S$R�)POf*9�zo��@D���`���E�NN�5U�HI Ѩ���m_�^>Q�^>�LS3
ͭh���{���J�֫z��
@a�Ap7�&�P$E��K��8^۲��ɤ��tO�33�i'N�q��q��x�,��Z(�J�.q_� �[����6}���"DYdF:gt��#� 
�W���}��߽e�"t����O'�(Q�#1�����.���s8s���9���R�d�r0�ژ&�[p�]wa��e�Ø��«���Ϋ�����_CDRM--hi���H�/�����"lr�}0<>����@ђVb�.g����ł0�(�X��W�Q�Y!���E�Te^c��}�<g�j��v��0�c�W�,��<�SL�29Z���!�u��.������Eh%Ծ���.�k�V�o���w�|=�iG,�avD�O�EyzJ��H���e�R�P��t�x��6����]�x��^O#�$���*|�ER��Ċeͨ��@>��[������>���4b�q�C��CRh���P�4���\�܁hl��w��<���h`T_� ���2EЉ��ttt�c�X�|淵���GX�P(���R).)�\}Ͻ�1���Rd�3��y�8� ��H�xB�~�l��.�
��:(�X)E�bQD ����[�(t�5b�`�C@�Ɛ����(w��E�,V�ݝ�'��]���������w�h�-�S4���?S��K�ΉS"'�������h�7�>��� }����e�R_��bu�4���O��m��;��?@�
��C/G^j��^W�n;��Ώ��Na��|�d���:a�i}���̀'��p棻.����S��hp#̀󜥢B�&&���d�)���!�{q2K�
�2����H�[��&�6��B4����$�B��G�+O �+z�n�t��:��ĝj7�%�dF!�K���r^�-Y������p5��Eä�'#!�r��
]DXz%��²^$�w�Xq𖔠�m�P���T��
/���ϸT�n#���IY�UE_Ozz{0�7���)TUU	�3󼻷%�0,Z��DyY���q��t����EE��j!�ҲR�75aŪ՘N���W��#����{NS:ti���$�P�A&Ma���‐�HD�A�W�o�!�ٳ���a�ktZ��nW�G�#�/ >���7���
*�U�I;]��7���e�csLo�ښݩ�|�?����x1�+��D��Y�b�T�I=��|�L��Ց������f��'����ŉ�\|\�\["$��9��;�Ƞ4d �w��00�;�l:��ߋ��*$Ә��#��i(��L��w7\�����%���V�Quw_�y8��Hy���Qo011���	)X����8�EG�w�В���OcS��D�Q5�*D���o���)F��\P�0����*�.�����׫oE�"��E�D�������f����Z�=C������(�˪c�\@���O���������8���dB<.d���
tc*���i4���&`��cD��Z,6Z�N����9�΀��^xj�IwN`Rb�U� ӫEN/�>}�f�aE�!`n�C��s8�>����ˡ�Mz��� ���E�љ,��֌�3.���������R�I���Μ�;恘wX�K"]�q��\Oq��Ⱁ�h�0�8PS�9gV�oSW�*�(Ͷ�rru@�p��%b,��=�W��
f{<`8Cf���ģ�Q��dR�r�v��#K�jF���8��SE�ĉp�k�$����=�E�4������u;��W����᰼n���rgO�F_?�.]&iqT˾��q�ONʌ|��͢P�aq��t��cp��t��j��^�.��?���Q�،�T��u�#1a=�8/��\�_7�N9��K#k�`��eL�2��U�:*�1��t�9 �uT�gev.6,�LU�b�Qʍ*E���s�\&� $]�q�IK-A�J�L�Y���^���^� c�M�΍�b9ю�(B��>�����r���
�q ��T2��P]���q��1�́�x�u�̕í���Xeg��*�d:x�����{��*�0���2��R����	.�SdPT ��ͽ�/�z��y�,+)�� E��g�Z���E�(���v�dXL+Cx�\��=jώ��������8*�%O�4Fb��O!�=z�>���Z`�b� �̍25��6�aV㌬��)�{趱�W�j��{��P��-�{?H���<VQ�'=�/�b@���S�x^_v�C�����
�hiyNJG@�4���p�_��3���#	�i�����h�{�M��	9s_����?d�]z��
d�;�ʐA�J;BU��I�H����Hgr�%�k�\�\J��8�9sp�<c+x�HЉIu�BbW��e�7 �[R��������%������hD ѩ�y���)%��H��	_�L��*M��	�keRțzI�IF���&��Lc���ϕe�״�=��S��q{�IYH��IN�X��U->���҄%���Ou�ZWb�(����X��m*��'*��u���5+��U���A��9����Ƃ��,	Hc:�~�s�Y�C���B�7�����c�2/引��Co�)B(D|r
#�\������p[}Mm�f?w�گ�Z�tRǉ-� ��k����|&7_+
!3)��q����L�TF^?����ټD�Jih��H"���Uo0�FAUZ�iv�Ȋ��:FI�+�����iJ[a���ρ!?[r�#-��+�>����z�=N�o��һ棵�Q2d����A��4�YE��߼~��D�w\Ņ��1C"I�R�.�����U��ò����觓4yʉ���S�����{�?��P��X ��i \�S&:���� ���+����[�w�u������m������X���������\d�DЮ��ʰ����:0:����8x�N�������������`�P�v8��,tښm�Z��lh6�T���k�wڣ�v��Ÿ኿��^�9:����)+����f���g\�1� �lx��/?x���G�hz��Z4��r/P6Z�X���@7�Ⱥ��rw�*�1�Еy�:�tw�B����b4�ca�͝q�>)�z���(�-܋���4*)qv 2�V�.+t[M/�"�i��).v+���\���"���|��dTE����
0]�R�iM(q	Y��������U��Fk�p�t�����&閹�k�N���x�ڹ�
��.�M1W+t� E(Y~�I���]�b*�(e�$N�JJ�`�JT��#�U��	L��afr��Iy�������d���+��[��f�"��θ����015)�g*��33ؿ{���+��QSY-��Tb��}��m���1��%��8�*�\����j}�?O��y�*W3��}�5�UW�o�, ��&��@c���z��켎�+]HZjA=�
� Ъ�����ך)4#�,�/[���z�[�H�.�l�F'����I\�Ԏ�+��uԎ���U�.��~/�{0�Fy8�G6�e��1E)�y�~�>�����*�{�Y�[�ګ���t�ؽ��ƹ��l�0-��b��>���A�
%�8X���{_Bc]�HSXoNǧ151�Tjn�b��z�� ����J����)�:��c��2+}���!+�4�{�ݘ�����|L�ˤEH�LXb,ÑLe�\
��d�De�!~�������\�tY���0�q���	�kk���߶��/��TG�������֑�H��Y�ׄ�R�֧�q��(�����!�u˘�2c�Ტ�C�] YDٝt1��Am���=�NA�݁�t��+m{�._+E��Â̞��X&e���S��q�q������K�^������b����`=��)^O�#@�E-����m�D��2 Yz�d�
�ء�+�@缓ǩ&���� 8/y�T��5�
��!��I�$�N������ǭvI��Ҙ<�9����\�hY���)˂��Q@^�GG��?ś�O\Bml�.�3K��Ɍ[��<��/D�.�g��sx�`�0��2��M��N�\�5��+<��A�t�e�5���q���9�;�Y�}҈J�/B(��T��t��/9MF��G�(�E-/��O�u��������~��c���z=�dJ'���,^�H����9W�
����rC���Y�]yhP��Ba��]���4��|����q��2�l��u��`��e�Fp��e��ԁ��~�I�����-��|^TEJ��ڂ֖:��F�V�q[�F�d]8}�<N�8���,>�|^,Cit#*`1#Q�3�?�`���
���u�l]���C�j��E�쬔׳$#���c�p��Q5r��T�S��Lgeu�L�P���Fme)�{�s8}����%��X�R��� F,@*����t��H�+���� ���A���_������p�:�G�`Y�#��;(�#�o2٤������߉������/���J���@td��車�<nǏ�D �kׯubd�j��PN]��%¶��FQ�o߾]
޾����׏3�O���j���b��TTT����G&�����&&�P_�Ҳr��_R	����e>��Ԉׯî]��g�^l��(�)����6oEyu���ӎ����7��0�2�&29�3��JDM��B��VE�k3L7�p�cȎ]�ӊ�̓,��_G�E���~�{kzt9k(�[#E�������Y�F��s!��FV��	?��`!E@�D;�qH�~��!�}�_���З�)N�d��[��mp/��������>�傿���e��D��#�,�YR����9����Rc#V��0����NN�%>Ueqg�w���9�G���E	ϝl��U�c�L-鲤p��6]�r4�qq眇<��z	���i9�j�]��婯o-�{X�G�K>.R�\���y�Q*�.�(7�?&&���
K�GM �
f�=ii_���Eͭ��
T��r+S@�������ty� ��BX�Ϗ�fx�a�>|rGPɬ6=Gb<���� �B���5��Aee��6Pj���R���
�s��L%14<�ё���ùS����AEy�z�ZZ.��(:���h�Z�!R]���/����^d���e�9rnN&Ǖ���ew��eK����dr,�Tgn���d�0����u}M5��4��n���G���u�T34&���4�N����$�Y���Y.R*5��h��LX    IDATg�ub2n	[��LT�98�,,��y�h[�*F,���힎Oab|�c�F��aq<���"L%Q	�+_�N?�}�v�$\��Ét6'Խd�s���/7��%��_�>��&��~^�MM��T��k�`��#��'`q��N���T͚��N��9��A3�e*�_����W(��Do�u��4�qÛo���P	**"�Ҏ�a���j��x�snz��o����j���KH$f�6>�{�9���3�K�L$��bc�TD�:o�o��$\Teй"w��q,]�Tv�_zi�a��-���{�{�.�ۻ�7=*l 36<�J+j0�����+ر� �8|i�_�.�kh/]e��5E�X��#�?��Phq������Wv�t5Tzu���U"X��'s6+s�	l��s;��J���x�,���첊�r@$%@>y������c))�m���e���g��?�;�Fܵ|�oe�����dm���US}s5V�-ߖ��ݵ���*%��9+@�!m�`��5H����Φb�9���U�*N����^�4e����Ú@ks������N`lb
�tV�eZ���H�La|,���(*�ję���<��t��u�Kp��y�SI��|�b4A���w!�Em��k�<x�@{�ttt!*AKS�"�u\��do�}c,,L��T�����>��܃C#��O	��{�2��6b��C���ŭ��c��M��E��)XM�ʛK�^3����,��{�ȣB>���m� �s22N���j�%A�|^����%��z�Z�F�1=6��XñQ�����{�^� ��I�-m<Š"�AbfF��]�ŋ���9���k�x�b��׉_6Et���(��QY[���פC��@֠���pgg��+���o�*,Y��Μ�����!������r���s�P����J��ݲ����v��X
�̉�n{�uY�b7�".k����7�S�܌pI�������7��$y�$�qV*d�PQi�]y�T����U���
p����� ���W� :9� ��+��H)~�+_ƙ�`����H@�(��$6���ل���kV�b�]M���ʊ246� ��c`(��]�֏��r�Ӷ=�en�"�+r@��`y[_��/���3t�M��qㆼ�#�(��xM����
\�h�bβҨ���������N�_�@@��_����ŀ~�B�R�鎏�#�
�ϛ7̗3bbr�)�k@���X�l�쫿��Kҥ��O����`�G��`�φ�7 \Q�	��N��{X ��.7|�U5���%{�C�NH�7b3e:Rpfb�1>��u@�1*�]W�"Z��ʆ�b�}���Ŵ�����^�\gw.�X�C�Clf@7?�� [  �i����� # ��Ng�c4����Ћf�r�.q���~O�߳Φ �+��* ��r���;t�C�Ժ��E�JI������3pi�)l޴k�Y�Sg��܅\��'_O�p��{P013E_�u?yw�\���,îp�J��v��W�^���*��O~��hTu�y�SsN��)�|�|�x������G��ҋ{�:�=� �Y�Z�L�;�����ݗq�{ ~�߿[�--xi�19v
]]]b������V�?���pcp^_ 3I���F(^�6c<��l�i�0�/ �����E���(������k�������_QOI	/�{A�8�DBa�z=d-����)��t7011.3���&,\� ���s.^���mA�O��T2���N�?{��r8s���W���q�O���چ&T�5�b�u��t�=��qv�U�,��>'P	a�]�$Fw����5�%nFv��Z�b:T�F&�ku�����Ds=��PQ]�@���eس� v�y�ixڧ2�m���'���Bs�������ci��[�p�?\+QmN�;WG�� ���DA:��KQ]݀u�ס���������a��i"��P)�/?�Ο>��{��эC��.���.����A9��^	�̼����Ҡe� ¥�X�lZ�a`t���6?��AV�v��1�XM�]�<�f��W�����֗� 1gd ����%,�[^?�� zeU��	�]��BQWx�o/�����ـ�uF�Ћ}lT�$�/@�;t:W"�˖.�����g�+� ���S�G����D���<����v����ȵ(
��N~���c�18=1�!���4,8�cȌ\R�.���������i���-p�߳bn3��~�f�}�V�sٲ���LAq� �F1SR�ڞ@������W�!��?r����Ec�u��,�nw��"���܋;��[����Ͻq���������=��!�CM ]CS1�k3=����=�ΥP��G����P[�޽�q��It�`��ؼi5�^ф�+W�\_�p��?|o>�z	�g%~���8z�bј�Aϛ߆t>�y���&��8�v��\o�A��:�x~=�z�~lٴJ���}����Ovc͚5X��ch��Ņsge)���Љ��"�ዟ�8�޻�����3��_܁������3_�֭[�?���ab*�?���!�I��^Xt]��lk�m�N�Z�7���}��ι":4��W�t��F�^����m~�y`��ȼp�����D]E�<.�d���5�_�zE��y��J�BhinFKs#�>��	�i"����TB��(���6���(�����uM�p��:N����k=����T��%��� ֮Z������>vT�K���,,]JPI���P�@5|�A��<n<n:�q��@��
�=�)�M&p��%�={YR���}����hn2���?��|�dr>X�p=+ ݝ��E��e;Bt
F��;��͓��H�d�枵X�x9�8t=ØL�@���5�����/}gN��ۥs�v�7X��xI�;T��>��$q�V�ix���XW^V���$�$�7������g�?y�iV� �u�;t�0�����J������r���g=�d2�:�[ �����ҡ����m�D���Ҍ���'�N�}�Ǥp�c@絕T;�Fr��1���0���"���5@	���ݝ�	й��Vj4��ׂ�f�=��J�ݟf�ewַ��m��������[�c����J&�&�0Ҧӈ�����&`��c� }��ee2_m�jQ�Y1���nՕ��YK��r'�~SUg����m@W��#>�=m�xT�'7�曙��7DF�`IDJ}x�����2�4�b�޳x��1��w����ע�ʃ�����нXy�2��w�K�ǒ%w��'�W^}׺:�k��%���]���o����q1�p�"6�y<+k�ji��}��hm)Cm��5���"�a/6m�"] �����$mpx�^�hl5�|��~%�<R�8�/^�m�_���h�����O�G7�G���(���� .ut�z�R:���C�����B�V�i�m�o5�����{_V)�y�8=n�(h��U4��{�=g
�B� �>�^����n�'&���0��LMM�@���H9���t�U�e������w�!>3���1�imn�3�E:�����;:��2-�q��'�_��n�]FR4��&G:���Om}A��T��(u�`�Խ��$fRL�#�+�?{g��μ���47���B���v���S��yG�5�u� :5��]�j9�n��>�G��¾=��Kg�NM?���ck�Zp�����k�@nb��ErM�ɌD��7��$\���<���L%,X�_O'�b�W���>q�xk֬F�$$�Iگ���NI��T)td0�p;r�rX�d/h�$U�V
�� 6?�o=��w@4�r�̎����}��z�o��_{}?¥%���{`v��%(P�E:�^x�%�������O��=u@���:���Af�o=^��	�<G�[�����������*P�7w�ga�
}ś@Q^J�&[�ҁ�`𐢤� )fͩ�	�V��ˢvW3t-^Uv�z����="P��m��7����,c[�j�V����D:���M���Е��0i��9�p�������t?��� }��ߴR�WGFG��m�o�P���~3���Z�n/��t��������� �vg(o ,$#e��"3ri+NK��C'V�Ռ��Z�5����/��׎������p��AM�4h�?�	<�v��wJdhCc�-_�}��������?�m\�����¥�nL�X��5rn��}�r�P�bAk�$�ŧ����ӟڀm�v�����Ǟ���V��2����pt
/�8���4Z�j�~��q��"�t^�W~�p��Y�����������#x��S�5��Ʈ��ʁ��T8�I��]Ń�F1z�g��7��Š=�	���At���u6��՞���AxKB0�~Q��q��"(���F/���Q���?�x,����q��c1LOO�Fs����P[++j�` A��>r��g�͍0y/���v��e�7+@��ՋS�g]� �`搙�D���'݌��R=.D�!)`(�:}�,zoalrY9��a:�$Ua:��]X�|	�,Y,�xW�5��H�<1���+W��[G1=���>��A-h�s�<*^�}=Q�@)+�W���E�N.'}�D%)��C:iathD|�Ï��$���b��`&I3�4��K��=���������>�U�ML`��8x���;��*i�B�dnj�5�g�����g�r���u���6����#Ǳ��a�e���92�y��C����� )�W_ۇpi��/_�\ tz��r羳M�Е(.)T���>�S�S�:�ﭭ��s�� �M�����6�4a�ڵ����͏�[sܤ(��p��Ul�{o!�S�f�vv�H"P���It��)i���V�K�
i)mf��M"=|�Ԩ �
�����2�D�)�n�
��͔���3����]sq�5{��9��v� G �l/�q��闥�I��vÆ��˾�+�a��=�G��i����F�X��v���x�n�V�Q7w��s;�� ��fI-f��]:�"@/�A�[��Sh���iV���x�z���q<��'���[��kW��Gq��������x��l���V����/����GcK~�?-!'O�����/��������>O&��`i�(���$���<��}�֍�����f�ؾ���e�}`���N�2Ė��r�j��b|"��H)V.m�;oDWW���'F�ʫ�p��9|��G�~����׿��H-V�� ���x��!�}�emJ�q��V�כ�v�-�^��6\j��w�Wء2U���]�q�k��4a�=px}����z��=��3zU�nT���.R��`	��I�n����u\�v�C���C�$�ý��+��,��B%�	����勗P]Y!BCn������ŋ��oBMc+گ����N5C7��XR�(��$�u��Z��{Vb��6�^�������+���Y���^��Ӥ'�Ei��7n�*���0o~Z�!�v�R{�9u��\��tRV��h&���ĲŭX��c�����#�^}�YV�kp,��c?�G��׃��&�8���_�~�	$�^�s������A��ed6�j��4�������`�TF���k�q�T>���y0�����v M#���u4�I��?~QV�֮[+�>�����02�C2��
V��}=��@gh��W��_AuM.]�T�5"�{7�o+t�6��:u
�P��5>1�X,*�@1��r��0;�������.��܈�<� }�~<��1XVV:g�J7蜡���^��0�f$��iRt�lt�}as�q���2#JGc�,uǊy#��r܀��CR`��[qU�о߹mㅈ۴N��U4��v�t���R����6��߯����7���Jutt���^<�(���~�����o���h�zfI� z"O�,Eq��D����s��\]|�� �PE>0���H�E�*��W�}����x�����1�<}N3���j,_֊5�ZE��}} �^:&9������z�\�##X���w���h?R�B�;�a�ĥ�=��}�1<��&tv\A:5�H���-ā�������0O vfj
��x��Mr0~����c~[�d�w]mG46�-�l��⋗���K���c�������&��X�~#�Zڰ��عk?@J��,i�¸D��M^�N��|t����"�}u���s�^'+�.�8�Q��U63�����?2�����y����P
���AY0��DldёaĢÈ�F1>����0����(��mHN��y�U�/nn���p���I\l�@u]�[q�zε_U*w�P�ۜ�S���,�o����fy|1��A#�i+K��*v���ᐙ��+N�,vu�t.��d7F008�h,.��C �UQ���˗�G[[��PZ�:W�f��m�S���"�T���h�ׂ�i���*K0M���(�v�b">�뗚&u{���*Ǣ��X0/��߃����I47�!e�1�F�cK�����z��/^�b���.ut�ҕL[NX9Su���C�����`ߠ�+2`g���(+'�W�
�^SC@���I�(�+f������s},�T�����B�~+@o[� ۶o�⌀�a�:����ُǶ~��A¢(n� ��)w�+4�.����ϣ����O�]�#�gRbP���4�:��h�����Pw��޳�_���r׶
:3B���b�����m1�K�/����'��?���U�Tŋ�_�����SL� ��#ס�X��7�)뫣�Y@�5.�V`�������{���~JK��x�g>X�R��z��:tQ�Dq
���}��!{)Z�5���,;�4�7��?�[6����x���:sg6R�~7�	\�܎ӧ.�r{��q�z�?��Z�p�� ���
^}���$���dv�4m��>�������afzJV��jK�dq)�=��_{N�%%%�yܘ��UK$!�Ͽ���b����ލ��qd��?"���j����6m^������#�Ě�֢�����:v����ä�-���hel���!��Ew�6����
{�3e�S�y��tֳ��0{׏CM�i������.)�YB��%�aT>;�u���P_Y��p)�>\��Owb�׺08؏�񘴊�5ܽb9JC%��nf���Q����A���DBm�]�QUۈ��ft���bG�ˤ3�u�+���kB���a�Ө.c��u�:1>�}��cxtV.� ]��s���2瞹<�|�cX�z��gϝ��g1�HJ> is�'�,��i�w��p604"�7�W�{�⥻���>��i���7�x��;���Ӑ�f�L����8~섬7N',8��&��|�����g�e�	�h�<4�U���W;��` �?X��n���)+1gss3FG���-� �s-�Z��N�\��<��[�܇	�=}콁HY����@/EMm5.^�X�Յ���.��I�����҉�������#���I�;�>�;�%�r'���)4����wz��6�Dw�E�>K���|Е6őIiV���!\��=��b����wX03���܎T��,)bW�v��UFS�2��])o�s�b��V�Y,�Va+�&ef���qmM|��}}�?�;�PЭ�F���Wf�E�~��A9������ ��<��������O�]��� Ew�2J���$�ſg����w~�SX��eA$��;?����a�9,YZ�%wՈaHr&���1��F�>q#��X�a�l]���J��_����և���p2A2���pd�r&�:�Zv���w/_�G���[o������b�������ue�N���?�U�Wbْ��￈��~Y�r�&��޵ ���ߋ���+�����ݵ5�8q�4�;��;�2��v���������{�^US���    IDAT�`��.*cYmިo`c� ]������Y:U5�����8˲���-.p��(��|yI	j#�G*4M�x�Z&'b������u�=�*Q$��.�;�
F�66�Sg��hlݽ�(��FYE5���i�B�neLt$e��%a:�𙆬f��TRv�)�b.NFx�~����'IQ&w�9�gVy|&��f��h��x�"����F6��?��������E׳�D���*]��9�� ��%Ia�F�P�+]��bI�m,��b�$kDfq�<���z���w�<�hV֡F'.S�ҕK�2�a�	W
�si�I�4)�\T�}m\��[�����0z�pC��cb�]�u5�p�BЫ��PYY)��� ���9�8y�$J��ʝ��s;���F�����G�d�Z[{y�$����� �6lڈP����������:x�s(�q�}w��7h��3�10��Q�M<���IdF(����bZ��|�i@72�f���V�����[5W����͝��w�r.��ж4���j���=t�s-��5�p���'�kW����e}5�Ѕr/�V�+�b`�]�}��]����SR�6�ϊ�f������֎�a��� �\�����2T��T��ÅѨ%9#���2�d�yCv�;����s���+E[[�JKp�dn�cr:���R������iFR<�I�rE���u5UX�Z���\�rUB^��Z���Yv���&%�xP(�HYgO_��D\���kkFUM�.��C���.v�"���4fō���挘�JLS��Ee��%�Uf<�d�U�- �3a(��x���`��Q�=�ˌG�ٙ�%���ϟD�A�W"������iR	��yV��J|>�������nI<�ON`�ƀ�U�t��Kz���gϞAii)��8㍍O��o .�_>z��0:6��tB=7�85��@����e/L��X��:�u͚R�)�eCOS�h�j�Ƴ�b��l0�X]�&���QoSv�R�RE�U>�bIӘT���g�)P���~�X���^ڭSv���Y�Q�T�D(@��'N��;@:]19,<x�;J���D�ʽ{���^S�J}3�X /Kb#,7�V������H�yx��}��3 � �ޝ(�������
WQQ	��f@߶�eYO���t�;~��xy�NY�khl���w��c�>	+�F"u'��^3Fƒ!)	��g�2q����(W0�=�k�rXpeƑ�N�:�kV�s�h'n�c"���?�pu����=�^��ܮ}����J��2�)g�5Z�:�XF�Sa܅:�|s��p�e_����A�����t���L��_�F�5C�� }n�~���g�6�#wH��y&XќC���+ݡ�x �i��s�F��x��t`2_�3�-�$��s4�$�ҋX��[��%]̒Ǣ��Ë��F��lz�e�ޔ��M�����Fp�r�$�b�b��g�p/Z�:y�9�5�w9d6���'(�o8MٻN�g�	�Ě��nwPv�)��� vU&s��|Tg�B�	�Qz�XF��s�⨚k~#�^��<Tvd|�fT:�-�榁�^��.�FI�NP��
x�_��.�Gv�9��nl�,����P]��@'a�	e�B�0���Fʲp��9�B!P�O�L�01G�� R���?v���^2�a����W�Ny!�Av�mɠ�0E����4EܔN�����ʚX����!ׇ#	1�U�g�y���*ŏ�+U�t��A(��*o�@g�����cfT���'y��A��>�ZF76�Χr�m�w�0��Q�$�)�x�O������͢�բ���%\��p��d@��9\Jt��D�0����u�@�;t�{��D���^����K�>�r��CW�2�ضm�M��O��[ZZnR�s����,\�m;v�𭡡7n��g�~|��'��=����I�'�#�\��}�q�֯Z�(w�!��ra���0w�S�i��a&E��)2)�i8S1`�j��^��2+��=��ӗ_'P��Z w�B����d�l@��_�w�y�T��p��;:y��q8��}}���p����GЗ��@�����X�eYB��4
�?���t���U�O����ڷӽ�H8��Pw�^@�֯RW���D{�R'q�{E�8U�|N�mg��������sx��K��l+M�p��]����p�{���*}�MF�|uvX&�Q��������[���*�-Cs���MI8W�\,$h.A�w�dsj�̵!9��H��]&s�U���Eݽȁ�3sz���seІ�o4z��r�ςT��6����dZu�seIM�Ց�ʨY@W�6�I�R��b@��{��֮a"�R�.�p�����~��p��9���l�P."��`NV��C�gc �TW������;��'����ffH[����+u��n�z��B�Y;u�=�ZNS��s���ڐz�$��P`."6�5@�=�4����"H���������;��� �����*�L{��SO�Wy�����(,��De���Ww�N���[����P�hAA5#��*����Q��p,���U�O��;rp��V�?��g1�a�)ndh�ʝ������2����̙3�;����Fv���n�UWWc��"�$���_�mR�e���Xfb�ܙ�G@�����Ώ��&q(<z�8�-X�۶o�.������
П�����t"�6�CYu����s/�=���րN�8]D�	xO�C�{�|�ϝ��`l*���&�f�fJvH��1v��X�JQIvLއꞰg��ښ�.��n7r6��;������m��;_��yM��cn�-�#~��27��Y��4xt�\�������+�V=��T�wcccMt{~nw�ŀ~������������c�6���o��tF��֪�6*?	?X�ы���y�C�+0�ָ(��r�1LX9C�.�kgX��u�Ŵ�׈�d"��9Kf�n��t��G*�2ù�4=FQ�,2��%���LmޑGIЏ%+cx�z�]�W�'��I��V_�-K�-M�'���TJ�^��n�NӐ�^���߹��	���x(Р�iW�5P�Z��Ի.����*dlʝ�U6H�u5n�I��yf`*���Հ�.��D�*�z�&Wֿ\t�3�����p卫m
�h���z��p{dN�q�%͍�(���s��ۍ U�	���(��Ie�����*�@�<�B"M�{mg5�K��� ��PQ���eǰj�"�`���(�W�+�k
z�a�k��8ΐ�,��Lj3�aOPx]%$C)�eUI��j����T�kk�2#S�
	'�z�A�D���>6�z���@���CJ/3znz���==��3�em|���<Z�f���-���Z����=;
z1�3��t���y6���f@?��Ҳw:}�b�N0�0��F@?r��-[����%��iӃع}7��ڏ'>�,n=$�X��:�V�b*��av�{���C�HP��W�-�#a?6<�Z��ɩ8�nD�?8�hlB�@R��,)�+0�)N��d�%3t���ʽ`��sK1~��Ă�(8�>���b���[A��e�
6��=6�Ɖ�%��q��U�l8)����p�z{;��;����?����S���{�V/�{��v��:$r\c����� �f���R����ʍ�t/�٦�(13����L�\����&���rb��� �	=�I������4�%^1B)����a��4�&f0����7����D2�Ao�$�'�%Ud��d'�x��P�'?�8�_8��G���L�a��R��:@sY�����\Q�,h���144��pU�����Ob݆{�h�b��?�FG� &�H�3C�Pip"��{�`��O�KW`�R�bB���3rJ8�(zա
�JJ�^Pր.��"�I9`(����i؀�q�!��v��7���`z���T�(CA���������d��U�!Ѫt��1�[+pvw��_���d)�Bg��J_!]l��2)|��%]Vmr^}�ʻ�3�ya4�-3eVn*TC7:2G�CS�,<IT����_Z��XFT�d](`ˈ͠O;y[*Y�Jh�^wNtA#�~�=�ʲ��W��t�c��a.d�����q!�,��^׳Y��T1E��=I��f2�ա�7�w蕑����Q�)w:�)/�t!�������v��C�)�b�ܻ���ݡ�E���M���g{�ۀ~���E�/�N�M���Sr�g	�{hJ+k0��Ӆ���M�����D'�6G9�4"eA<�e~/�'&�y} ��y�Ƥ�p�9���_�;��h�j��@ȥ�:�E�ˮ�t�vдY׹3r!�v����s� ͎\��v{��)-��i���A�-���ء{=f��0������ �NJ�e�6�z:m�n,k~���=n1Uo��sm�{����i,Cʝ6���*� �)@:��QY��=�	m͕(9�+q�R�;~'N]�}�<��m�3��	
I�y�G��Dtl?��0��	�?^����x��9Q���U�g�[���0�{���ݎ��q��$}γ�+;HO��ի���{�q��YDG��7�1�N?�R�ӉƢxᥟ`������������}oc^S#�ϛ'��=�c�]� 6my��'Ί���y���s_�k���dX�t�PTia�.��b�^��r��֒��.��jC��H���A]2���̶�Uj)Гn݅��:�w*~m�5L��z��4�R�q�� >�4�crI9����X�Y9�N�o;��w-��1���(���j���}��ke6�1��h?�ܨ���4<���Jxz�n(�d�lVU�x�¦�MbbrF�ʥ�Ub9�c��d��_N�Y,�h��V�*���AG
F�|�|���<�@��dZ�Yc�qY�R4<��\���n�F=�x����.3{�rw؀^�?����Vԡ�)���ZeE|^7v�#T���>9��
��X������W(��*E���v�n��rg 3љ����^Q�#B�/Ţŋ����*Z�P��o�}��}x��O�O��`���(��Ŵ�( �����)��T����>'֬Z"l	M�2Y�G�0v���8rQ���=t�pl�2vR�n�ikB�(a�};�������@�V��<ܵ��a�� %�-M��3����h�]q�NG����:��ovu]�֝�����}���5�"�G[�=�^�sA��t��C����a��gЇ�е�p���CA�����	|�*K�ѽ����0-o�����p��-��נ��:��0����o<�k�;�[���#1t]����-�e9�7}�7*+��{�`��E�o���T��;{q��5����H�I�ǧ?�ٺ��i���p�)����yDG�p�h;FF�0�HI�}��|���g���9�w��G�J���YR̾�O������a�&�JC����}�0\�OrХT=+S�E`Ut{�O�K'��v���.�[a�Mg��l�/�|��AKB����]���b����
H��".�S�E�`u{$^6�L���YdSi�0��X����X��N�i1���C:���]�������~+0�멩��//ÓY�a���ي^#��T�����y>76�z��������-G"������.^���J�)��S�iap~�XY��T@Kał��w����Sk��ۚ��T�Hy��)����.��_v��v��U��O��X����XȞ�r>�y��~g
��i@�]S�"��{�4bQ�s�B�N@�;�H�� �}}�7u��I�?��32C?q�J�t��@G��qաs^�N�����.� �!,[Nʝ�	ۥ���ÖMa�]ؽs�|�i�Ri�\�HM�3����:�d�ny�r\8k�*��4֖���uA�20��8���㕄;G2
�u
�NêB1-�9��-�й�8���;�:2{��\���z/P�K��kk�A�P��[<�W�2J��"��4�>���p���:�w4H���}D=�;�h������-��{!n泇��Q��|p��0CWz���U:)wӕə�t�l��;OR�� �7�|~=��]HL�����eK�f����>y�"U�~�H`A򝓧p�����_���{��ێ�y�������445�����I���%�kǛ����ū0܌D�j=#ï��'��oķ��]��PW��/�����A��FllR��g��4>�O�����f0��̉S���A ¿��'p�J�j�j|����}����	�`�puM-')p��lPD���� dwY�fig[�(W^S�b�S�X׳�xύEK�]�2-t���mi9�ƪK/<o�R~<H��|8Ҝ��ma
�c#�l]mZ[3*>'q��3����A�`e嫂[�6G��
��!i��_������S�{J}����#���n\������X�BL�m�L|�[�����`������5㍷���ނ��U:��R�NhJ<M?K]�9�H��g5�pf���Qp���ܻ�7�4�E��� >5�/���ZTW� ����s8x�nD�œ��K���x9}oqK@�Cn�����������}��_�֪++з�x�0C�������x}>�����N�W������bbE@ggϳ��Q(Gv���9Cy�v�4 �o��0vl�%�'� �zyu-�i������������Is��QO��+3,��(�5��a#(���ψ�[�|Ѐ>�rW� ��еS��g5�V��� ݶj��t���ۀ^��L�ҳ��]?_���=�*��t$�^O�a��u��w���~}㯦���D�Q��E�JW|���ߎ�����ߙ(n.��r����݀n�����l)pӝ�a:ᤊI�3ؼq5�� �C�r�¡�0=�A}m-~�sObْz8]i�{������O}{v���Ͽ���/ţ�nE]C=����s,[�ڀ�'�B}}�/X��)��z���6�D�G���Ώᗟ{����׿��b�����}e%AL��e��ͷNaﾣ�����$>��G�������4�a��=(G$��{��7�����ݍ/}�)�y�0��O;�f�h��Ճl^Y���Vy鎽 �Ҁnw��.�i�Ͷ�g>E'ˣu�k��YJ�]��AV�4��bV����Fv{�M�9�e����;Q�ZeΚ��"����3�4#{�2�)��]���m3�qά�{X��������X��|��]DI��R2ba�����hF9�RdF��h�����>��Kbp�]W�05ǽ����'���7�p���pʺ���u�E�p^�v-g��0T(	W.��7܏׮���:.�C��k����?c�Q�H����(H{`�*�.l�������vt� g�UqCF��)�kc������/:t3)wҹ��i,C@��x���r��1m�ō �xL�46
���� :i��[Q;�O>�:���6n~�Hb��<v�^=�C��!a��憷��z�[p:��G0�����)$-j!h�`�c�d;'9xNKS�Zp�"�_�����+�Fj7C{�=��w���k�!~+��ȇ[D��*
�!�%m(���[B�]�=d�}�].㯯^=��?h�����Hz�J���@�_$[�>�"S2�{�>��*w���	�R��C�ۡ��Iu��Y%���I��A�zZ }Œ���"�Ϋ@.�@w����똜H�����`ѢzTT�`p4���`*>�/|������O�a��ؼ�a����O��ҝ?��&���u�J�1�"�G"xiǛ���3�҅:�4ܹq��W>�-[��|������j���Y�)\�p��Q\�|.^Ǎ���KO�Oo�w��ee,^4S��~����7ٙ_�j���Sؽ� ��O�šJ���9v�*+Y���|�+��,�mw�jVW�C�oO͙�b:5%/:@
0��-�Q�z����v�R���X�^S�.�)��>�%�H&+�;{Z��E+�-H�
���ja�    IDAT�L:���3z�L��
�UW��
�3[�(3�µ�Y���}�5سK��b̮LF`�Uƹ�B�(LjJ�n�Z���[��x��݈O%p�ڍ8u��<tNOP�`,�/��O�֊ I���R�����I&�[}7j+�����I%1������ÎE���������x�{|�>�F��?��]=��!e����v�p垃�i�V�����zPSU%B�m/�P�Ћ��4,�N�[�M�s�.�^R*� �o
��@�;tR���m�ݞ��C���e����M�C߹O?�)}�	p�CPVU�)�ikװm�[8��E4�.F<��Pt��i��a*��jj����B�/\��T<%�)�r�O5�c�R�.3��V�3�ZR� gc��!���4�]l6%~;�^|�w���,e����ܦ����t����r��ի���v������&����0:::�������mP�������/{��u����g0�D# $H �{��)�QŲK�$�$N�8��ܴg;��K�/�_��I|��KT�D�IQ$XA$���O�yo���9��b���B���̙S�^�*��������v�C�:����E�US��J5t���hL���Jq�%�E��E�h�<,_�>o��o��ٹ�3�12؅9�EX�t!�/��w����o��Wq��q���~�]����K�3/<�;��Ķm��kG�9X�b��r�}�����%�J��X�����������܎�����W>���6�{�45^A0Hқ	��'������?x�7��Bl߶�Hg���߾�S8\iX�j%��v���{��O_�4,:1���R���b���V�z�� ��U�q;���\-G����#У.��RD��� tK)@0�P!R�z�$�"Lpa|���R|㱺*�g�Fd1J���TDc�]�X�"~����9�Dͨ�r��~"��jf�ڹ���&�s�N0�۝��S*o<̂"iz_�xPX�6</��r2�p�][�q��������imK��Aݥ&;Y��̓`,�]��)����<�����@��a #͉�s���{��֊��!==�%��������p��C(+���%3�?#�h��g�r�������b��y@e�ԕ�G�n�~����}x��>������0X�0����E��ԇ��܌5*B�D022�)�,�Ď'�E`>ЅWYU��{_���(f���wѴD���G�w7o@^�غPS��3�?<U�-;�Ag� �����aG��vs5�"t�ǉ���QR\�����5��a@'����">�	�p˸�r�}�KT ���=*�(l�����g�(;��m�i��$;��5�:�ٵ�������X&[���j�̕�n�}�F�������tS����k���c�Э �
̓���z��m-A,wt���L$��U�D"'�&A}��ސ��C���bQU~㳛1�7��+�7w6f�,��x����X��[�����y�4MV���x�������;�yvwvbi�������x�JKx�ʁ}�04H)�|�yh7��ub�����gxZ����x�S{�{�v���._���4��ǐ������p������7�u�Jlݶ�=w'O�la���=�''N4����O(�U��[w`~y�x� ^z�8���ȜZ����7�Ur/�%ʔ^h���)@g���q���9�U���Bsɨ�ۙ-/���?�c6:B���x�G�R"���w���J��KRF��\P�_&�)\���+҃͢��j׍�R�fu b��{<!�����`��Amz�{�@<"�t-.�m�IYW���8��
r3�'EwG.�����@�f�)��X�:z��څ�`��4/י#��㘐E� "R�ĜvE��y�j�[�����zp���{04de=��S�e=WW <>���v�cX�t1�Ν�w���E�V`^�B|�?Cg�0l.J/S�!��>�����QzK�
�_x�Y���@ɬb?~���|m���I���)�n
˄�&�i@'G�R�T>`@�GVV����J��R��+@_� {_{�##<���;�����<�:�׷�܌����3-x��q��kB��U��\m�닰�$�p�0�32��]<m���G��Aw� w��
�8�<􋰇z�L�Ô��G���(�(UZo� �^�ﱂ���n����T�T)|�n)G:�Μ�t+�n����/_>�_��`���[~U�|���SRuzV@OV���t��c��I).�&ү�%����Ѝ�<el9"�^Q�b	L�&C��cǬ�x`�R�9�"���@`<���;q*K�bE%F�B�OI��=}�8VS��k��y��#��C�߇��p��5�)�����X �uW0:<z:�o\�䤦km8]{	�����xۖ�H'Ǐ�@�<�g�3�P�G���c�<���+��ĉf\�܌p4���� �׏��^|�=�q�l۾���q��I�>{vR���Z'��X&�)���gn��zȃ1�D��5NQ�P�R�Е�-���<��h��o���痕�!K��j6=sE�c�(�e���@Z_�N�������RGW�5#RQD8nˋ�+�r�4g�`��+GSz��z�*@��z���9�-�M{�ڑ����Y�t��"�J�`Ú%��Dg[�ry��������`�}���,���z��N�,�����Aٮ(�{֬\�_y��d��Ļ������H�Y�	:�L?v�މ��K8]s�h�V�������ى��lx|�8][�+-���2O�2��Y�$y�R�J)n>��� ��
)���E3��O��/>���LH�9~Lz~;�~� �V�{��W8�nzг��ё�� ]G�V@?r�0-Z��{_%@�ow3���5�O<�IΤ����kn���8v�o�|���\�Cca��u���JT�G�:_23Ұq�
dge`l<�ӧ��;0� �׍'�qD�N�"�C��ǀ.ѹN���8���J]%Өԗ
�y�Zu%�ʭ�0��5����ʩ ���|7	���[ =���vٿSWw�_o�>��ގ)�_�D¿���;?�)w�B�j$��\��L�i�G�"|��O*P�z�S=zo�X�� ��M\��
нb�uʇ�Mf���9)RK�&x b�=�م�(-�Ea^�������!q�a���9�J�q�M�����7JKg�����A\�����ee���G5��KAR��(�u�ñ:z0>D"��nG��YX��
����c�ۇPZTy��0�h��x[G?|iY�gs���8O���ʀ�MF!�Pp�޻�Gn��?>���VeIic����0ɉ0C�,�s(����QN������U��Y�l2�V���
ᔮ���]#Z��1D���P:SѸ���?���='���*(�x�j��%�Y�M>IJj�P�.+�ܪ�x�����u��.����mXUK���OS,ked�X g�Y
�*�iv����d��h L"���t��c��b��0>:
�;�Xx�p ^��Ò|1��Rz��E(�73�=�#��؂��ǥG����v&�9(�M�][ףr�\��'?C���=�
Ͽ��C��y�8b�Y��Ǟ�4jϜ���^g���%3�t�lݲ--Wq�Rf͚�3��p�D-�.?b4��	�Lq�G ��JqԶ��Kry�(-�ޞn���U\Dl�t<�<z.JJ�q���z{�mΗ&�.z��C/�+����䓟�;:E䔪�H|pp �())Ay9�܁�Q�~żye��/��C$,C�� {����!�,,������W�
�?�(���[�`a�� PS{��;�����X���A���<����I>����� ��1qv��eb�!�"C@�8��*�F�s	+�S	i��p���Ab��֔��^�J�'/l]#פ8RĔ��ɽ�=�]pN�}<+#��������j�m*L������_��#_���+'@7��*!ʅ�-�L(�2er����D��@}�0��C��{q�ÕYWzƣ~�@�`�LS�n �b�FD�n�x�d���e�a�y�8e&3-JVeR��͵M�I��(��q���_��	b ���u����a-/��^O�It��D���Tr�R���������L��Ӽn2`�D#a�"d�IG�°;ܼ�	�D��@J�Vh���Ì�t�}^tu�BQ'�Z�x�+��$	Kuu��J�0I���G��'Պ�4d����5(Q	"h0�������7{�qT!��M��:�ovH�d4�z O$Mx��lL�p�B+�Rk��'	e���HTr�����b:$�7��'@�,7���~`2���&��\�f[�D�!�9����$r�f��	�y�ȝ���U%���mĹ�+x�DBc�GB2 G+�����)�O��l.6o_��2�󿾄+�휶��I�8 �
03�n��*CI~6Ҽ���P�������FÛ�Aqq!�mی����Cp�ƭ&0oN!~�w��p�x-���0�;\�^ypg"��"Fk���j\k"�=���r�_{
�ra'5G��с��F\mkE��������?y���3{N�|��R���/(�a<�](+�����{��-#��'�|
������ə�X,�u���~&��0���j^oԟ>88���J���a�jTW/��/��N@aA��.t���#��{LCU�غY�� 
A͙f�u�(j�\BaI���q���=r.��� ���\X�r��s9�:w�:::1<:�Ι-�=�[#���K:]�;I��5)�	�>�i}�â���穀�M�?�$bD�����-p<`H9������ٙ���SY�� =�徾���N�������DEn��/����Α�����Z8B��q�Ý1��"�~D���n�Q�CL
�~L��!��A�TɈ�U�7������B<N$����+$���zE������i�vq�PB���~$�J�8ENnI�1pq�$HC��*	ٺ]��KbÃ#���ty[�&*n1��H)�>��+�/j���éR���ԃ��ش�3r�K󣳣Q���|f�$G�I�;���HbҮ"[Iˢ<~S�|����x�06B$J� ��9�t�4B�2	���m^*�frE��T)qJ��B�]2�9R�|(ZT�p��]"j�ҟד�8��*/6�ɩ%M�P+R���sW�"���z���2q9��^��� Ȁ������"�9��H��������p���{�TU���Z���)-�6:<���TUUp-�����p�,]���ݟ���W��r�E�g;1��{�ay5|�	afQ>�ǃhi�������f�E�!���EeU��<�t�.�]�����(�KǗ����\F��<��/��x�}����y$�"0��Ģ���מ@��<�h���nG��&447�x�,dd���g^B~n>f������0������q#/���m}���SN�h���*cuu5�x�	466q�N}�\Ce�N��Q\\���*���Ap�� ���w�l�b,ZT�^؋�a��{��+/���2>�(sFAܹer�gb<lñ��xm�a�<[��+��;���6B��r�rpb��(.�F��́Cw� ��\gs�\� �~�� ��rW�!>Jw	�=&����;N��N/MUV����d��]^O\��|���b�@��Kn��Ν�����k�g�wg>�o��À���{Ԉ��t
������D%&$]����\M����;���,��_�`,1�#N�N�A3����K�Х�*"Ru1k�"Y;<���wsڎ�Y�`���յ�8k	<$x���Z'����X������r���LN�D���H�	p�8E�"~B��� � ��r�����#��aD#�p@Qn�ٸ�������S��iL��Y�����e����p����D�X*��x��� M w#�#2���F,�2���ِ����7��h�#���0�(Ba}};F��x\&4�.�Y�8����Z�Nd�2�9y���$`#���E��tI���Ƃ!x�vd�I�'N���(J0ًƮ����s�0�Вm�'�Ex�Z��#���u��j�T���ݛ(�:�Tʟ����&���'��QMR㱿���B�||�m�R_�˗���������<�{����BhkmEWW7|h7֬Y��}��P2��,�˯����Q��G@�y�Ģ�����z>�1D#�XP5C#�h�ځ��D�C� V�^������Ԉ斫����!iy۹k���ۋ-�w�ܹ�8t�	���Q�z(�Q�L�=��e3�ͯ>��Rt�C��׍����k����9��+�޽o!F>Jf�D��cth@�݁��\ddfbhx�EE�]y{���hS�~�}������_�?-����)�������̝[�H�dm��w�Ki|j.G�UU��(��w�9ȑ}AAv�،�－��`ǎ�02�E蛷"�����h�˯���zܹ�.t��\]#����De/Z;�)��Qn
0b!��I8݈Q�T���AtWdnb���'H�.�˔�d��_�'+��Q�n���9'��Z��}�\Be)cE�����>>#;���r�cm�ߟ&ܪ��v��t՝�G~����<��L����aM``S5�K=v�bz�'�,��_�Nj�n�m
�3���#n�#a����yjMq���R[�����XܮC�	��v���cQu��K��s��\�k��@��-Y9~ܷg��Gp��\��@(ǌ��|�z��E<A��shh�µ;[����T��b.��q�lzcG(|�el���!�ڱkV��{��`��2����^�E���ý�gΞa�m_��g�����X0��.�P�Yآ�|���]8C�%з��o��?���r�^�=��x��|p�Q7�L�r��I��xe��d�|����� ^�����:QSS��ￃ��[6o�w��
��;&'>*}�|�>�^^[�X qv�h3{$ʦlF4(cl�D>$\$�Aҥ�	1I�e�!;Ӈ��b|�s����ĉ.<�����ѡ�5E#�`s�dD�{���7����Ip*�V0l4��Ϭo`�f�B�3=]���$XoC�;��Ѩ�n�t�lH�:���E�߃ܜLTVV�|�Y���aúu\������V<���X�q-��W�Co�8ܾt&UQ�����F�'�J<��Z�l�����!DC����2ς��h�� ��#;Ǐ��4frS�8�*f$�C\��De�gK��L1���Y����M�נ�O<�-��$��UI���A��F02L�]��x�U�W^���� '+E��nkA4 ɚ��p{}�l���s=����ϝg>�������A!}�0�̙;�?Ǥ3���d�p���&G)}��eYSi���%K������X�h.�7����7nDAq;1�/��jN��~�� :�۩� �ǧz�|I5�� �Xձgp��;�p;i�3���s��;2t)I:�C)��<������j�Su9Y��(��q{��;w��,�w
@˛�W��x�{�ԡ�*���qo?@_���P��=����H2�K�[L���R�ZHc��>9n"�{����2�EL���H	�+FB:'����cN]*ږ�	'�,J��aϽ�8���%��������3�y�J�XU���k8r�4�}X��|"�-ł�2�D,@ZZG����Ʊf�V�+�(�V���/��cx�̪�f%�G���u��۰�j��{?�\,_��9����a�]��b�;w���`p�n�jlܰ���/64�{?z�ݘ;� _���"/����8}��c1��b�khF�YX�zV-��>��/@�p��{NsD:/���_�U�`��jI�650�gg��ճ��{�ߎ����o��g���GF�s�
����ѿX׊��A�H+�!� �e<��Ch�҄��.,_T���\�4�;Q�Њ�-ה�%��d��93�zy�ٱ9ٹ����    IDATvm��γ��6�o�BP����3�����!�bkKC�
�u�=�Gj���8]�kf��u��R2d�L�A'0��$�@�8��K�戇0n	�����t����]X�f�,���p��	wݽ�7�Ǐ�"���P�����@c�	�KL켋F�=D^�9�^���#	��뢪%adxs��DwO���p�y~��.����&��3�����mW�K�������t�_���\t��G�<�=�E�s�}�r�1�׋�k��P�y��*.Dłj�:q���4:wl�y�3xlj�����02�z��"�h��9)��(w�w0�Q�����NR���,6Cuuj������!��ds�:��i�*
�t��:�������	��X�zf���(�����T�%�\�	=���o����qD�j� ���#�r_�fO�#����]��d'�e��F���#txj�C:-~���z�Ŷ8Թ^�i��L�K���6r�	�isj����Q��g���u�8R�Wp��v�ˉ��t:�{��s���՛?
G���C�!]F�C��,.#s�ʄT��)�i�(�=�I�j]K�`�?C�����ܶ��"�71��[at˴fh�:�iL]g�5m�@bDSt<�8��w�&:]�،�ys0���p���Ŧ;����AQq���c߾�8�N6n��w߅��Qtt�"Ã����?�O~�:�صk7�7���Q\�ҍ����E2��Xg�R�n�^]��#+#����kp�}����	'O�����7����O�B`|�vm��w��,Dvn��C�����eag��o��e���9}O?�:zGI�1�3ih�y���� ><z?��\��Xĉe<���*a�#c���[���[Y-lߛ��}o3�`�ƍ��*��מý����m[�o�#�Av6o]���B���}����9�K�ݏ�e%�4w�����~�	_x�(+��ݍ����y��=�גp8i��86�^�m[p*g!ݟ����먫�d�V8nC���Q��K�XJ�SF@�)S��_�OU/�2���(� �$��fD[�Ug���Qtq>Y�N�$��S�{<�%���_�ζ6���"`͚UXm��T6l��u�q��)44_Ego��E�j�)\3Η�5����yܮ9:ҋѡAI��ß@kK;���k��={
o����w�܍�k7a����g"�p&ڻ[�ˠr�o�}��2�];J�	t:�,#-�|�0��ŷ��9���hojF���U\������R��ee(�]�����Hc�}XX� *+��م֎�!Nirgj՛?�����������������! �q�S:gkϲ�����`����Biwu�߃��vtww!'�R/\4���g��r�l�Zt�����������`5��o���Ѐ�e+�?2��k���x(,�="��c���X�b	r�I�.���ftvwcht�
�ܝ�#N� ����z�˺���kE����Z����������qQIQ��[De�c��	�n�Q����G}�����}��*���qo{@���� ]�yS��o�ִK��N[�����8��TmkaV�#Mr��<*����?fG	s��F�#]�(\�Ҽq���P����%��MB.���x��/##�zǗ��G��=�^��y{�ۊ����[o�F��Z�l��>������E۵~�ڹ��l��GQ���3s�?z
�;G�>�K�Q6�Ã��ѿ��Xdf~E���^�BWgN�>���L�{��q�]�����l~J�W���ƩSgYx�/��K(-��@��շ���4�t�DmB���J�?}gk�𓟿���I��T�H�nj�� �����Ps�G�?���k���tQ�0��@/~�3b��-����������BYy�b��f��k�j/bd�_��]
��&��v���in~�K����8N�nBkw�.\���Wy�,��� ��{v`�Ux��P^V�%����r/9�,b8���p��	N�s�kT�2�u11�m	�Ud��]���o��O��Xx$J���s]�~���r�(v��,���(x<{ �ڕKP1o.�>���N���j�
~�WCc#*���l�*V�;q�,N��e2�,��U--L<���p��(f�`P_�j1��Գ���#������(}�~�4_��3'y(��+QT4���FG� \^/6nވ��8.�_AM���[<���#���9�Ԛ�A�sr���y�la4]���+�X�l1֬Y���8:��������I���/^����lΜ��	��/�̩���ҙYYL��UR����z�V���C=�2���F�w 0�P(���N��(9�<�� �����aݺ;�M��9��	�Cc!Ԝ����9�ں,Y��#chliCO/��ׄ�9�1G�b�<^cc�`���asw��&)�D����X���	�@W�R�T�h2p�S�C�n��:��CLFwMQ�\E��!�N��]9�Q��kpvI������<����[���п���[G�t��ص*�������mi
�g��U�P��3��U���!e�)��9|����e̔v9bp�B�{Q>�+�.���K��_���Ǣ%���?�e������{x���x��]x�p���H$F���e4^i���j`������y\_�x�b,]����~|x�
�;i�Sz>�هP�����v���/������s˲�OO�ϛ�����7���:D#�{��]�/<��EsP^�Mm�x{��_m�_|�P�����N��W����gMm]LJYPY�o��gq�R+�}�j��0���0��vB�ap�ytύ�?�y=�D��ĺ�騿|�|��ܹ��πZ����Ƃ���ͣHƏxԇ��B�<��df�p]�i����i4_i���m�?-��q�]�;�_@$�D�HR����ߍ=�nƱ�'�����sJ����������f&u�R}4�IqT��J�N�'	ٍ�zgU+�����1.V��&b�q���a @�Ɨӑb^��H�0�06�]�}��}�������j�J�4���9�NQr���X�x)��:���K��R���Re=J�Ga�0gv�,���V�ZK��[�Ȟ{�Xߌ��/c�~�uu�Y�������=߈����'��S����^|p�$��!$r�W�ɠ��u)Pe=�=�������<��t��z02Џ��(-��(������ő�Ӗ@pt9Y���HGw_��ґ���)sR��EI�}����r��x=n�2cF��H�b�����d������cC�:J��ׄ�-|#jm��s��((��/�#v����&���A��P����D���ڻz���P�$�����+Wq�o`@�z��9�N�kKCY���r��Hq�Pʝ֌ :�:��U!H;'A��R�S�'g�x8� �p��EΎ��3��ҍ�i
�;��.}'ݟ������2������v��r͖�CQ��p8�质$���9@GB�tV�se� �� F�$Ig��g��2IB�sp�Y�v�=�	�M=��(�� ���Q6;��ga����?,�o�ٷydi�R|�/����1���1���{x`�.<��n��v>8z����_����p��y,Y�
������ԙ�X�~1��Z�W�_¾Dl�7��EC��MÓO<���t����P ��,?�rr2PQ1?� �zGp��e��b��jT�����×����9�������2�������!�_�ϟ�]�����p�QQ^�?��ϡ��/�t��Z0�#j�"J=��%�
��m�pώ��8#x��8��!���X�~攕�gO�o�}��ܹ�럟�o�W/Gբ"n��[����� �oX���a�������Ͽ���ߏ%�sQYQ���[5ϼx����F<{a�l?{t�۽��c<=+Ӊ��4��g�?x��g�̦�P[�Z���Wٶ�b�4V���꯷�Y_ǛS����$�n�&6�\37�k�ll��U����8h���X�x�x�u";+�[��hq��6&�͞;[�o������'�t�6=M\��狤�? ���D��2TW���@�Gq�%����=�,t�_���H$�4��v���1�_z��=8q���C�L�\^.��>_���!s�QxqT���7��1�+)���095~����Cʵ�sw�悚G�8&���w�x�n�CԺec;@�e�.�&	��6F�dL�C#ܡ�q214�s{'��F�U�
F��p���t ��U��&�9���X�k���;�p��el޶]��8w�"�z9kbwI����w����LĽ��1t��1)����l�^�i:���n3��5�� �T��ɲ�&�� ���̯�XT�E׀Nk��K}�H����s羙����}�^z�V�TǾ}�gÑȗzzz�C��_�5t�.�sY�VR�d�������o�T�=�C �u�ĩ��Jq�%�b-w�0���M=OZ1)��Պ��I��fC�����۷�Fc�Y�=�r������`Պe�ӯ�#ZZZ1o~	���{���k{���m�p�����J=jkO"����8��9���<�ħPXX�������>8��\��K{`��#��	\�(����>��S������~�a��ոt���.�}��S_@4���Sv{�s0����=p�ܬ(�W��sϾ�#O���x�js�5���{�����^��(���o|��q��5���#��؎�PQ���B���3AUY	�\��}���.�9sy3fbvi!������-�o�;���w��̟� w޹�� ������s����؀��6�5��a��V����⽃�X�b!�>��(6�\�����~z}�Q�}�d����MX��>'���񗥥�x葕���?���6a4H�^��I�D<K�T6�g���?��+yͲ��'SS�B��%ͯ]�\�s �� �<��.�s�\mi��I��,��q꩎�3��tcvi������Oބ+#��� ��Ka~A����c1�|.�|n��j1���l�Y�SE8J����B(d��A!�3������]�9\"f���=+�Iʝ뻱|;���7�QT��G���pɘ9tc�8N*�P�<�9s�_�E(�A`��E�mC(��⤟ �>�9��QXD	gY"X=��XMјL'�?z�H(HJ~��@NG��(��G8g�<	8Eb1�����ҍ��uh��ƪ�k8�w��	]=����"��s��� &#�\�LB!��(]�=gl��z5>5@O9�j
V�YJe_��L^Γe��@e���[�e��L�����S'KI�z<����7233���Ͼ>�w�����е���I䑺�>]@[5��6�C#�2�O%-��xrJ���Q�S4�5��Ȍb&S[2i�t���$7�(�9�x�.$�C��iFz����a����g�m��5غs�� .]j��wN��IgR�칅�����s�pMM-��'>���鑨���FZv62������7pk�Wf�+��c�ˑ?#���GQa)֯[�;�ѱav*ʫ�x�	͍M�'M���0��9����U��D��;}޽9���t��H��(�N�Dfu�||��8x�4~����r��Z�L�u=g,��t/��`��J֭���p���g�-x��7�|�2,_���=�3
XM+3��$8J���Y�r��Ӛ��,��M��a���p��	�M�X���m8A��\;݀C�#��%��/6oZ��,Bc�h�x�@�yع{���q��5Ԟ��� ��I�� <D d�*�ΚL��u�ۺV��R}"9����k�KF�ʔ��!�E�IkK�T`�J�*��}�"�^QۋF	X���p����q��%�<� �U�y�:8EOݐKV<���O����e�ih���"�b����E�����t��OA$pD���90!���Q�fy�a�b�f8Xޔ��\X^(Nr�֜] /�C`iO�gA-��3u��+I���w�v-f�7���������T��I���z���NYS\'f\���ڳ	{�X�p������QX<�`CC��G~�~ޚ�I�w9Tr!�8��H�!A��Qxl#v���Ԯ�gXHZ�l'��xb�@̲Q*��ͺ�~#�7��v^��t]C�u�<Woż�W233��k�컕�=ձoK@E¿��ӷ�"t=p�kA$����ݚ"1�+�e�kjMaO0x7�W�,w"�9%�d3�)���M�ĽJ�����ð�EΖ�81��1�e�c��MXP^���4x=@sS;N�����5X�v-�ڽ6G�# Oy�lkT�����{v����vΟ����F���}��9s�}�[��i�(�=wl߅���q��1t2�.Gi�>��N�[���Ocl$�ٳga���<&�,TwO�9��+�عs�����������<�ؽ��j�ڮ�����$K#S�qFFq��y�WTb�����`�[G��kGX�3� "��Y�s�y���+��</k� ���իhii��P?Jf����͍mlp��3��j>�Oww/�r���;��[s��9�9!R\OO7"� ��J�����Z{�p��]��p�s��$�^Z��D4���!������U���r0ۿ�s� Er$[K�4B�#�9V4 }��2zO �) 6ַr$�2*������)p:�+�^��$SBE�+9mp�h���5J
i��H�����hE�D��IɱS�J_��i�%��S����)e@5���h�E���h��\vGҜ^g�$�R��R�+��|@4�]~���"�Qn�c	*��H-������ :�P��Y��8.t{���B6��/	�H۔L���I��B�}rZ.I�&�~~.�P;VD�D��Jΰd8��L#�Y3�A���B9�RS�=+d� ��<�0�12R�2��1x��:�t�Y����\�KN���!B��Y*+p�k*�mmW���ځ��t,�����#t�Y����=����d����/���t�ϭz�m���n}*�foo�"�r�$�v��3�~.�B{�&�Bfb��e#��${�фa�YEpg�@'�8��$�V�i�#1C=Bo0��m�m�X.[Y~7<.���iP�H(H*hA��|H������ �paJ�%HK�r�Iu�@ �R��:y��VR��!�nx2�16��R��V�8��ܱq֭]�����CC�z�� ):�%�+}Gff��}+�F�Q�b�c����9���	c@8M��x�R����hjjE_��qQ���$��C#�4S>���d�v$f�/]b�R�/���{@�<������h�D~D�~ϵ�p���>���݆@4�`$�*Z�ya#�#��]$E+�N�D�r$���9�#��p�ȝ�v�-.DO�ؐ�㮣�dC&������*�O�%�A��$��ۧ!s��q��D�F�I��[�yJt'�!�v �f��&ҩ'����Q:T"=C̈K�T ��9�$@효���:�#�;䲤'V�M�_`瀜E�ϒ�0�M�	�H�U��ّ�6&�YRʊ�� Z�W���b� V�j���SG��$+����x�p�� �쏐�\��'Ar��a@}�f�C����K�lHm��`h��8<���A�`���!�u����v�,��f5 I;������ԥQ����3���e-�2n0���r;�.�����Ͼ�N��n��n;@_�vۓ�P�7�z�CA���ĭn����cU��䔻�P�)K�ħ�[�&�Y���r׀�tx�f�C}�y�1�V�|&�Q���1ǔX�����l
D����8
#��j���{!%J��*���W���=���M&���k��	�h��ɜ1������f��du9�<�h�D{G�p�>�c[�5�x��_=+~�E�	=ĎuR=1�ҹsQP8믰sA�YxȘn�"C�����p�AOFEh�yK��.8�����a�<]�fx�jܪ�8��    IDAT%����J�҉|�2E=N�C�EE��g\,�(��5QG]���rՀ���*(����֫��R�:5��\��顚�X��m�� �4(JR�������A�!ʍ��1
�؉3d�Lf��Wd/�N^���,�a�u�K0y��g��H/8:7��H�X=1����JRTR���$d$@����7�g��U�P����=��d��$ ������}��y��,aN'�2 9?�zb�Y�Yw�j_�cY��s�m Q6u9����B.[�� "CͰG�H���#�a�E0�Ҍw����d.�I�Vr��.c��f��[���;��v9�U/�Ynn�s�<�s^��=���^���`(�=��Kt�>�I�P�� k��'?��=�Fߨ��[��8)�����(�o=����.�7��!��)�2��kf4O��ElZ��h�3�Wo.�E@pɍ"��� /h\;G�b�tC�;�#ߟFa������j���G �l'���6	�f<��D�xC�˘2$���kEͦ�,�L4K0��}}4sf�ǥ�L�	M�����2��R]���͛'������1uO���X�J���"�"F�T�2�D陑��6�<7\���P����*��"z�B�g�S�Tv��N�Ѕ��ݼW�4*�P��1Q��Is7�'�d>��x�����i�3�{�ӨN���ѵ*�@��:c\�v�@�X���	��Ƨ/��8D�Ҁnk�oIo�p:�!-p��Wy�V)��υ��
�8�T�M�V?O���I�����d��0h�30֗%�����?�X��i]��β��hI� �����������Cr�db��/�	��2g��~��㲑=�=:��H+��a�"���@�qfE��H�Z��:�����z��,..�p��b���k�Wk	W�Cq�л�,\������~��G�}B��������D(����P(����U�K(FG���"���5��z��L* O��;hF���T�)@A ݗ]��͏P܅���\��v�"B�h>J���m4M�減{�	d��yp�Me���,&I?�&co[��l�( ���F�pO	�KK��6�DJ�R폧����I��H=R��[�����UZ�}	���'N�y<f�
���J���y�k�R��1Wy��pG�*2�肙F|����QE�:j@`��`��G2�:��Ӱ�DU�'FG�b���K��L_����l��PJ�ҀU)���Ҡ������t���J{�4��\-Vf�vQ?X_K����@Ɋ!��hkX�_��d����%�	g��͠`f@ ���N�.Qk���53_�J�UΎ��R�ӌi�ԨO��=gy�\p�y-�9[������o�D��kn%d}t�1�c��W"B���a�h�瓲)v���H�A�O���i�B��Y�_�w�nُ��)7a#�K�((����c]��Fa�S�"~G�2SRyN���skV���Э�S�����g���j莎eK�~�0��������!o;@_�q�gB��wuw/��Y�Yz	�$�SL��T�m���ߎ��7�u�蔱�n�.����8i�τ/�qG:K��܆Nőw���t�	Й��;����
r��ĚS�Z����G����P��TA�*Yt5�]G��;W�Sbҋ �%!�P���g����+0]��0l"U*�/J������SSm8����}H>@@�PG�<Q٘�ŧ�"D�R�+��E0�*�����AM�r@��3��5O�1�$�!�L�#u�?7� r�R|'�bsN����N�z&o�H�e,S��	�[��lr��?�G�ǳNbk��M�|.uX>qe4��h]:�F�5l���kf��F��;_֔�]��^�ۅn����ja�i���W��.��~�l�v,��R̮f�.y�fT��!�S1��9ɽN����s���v�G���z`(��y0�'5��I�2^X�";-�`S6��'Ǚ�QV�KD�@t��G�l?�%��S��š�hY\?�����v�4RJ���Z�?t-�օ5B'w�
�py\�-�_%%%{��_���͟�������o�����wtt/��"tŶ���*���	��u!�qw�s�Fk{D���Rm�1�}p�����8��s����iYjw���0)P�c��"LF!������^��Ű��qK	^�e3��&�q�Q�WKqj-��ȁ1�K�f�k��{EO���ч�NV�'�C�y�k;;h2��ʔ.�%���(�~WQ���Q�F��a��FwăH0�X8N��3����uQɀ��|���@N��I�d&�j�`+�d й�A��a������*ȇ����̺Y�dS�N�"�Po�~*L��#D��W��S�$����zV�D,6AK��I�P�R�ڵ��5_��:`���}��V�|�ݢ��V}��'�w���uo��!�~ni&��5yK�o�=��(�'�9]k�/�� j�D��m��nL�^t˘��z�-RW�Q�b�+�T��Tӽ̒[�?��T�����T�ȩ��65nv�Q��e<O`���f�bב�N�K�K�p�&j2�0�ݴ��K�W�o�`L�Y��$�$�D�F:�(�lE�TR#�O�D�B��ڍ�ˣ�����Ӿb�a8�7�7J�Gӓ:Yut"��(=U���q��Z���ϝ�ڷ��go��>�Oܦ��bGG�
k��=+���&DϚ	��W�-�Я��Ǵ����D���t���]px���f�τ���&�9��C�<�S�?��$]�p!�6���d��1͘�%�cZ�Dϲ�9�� �e)A A��b��U�����h�~����uo��2}mF�຤!-,»�\!}��4^��51G��N�~��z���gT�4JWI�NN�sox$��&[�����R� ؐ��@�C�@��[3B�{g!Rǁ���uT�y;1r6�Of�<�xf>�i!kqv�z��i���%r�����5��&b�ԬuT*lh�I�?T̫Ɏ2>ռ�����*p&�[�^��	�nF�r������]<u/4t\m���j����9�i����@ڥ�������]9�
�,�����:�m�_���.$���O�~V�3exX��%Rf��0���5��+1J V�b�Qr�W&��F�^��1��,�λ��P�$��s';�]f�h���]	4\��OM�Y�O �!����1.P���+�>H5t1���pZhȬX�2���r�*�פ8���:�t��㺶f�꿟?��Ϳ���y~Z'w��t�����>�}���cE0��M��d|�xՖK�jO��'o�$��F���'���$�Q�)	J���6�J�7�7�XVv�<D;ň�M�)w�F�rC�!��
��B�����l�Xw���D,F�\�A>1AM����	�k4��&����*�"4�_��g�W�6ø����T�^�e��\Ȓ�#gC����1A%��DG�d'?3� �N�=:�����:����:ܦ!1#.ӢZ֐ʊpU��ZU�N��"uM�s���؄.lߨ�c��=���($��5��0������+{E��pJՀ!6���`�)�8���u�����7Șd�]�dHZ׌�ћZ�j5Q	C�m�Q���$��0a������]��H�+���ˢ"Fyv����<:k�b�;A�Ԧg8oL6S)�$U4��o��k�4AV�QȖ��C(�Ù4��9������-����3�I��!Ā��@�K{��J��(�2�\;5��h�ߩמ�O�� ~9��������p�P8��: =wj[��s^�@7�\u���2$�Н�֯]�7UU�o}�_�8��o�� ��-�>66�����U�P(CG�Nn��c-�:!e��j/X���vL7�.7��L@CŢ	Z���M-=�l���hp�v�%s�� Z ]j��P�N ]Of�X	F��uDʄ!zYU�%'όn�,T#KjQ��� DY���ay�0��0.�����
е�����]&�q�R�J֫�iB�rD����$�;մn�*�����%Gn��OCGhVGΚj�\GgV���ZA��x��U7Evc!0���)wM��Y�e8� ��)P�i{�q���8���8�=$D��[7u�F�����g�Pev�kBg��� ��H�''Y4�XpP�w�c��B�(�R��{f�x��%Rֳ��Sd�5�	L��T�=;y@ם"l�e��=o-��ب�!��'@Wm��(��]����7�:�N�3ׁ��A����5+Q�~cVG��m>͢��Ѽ���xJyM�yF9���˾ր�6�]��4ݜUnU��I��t�е�s���6n����;}�]�?y^|,]� d�n�mp�XjE��:;{�I��oK��mkn���7�ղ%�����?���~�９����G8��m{>5���W���B�V@'P��^���n|��.�;�R�zr��J����x?[Z��rj��BE�bNh�07z��b"J�P!���U�ΠL���7���߭ԤX�J�"œ$Q�~*�^���z�"�蛡+��݇m����$�Jz謰ŭc>8n؝6D��kvd�&����i�����r�!�Q�4*����#D�X�P�mh�&��(F�J��r�+�����/9�fN�b����z�8If�#Q����3? �k��C1f?�F&�	��s�Ιzd��<�E;褕�σ6�������$�2պ�%��% 1�0�Y� T��ߣ ]��脯)쒴��yUո�������9:5-n�N�S~ǌ^\u/����#��R-S*���b]B҄��,�w|}?�t+C�������k��I�e(	39�Dj��K?�-�n'=v�O<A�
S�+g� �7i'�z�u6E��@����K9�zo�d�9��s��FS�L@�Q�����]U6J�!::�tVO��J����1R�S�.�N���:�&�DzT�$�O���LV���b�G�� Ld�'����	��m8Z6m��ͥ�������nC�c�g�6�{�u>S~��|b|l��W�^�#e�&CLh6��6$�+�T�Ƭ�al�7Z��-3I$d}����NeN��bqD�E'� �W��C&Bi	��gB8-s3-F�b�ᰦ-#y����m���E@�Z�l\E 3J*z� eLy�q�Rm|E�������7�Rp�{�Sr�d�d肤�Tou���i�E�/�'?�&��ye� �}�F+%Y5z��]$���B ]�&�˩�,��[kd�IDt>���hB�D����Tρ�l�X���J���%F�<Yn�Q�;"
�N �e^�F��*�#�y��%��dΩvHy=��������(^@@���Y�aF�P[�3��ZT�,k�uM���,s�?�;��PC�F9�*~���w��J�j��6h��K�4�y��W�'z��TR��kD�jcg�75 t��EȈ] &�ʹp;�j�crr�9Z2 וN,����RgM��'j�&N�tuo�4d���<=FF���N�G�2:����β�P��jؕP��T�7"��
�ӽ���g7\�L��
<R��'|�2��,�%�Ζ(9J��ܕR\���|��%����?�2�y����v��m�����=��ܲ-
e��U�8B�zx����p���	����u���?����L6�zAX#x/� �r��#��N:�v�G�h"$B�oL�`>��~��-+��
A��)#E6cr�2|���'�;E�B׃#�>nI���/�ĩ׃@F���X�|iV4e ��=���f��]�@�ɨ��<
e\��f�+iY�e�t��(��f���%=�(��L �Ԯ�QV�d���`��F]j���qBÆt~��ڸF��2�G��9��<*FB��m��R�%�IL�d�Q��q	��rg@#�q�u�l�צ��1ٺ����*�:^tnr?%��=t��R���.!a�u�S:��]����zsM[���6 _S���Uq�����ߵ��Zo��m�M���v���:%/�A֙"��e��1Di@�coR��ڴ\*�BK���t$g�0F�]�GTiQ�G�F���%wVn���,邃ʆP�.4p�=8I��2w(���\ia�Hl���!�\R��+�C;O�d�Wèt����y+�����S���/��;-Х�Ht���/�����\��M�6��K�<����N�G8���#���}ߣ��<��Դ-�PʌIO�8e��~jHq�r����e�'�T~2c��⬟�l��ЦN�hk�+E>�̈2��cTƵ�Z�ixUo��)�u0��eck�F���!��V�ߗ�f�?�"���B�㯻�m���(+�eD���yUC���u��uGH]P�K>�+Uz�fç�Ӓ}7HP�]V-t�isj�bU*X�gdOu�Xz���Q�]������U�;��� ��Й��v�t ]�Qktnd��ԮvrM@WH!k�S��L�o�B�	;ϲ��]�%�e! ��"�QY�2�E� SΔ.�^����븬֥��qjU:��4 =�\�+�� ��u�ŷ�2-��(е)G[����YA=��:Y����W�x�e��w�SL6�bO�����AL4Y��ߕ�2;�&˝A���/W����F����i-i�����wzU�`Me�e[��)����X�j}�{9�J��K�6�q��X�|��?���h�j����������1�c������=Q��@ 0�@U������\"tz ץ�����<��6H�(����ꙓ]�D�4y�*.��1��gd����hn�ІA?Vl��0��ģ�&���L�2L�V�-e -x`87N��Pa�N<�O��f`���X��]+?Q�O�u�ބ)#Q΀��bdU�M��P���'�a��Z!��r-�Zn�I03�W;0�ø�̑�1'g���,Li��U�غ��}ڤ�]"SG=ׯ~㖪��Z�~�YNs��k���n=wZ�:秮C?�M�D�^�}���k�;�3���:���7��o9��OR�#U��z/&��^��ژ�gY֠^����M�U��	�z��Y\V��kс0��	MD�h��e�np�&���uv�f������`�>��Hѹ��R�,�ڴiㆯ�Y��?���~�f�������?�ɧ��|����=�@ 7#@un[�(H�L��>1B6=�d�w3���`�Ɍ��<�� k2P�ę�Fd�}�t��^����j�s�����ޛ����YK� �z��L�d�r�kԿK�7����t@s�{0�H�dͩ ]wr[��N�|��9��:�~�x�׭�%���k�﵂d2���X����N�I՞:��c�/���?�S<�}M��gm}V�=�_ľ$?�����?s#@�ף]�&�έk�I�1�ҀNN���hڴn���v�������8�z����׶���}���s���Љ�,��l<wk��\��ד��Mĩ6|*p��o*@��CL7� � �F�g:@����������n�إ2��Y�S���O=w:���c������x�:��%�36Gb�u;�z��������8=�s9ճ��Sp#@O�c� �z���u/�2�V`��1K>~*���>�] ];3��?�O���hmܬ͘�:�sM���}��#��)Pff!賺��ʪ�(ן�}����vՆ��G_��}��b���?��wttv}�L��O���F�t��t�y�,��9�GV�]��J?��.7�PV��F�u��Y����z2x${ҩ��sI��8�ޓj#';��f���	��Xz��)��Q��4�w��yO�7Zg��X�J�H$_M����9�:Q@���m�u�*�|oƩ�7����um����������N��x3���<�d�r#���t����}��.���S��R� �g�[�;S��մi���m\�����ޗ�ݬ��8��E����������S��������.���C	�)Z�A D����Cb������ʰ[ȍ��nPkt��B�����n���5������ޟTV?7}��hk�{0�Q�V���J�������׺    IDAT��57���|�V �����_�kL���(�p���� �*@��h��2�sJ�z.S�/ճ���{p˪�\t5{�s�
�*(�&1*�(��h�^}�>�1�7�����kL4Ϙ���{yI�I4FPD� 6l�`�������A�NQ�����n�k�5��c�9�>� �w��p��s�5�h����>��m^�/��5;
k�v�Ҹ��?p7�*�]�dJg����f7a_п�N:������W��w��K^�=�[����۷�ޞ={B��5��@�8����"s���y�h��9q��搲N_ǭ�M�˝�"��m�qH~�M�T�(w@�@^��"�]��f+�y������wI�l#�C^���R��-���o�)F���r;����dH~쓏$u�-���o˾�@F�/F��,´ꙗ�5{��G�@6���2��g�˭n�k�5=���d
��V��,z�|�	'��)O�/_}�+_pgl{V�ܚ��_��|�ߺ��w�p�~0:��z�d4��5��b�E��E�)�I]���!`�J��N�뜱��9���kDRF�=б}�d�N䥾y.�ϗ=��F�Z�e0���bl�GRV��s���M�K��9��d�c�M��gw�]������z,�[���<D����@"J[�~��{��:03��N[w؂̚�Ŷ�6����W����E�/{��x��>k��/����p�8̡��ܹ�����#�}��n�$ ����##_>7��3��Ϲ�g!R���������g2��/ ��زh���֘�B�!}K��IHw�C����p��H��Ε$tMn�е`U�S�^#4)+��H6�!t��5�B�@Ӳ[�6%N�@Y�l!�WB��Z�s����X�a��3Qʺ}�?�b8���q��'O|�/�5�y��Շ�z�^��~ۭ�ھ�M�t9�z�!x �}���w0B{w34�c��Z�e9{�2-P���<��DÝ��e��yoLIg`�wr�	�b��!���)�ޤ��L̢Jhkur��y�`#�p��ו�cV��w��9�[�����4�s[���ؕe�k�Э�3�O��C�]8�� t�Ћ����yt ���~��ǿ�ɿ�����_���6�F�5G�'��5'�y۝��s��R���h:�O�����5 �GU6���}��rC������y�*���J9�rZm2''U�m��+E�>�����i��A`��ڦ���Rn]�g�FB'�Ҷh�wܴ��B��'��-��H?�N�k��%>σe�ԥ;���D7��a:̡ӑ��J ��7�;��uB�G1/~��p�n�W4�����L�!Bo;
�o���I���Z��K��gB���ު�',(�2*	v1�7�H��{��tY��ڻ5����Z[-R���me�6B�|��Gڶl�6�����k���	�s����
�B�"�p:ו��|��|��\2��XCd�*��"yw���!o7���Q�t�|��@�;���?�)OZ_�Ё����_۱c�ɔ���"�����M	*���!-��N�3@�� t��Ry���2<�ҢP.���/���q�I]�If~!���.LBd+c_6kٌ/㊱3n+.C��jd��C���C���(��%0��'���-����5椸X}��a��J���,�ϩ?r����]��e���I��F�|�����v���("�ꖽ����w�/>�����N��k_���V�_�ֱ��_��?>��o�
��"I�<CG�n�an�^�"tN�2+�7��Qփ�л��r��9�6I�%t��,`�	������|��J�9��gĜ���m���sP�R���>��~��krYN�b��^c|Fڮ�����l�[��������#6�ﲞ���f�=p7̡��{|ȝ��?�������׿��o�y5�_��~�n{�Ν�_���Ѿs�Л[��*��W�h$�	��:����2v-sY�5G�����/�i���LV+���<��IyZ��\=����FbȀ���\��P���-B�2�y����wm��zL8o;-��1���=�E��{�X���DR�G���*�i[r�{�<�����1v��w���ݻ���8Z��	��ܶV.;)Ns��Pf.I�X����W�31�γ	��pS���hG�#�PL�+A���D����`k�U�<���de�Z{�;�yH�Z`$3Dn��7�S7h�l��/���@���ݟ��������b���6��Mk>B�9t t:)�V�����_�ԧ��K^���ݵ+Y~�e�xş�p�������qI�*\̀���>5D�,��@�ҹ��̄n�w�-���0������i@LC�� ��FTB﴾��(�K(�{��E�2X��E����j�bh���.+C�z�O�B���>���|�P���g3t�C����������G=���xƯ_��W<�����r�_����۾�,ڶ�A*B����P�P9��r��g7]3tx6��}e}��.o3w䐓�(���%Ƙ�	|9yk�q2���< A�խV^�Hܮ��G��r2�P�u��ֲm.�=�l��!���mȕ9�ߗ�_��?�	]���bGbl@�	��)���W�5�-� ዻm.f���Y�D�~�ƣ�?xړ�v�z�Ҝ��2��;v���e�<����!tn$ڰo
�]mB��qjM-�� ���|��|�+u4�z�Q-C_�E=���������/����v!G�g�!��!�X��m�[cH#����\��<AL;�C�}[AO������r2t.�X����Xl��4B���:��V�����L�ȼK�\������c�}�S��_ևܻ*���v8X��֐;E[H�(q�3�%C��n%'�P�!� ��Z�C�N��;���k��2㑸Uw���i�����z�<���C蜈�K���L:�g�m�d�e���'�/˭���\)�����z(q�zv����5�"t�t������p̣�~�Ӟ��K_��(�_W��rB��3w��鶭Ѣ8TN����kΣe�����a9qL��(bI,�����%?	��B�����|1��k��߄��
 -�t��O�V�R��~�'s)�ƚ!Y�x�kW�-��-�od�>BR2�|e���IV���qGu�	�-��Q����=)K�I�^?���?���O��䓟���"�z�����r�m߾��;w�x񞥥C8���U��"3t�B(��n�(�WO(��n�1���S��$$g��d�HG9F��]��G��aL���hdae�Ф%�w�_L��eT����Ƀe,B'P�.�����3�c�H���\�=ked�I>>��:�-Yx�!��/�j�y���	[B�W��z�uG����������}1mZ�2k��_�'��vǭ�رc�K�Z�N��T'<�6��!�PV�s�y��uBoK�)�'Z=�1`#C(�e����`N0���V��T#t��1~�#|jiO���&�S�K�]�ؕ$�OB�0o^B��\LywB\��kyy��C��^�C��~�w�������Ͽ�����t��J�_{�^e�;�o�2t
�q��0u��(���8���?4����S�H賀��.��1{]�u5���W��})��q�C c��Zo��~י��t5�'���B>�.�
i7��44]F�BYT�{l+���J�k|�rA�X���\��n���1�&����xs�Nݡi�N��iz�*[��!���g� ,�>�P��>�}i����R�.u��-����}X����T�t@n,My��\>Tw�n"Ǔ��h\V� ��Ce�U�y�M����#��ٗ�ş��O�ӇM[�"k�����⸛o��3/���_<�q�ۃ�s����U���Dw��G��c��P6'�5`�v��q�6�b|u��$�F���ug��a�'u<+�#�3F1o7��<<�L���$��MT�/T8��!��/�*�J��Z��8�jSCvai�ŁF��m"x�^,m���sv�ʈ	u@R�ځ���֧.A�+[�=���@�F<h�8:(����;�59?o�h��τ?3|�D��-a�Տ�ύ���
� ��
�%i��߭��*���ȸq��gM�C:A���B5@���2m�YY)fו���6*��.R��9\���뷝��U�[�>v$?�^6��{W���/z����W=��O���?}���u�;����7��\���h2��m���#t<��EV-�E�h�V�LCd��� �U���k��9�pYX�UF�Q�'+���&M1A���*���5]�lɗ��!\�V�+�(I��mY�� �]�8���u�������L0���F-0TFpX4�ӗO�:��Bz�K�۔��X���q$��S����E0d��b���@���v�@R��Q^��tקB�8���Ї�^~�>��>���g\s�)������Ys�����ţo���_z�e�ZZC"eBzsJ�#t���̜z�`y�B��N�sQ���K���"C���е�����2�.�%AN��3���Y�htLPP�y�,B��٘FR>�lg��8�;ձNL��z<�Cs�s$d��3d���%t���F��G�O���̺�2l ���܆I�\�O:��c,�L��o�>���dY����#��#Y⸥Z��*�b2q�>�N�w�^��g������u�U�v���.�&	��[���K/���=K{s�	J�C�ȪZԐ&ɤ@��"���F������I�Gf�����vU�|�J+@辠c�	=$�� 1D�m'm_\j����V�S,��:c�����T���yGB��	w�MW�	�L�s�	0��c��|*�o��DdD{��`����b���}͝։�W�~|��i��r��p�����/x2trw�\�����N��d�2tx&�ӥ<�v��'�z��2�}�_<�[����^�����>t:-���RdլR��D�`fx1=���y����}l��+A�1�Yn�A�����󴯎��!AM�2���O�&��&x�| �x�.���v��	��kF'!�G�]	xx�f'!���C�!tx���&�L�o�>B�����L;Y�.�@#t�)sb�6�1����p���I��/K~���%��k7݂u4F3ud��s������$+_x�-7\��Tp�e�|�뎽��۟�c��/ݽ{�!@襛C�c_�qBϒf��1T��I�C��At%i(rp+�o_WB�
�1 ��v�E�Z�jg���Ր;E��Z�jk���#��C�����]u�I����s�@riH��^:���UK�4�f���U�F�gV��x���q=h6A���W�u��c�)dG>�s;�� eo���m��!w-�a�i���_CA�����X�(���eר�8��rO�&�g�t�Ѓ �x�K_s����̝�_�"8X=M{�PI�(`�L���u�	=6���KW��q�vB��+��sR1�ސ}C��|��څ1��k_�t�JB��Jzl��P,�jm��\L��&��Y�w$����g�\�+M����j:'sm���6�K}��m��^Bv"�V��sL��&Co5�	nc+��!CO�rg^d'�~�z��������;���.����YZ:.�l3���I��2!�G�p�Qd��:^�3]	�z���X���6�Ӗ��CHN�~�'�f�;oy��dL9x=6�%���Hq��2t_{��|��zȶB����?��ҡ�{_�n�E,��Vbt:/�k��\&2ؑ2�ɚ�����H7��5��]��g�T��$�'��}n�;�IGB�ry�ޗ��t����ۯ�~^�Z���ܐ���ʓ�뻿~��W=i��A �,�WC%͡ ��i9���C�(�xBE�1
	����P��z���8���� ����{��c���#}q�����|��+����䓏�q@l�;���>m[��N�L��}�:ۖH}���Zmd���\��(
�4��J�7�vJ�sL�!t+��gݾ|:�� ����@���B�n�:���F}���I�����K��Y��o^'�l�y�s_�Kw������kg8\:�-8Bw�;at�V�gi2�}�(���DwB�!�S1�K�#���8>p��{'T^�Љ�b���EeHB��q��:�[D,���'& ���c�ە1�Э�ɳ܉ %q�le;b���:��p��z�F'`���$�s�i���컖M�Kܒ6+(�/��}溋]���A�ܫ!�4���^<	��;hF~���^?�q�߻�L�W�v�u7t&�~`�e��y�K�����7����g���"�~}/�y��w����$S8��E؅ra{�+��'���u~�T _���$t+P�U���g��9��`�T�'������� Z K�����w�
8-�[O�\�ЛyϘ���wZ�wȯ]�*>j�K��
��4yʠĉ��Ϯ#<���%�z�:�z��Ԓ�H��D�ݐ��>¶5�(�O�ߝ�T���D��?B/��n���c�f5ˬ9B���?����ǕW_��h| ���d>�,ϒ�K�ݵw<Co�$�n���e����ei����9�&qu�f�ǻH>`������:��!�P�kzΗ1��蘡�d!��� ��9ط�g� ��D���#t7�sˣNg�Z�����X�Π���G��Xf�Z����X�����
tb��H�t���5��OXd
���lG�����`Bk�e>bBo�\��/f��Ы�0�]K�~�������:�Ǡ�(�~�~���\}ݳ���N��ʽ*q�^[v�(�ϡ7U���}�I�sǏ�<CѼ�,�I�r<�]�����v�^G��j���b�c�C�-��iH6�L��*�v t�}2��2�,dv�*q��/Cӂ�5�j�G?l��аE�f�����h}�A�ϖ��q_e��V�b��J�]�=�h�<���Ҵ�I���X�gjo'��F�|A,L�� 8YZ����ҿ�s�GO
7������{�ד,yͭ߼�滪E�$��M�V�s���'|��w���\���hx \��$H���U�8X��C$m������]�x|`���+�j��F}7I����ݮ��C������)mj9x��'O���Fx| �و̺B )�[$�d#UOِ5|"�"	�G0$;/�+���p�Y�'��Iqu��Ņ�m1��F^]	�}7I�>e����1�(Nkk������v��B�Qi�\�@�Tݸ��4�y�D��־�7v"ߤ��{�ד,['��´��ܓ�{߿��_}���.-�:��"�$I�Ÿ�}�ϡ[`Y C���΃
-��g}��)""|��Yir�!��R;�OB�sĚ�9Y�H=6������>e���5�t)AU�;�~c��G��ή�C:� (hX2XBg#H^���ob�e��O.�`�U/�'��2XՂYR��]�ҫnZ��8(��'���׃Q�,���irW��}���׮g���������ݻ���e�b:Fᄎ���pS�k@&)�pc�H7�k��r���cڠ�<�]��y�rr��y�"���}de:�b����<���G�w�K��^f{��M,).�ЭL���տ�@�G`��FR^H���G6+	�HR������mk����=hAN(���YZPk�,L�¿�h���Cw��M��Ņ�'?�	�1���4y�w�q�7Cm^���ܐ�����_��?���^s��.���*C�g�����ܶV�2V�?P�.�G�>��j4Q �,��. �X40��Dc���=��C�i[GkJ0�!ܐN(B�O�����P 1�ˬN�GL@��G�@(&�j�'�,�XB��;�'d�V���hv���w�����oc���Jn ��p�������dÆ��{�I���s0�}�H�ׯzW�N�D:̡�ѯD�x�f�����9t��Y��j��5ۘ�`����?� ���e�o�-ʠ��5Fu]��\�Q�LD���V��g�mPk�K>�������U#    IDAT×�H���HL[AbD���>�=��A�/ov幈����K�p[
�گ]��71���Ī��8zW^XC�!�	�@y��ٚ$Q�{^
M𽵋D�݊��A|�ǉ��jX�ߍ�c���mk7.&���Yz�$)�d���n ����7�������!w t��Y�:,�ʛ=X_�^��~��q^�������z�v��~5���z(��\�v�.	ݺ�ے�E4>�О����"����]%�_��!�Ѿ�ɪ+ԗ]T���.�.���
,��ʆv�H�XSq�"ܵ��i�YMB�tk?��5��.�ӂgw � e{�����?'��}�?���������+����o��ؾ�V�57�����~��߸���7\Z:�m1H!��{�O��ë�9;�hj���Z�2:���g�9�-d��Ź��Uv�r�:X�!�y�?�e�1Y��O��53�߁���%��B�w��̡}>B������K��ʭ:��U�|,̱��
���(d'3�*��H�ے9��}�0H���m:Mz��{و[p���d4J�޶?�A�Ņ������uB�ͪ�s�����{������ޝ厄��9�s{�]NޞC�mk�@�:`Ͷ��ľL�j��"�X�>ЄC���tx_W��5��Da,�2��l�G2�%t��!w-�j��1��k��U�'C����H��El��I]�d���}���:���=)�%{���` t�j��4B��/%B���n�˼���-��w��K�č��Y����_��?���]7�b�j�[s������y���u�u��ޞ=K������,�I1��]ƬrOݢ�	��T�j���5��� 5����r����2kʡvk�"G$������۸�o�+E�]�w�=�!q���H��P�8>2�d��Q�[��i��~�Ƭ�"t��p�PY�j�	�TKg����B� �.�����EN��v��Iw��~x�B�������q�#��h����cѳ��$Yڽ�-�2l���w��M'oX���S����p�]?��k�����{�`������T����>B��)	=��E������ݬ�Ӝ
'IQ�<����,���d{}ν2�>{��<2�XEl2Z&�	QV���й}��4ߪ}�R���}�i�-mlB�ȅlB��kA��i6U6�i�d�aB��c��ޅ�59j<3��}�x'_���s���E��� ��.���;��d���&Y���,�\лu������I}�����=���{�{���^�b����#�a����Ē2��e��B7~�k�x@�q��s$	�]�5$N��=�(c�C#Q�m�2.�O�[]B�M���gz��Q��^�ɮď��n[���?%NQ;�����T�V�.DvӪ˽�����T���Y�b0V�K��.���mi:�-���C䜀eP+�)js��G�Z٢%/�l��v-���F [FYw�쳹� V{C6��������HV�Uɑ/@'����N���S��m��登�(빹t mZlg���>wMu������..,|9�do���K��u������y�ϸ�ʫ_��4<�}0XHpރ�Jv�r7��V���9�@@^�޵�Zy+�������:��\� �;�[��ٯB!򛕢#�Zo�)g�S��l��#�8�9�͎H�6*�(H!2N�������G�.�i��&D�]�#E-��#�g4����z�懜��� Q�G�|9'd@��wIj�t��/����O s8��۶�O׮l�K��k���-�E�钂-D��\��W�:�ZS^�=9����������*w�W�daqp��_N��ϯ�u��z��S���{����˯|�p8<�1O����e���O�,��O%���
|����#s�>����ड़cH����:��2fZ&��D:�fo�s�I@Հ(��q��tz�ͪC.�B��gCA#�\3�B�"���n��f-�Z�oqR��P�sHO��*�S�;���	N,���}hm�W��wno��S��ߢ�ZvR��H�}p�!�@r��.�YX\�u���/�i�uB��8V�U�z��o�������;~8d\&x  �p�����a��&C'���������9IHP�N��n�R�ifUsz3$V�+M�6X�Y(��k�Đf�}1���}�Z���b	=$���X��j�F�]��y���ZTi��V?ԧɇ����$���J���'F<���~�����WI��s7�����A�sܫ�Y�Mk%^���a��w6m��,�b�z�ޝ�������뮻�i�\��u���̮{��P# ��NQ͡?�2l�%A�IS]"_��k`��|��O<&���g[2�����E��b����� ���o��/��e�>¥:c��
>�zl��>9Yz'le�	�vi��F8Q���\^��|��5;��ѰBf�<s�l$�W��0�.��O�Җx�*q��/˒)�-w�0!�� G��z�ܡ�ƍ���kӦ�H���ڵ�K�C�ʧrox����]��{�%�^����g�g�
��@q��4O���?���1Gcx`2tiPҐ}Dce!V�H� �^�zW�.��u�4��jR(�u��[����j:��7$.�ie{�� ��j���E,�k�[r��"���r��}��",IF�Z� �	��b�*����pI�<��)��B�.ej%4P�
�ӳ���.��IZ���!C���a�	}÷��{ӗ�^��v]�N�1�����f��]O���_?e<��$���4�G�Ð{���M�����9���:�E�T��1�!�X@���u�>��r�y��J�&(p�j`��L,�[ �Ͷ$Q�21�ǉ*��]��A�V��s�f}��4S�oe�$i��l��Ҏ�{�{m^[H��^~f%�y3�s�Drd��yg����+��!��)���	�׍�������:p:�a�M��y���1Mҿ\'�94��~�\����2��C$����4��h:bs�:�cVXm�	��r�Pw,B����Dx=�]TW�Y���ק�d�"D�2N"��V��C���C�YeI" �)��J��cݒyȖ|��E21�"�\�����N�\�A�1�"���e�Y�\�������G~rq�����]L����x0�}O>Ʊ�E�{b����<ZW�2t���U���{�閭�n��ֿ�����f������S�FB��W.��%�Н�����!��ĝ�΅Z͐{S�}��|�ϐbE`�$,+Z�}�/D,��`��J�^;����!urd�,倫��]�[��� D@Ieh�����-ғ���k/]��"���q�lV�
z�C�V����Ez�����{�$/�Х=������W��Tg�L,=�p��OI9K���O�Ӵ��Mb(��!�}����m۶|>+˿���k�X�g�&�_~�\�կ�����`Xu��H�f�e�r%):�g���fo����c��#t����j�`�7DL�-Q}\Bo��c�n���Fh�h.�@A���1���>�8 �Nx�6�ǒ9�9x�Z��V�"�.$���g�wk������]�R��-p�m��V~.��q�ХLd}���g!���?����C�`�ZwE���pq�t2�Y�e�>��۶/'��\tѧ�	=��{r����q4�,$�E���e`:l/ �&xҏ#j7�a:$�h�G�!��EaX�%��0��	=$+-ːm��mF(x=�iN�g�12��
��s]�=D�>R�	Cr�������� t�.|�������4@H�X������ΐ�cecK��I&�=�r�_��=�Yz'���g��
�<��U�[�n�����"K����v��clx5ˬ��/��G\qՎ_���K���h��d�$���6�}<��8�>U��³��9Y���kDڕ�B��޿V}F�e�E�{�.���}��d�	�ʄ삲��I#z^���B� ���� U�'dwZ�1 �ksL�{�wZ��կ}F٨���cd$�#���~�gZ��iW�syH[�C�2е���I���w����Fmֶ ��n��`@�ٹ$t8˽��d�*��[6�p�A��:������Moz�a]|�/_z�5�ק��,D�d��j8�G�R�ޮ�r�!w\��3�.Q��q�����%-���4��s�n��:B�h��F�b�M�Q�Z�%8�H��-D��x�$���K)��`��|��J���H���99���.����l�"XM&��	�L,�/�У��[��8SNL���\[Wa��կ�~9�����{moz�N}~���5=+�����+`�sx48,rK���sk��>:`W��˸�dq�;�lݺ冃��ߦy���=ƃE�7�����K�����=.���e������v��>tr�>�+��7�/g��ⶭq���b@[��s[e��Թ�h�@"r�7��vX�tf�� G�ʒ�b�<_E��34WN��m& �����BJK��=���<АA�ր�˄��aj���!B�t.���[��x�-З6�e�ϱ B�H3��-���,c�q�;4��l����쇗��.*�+x�o��Έ�ɗ����C�o�+ i@�Eur��s�^g�%0�~M]�e�k:��<��/]������j�YsC�@�_���O�l�ο�?:,ק�5w�0���K�C�}蜰Q����,)���pc�`Y��UF�>���}m���!��}�ߵ9n�i��=�����ѕ���&j�Nҡ̦�Ͼ纒NL]Ɇ��ɕ봋�:���`�o͒�ޅ<e@�VMZ`a}|XAn�}pB�d�qI�����H,����ʑ,�蝾5!�����s+��x!�����IZ���oݺ���:��2��~���U�_r�.�t����(�m[����#��*�&�\ۄΝ����_#JrID�4 \MB�5	�?�:b����J��/Ђ���#׳�1|Ƿ"�C�!Q]V��Bׂ(�I���\�Iʪ��Ɩ�D�Vy{�k�R7�4}��ဆ3<����r��m�얗�~N�i#m���0���i	�H�}�D<��e�[�?�>7M�7���Z;+�~�ŗ>�˶����ih��0-1Cw���	��<ۃ22*��PWB�C��#!B��rd��9<�V�p�5���fp�T$�z4���|�N �J�>B�!\Y�k��'��o�NCA��Jfn���^���<k���%gn��?����<����G�$���K�sM��s��d&��#t�.Yg���8:�Z�C��R%͡W��>�c͞2�!wN�nȽ�<T�.���!�=�y�[�B��E�1F(˄HM��%N�vv!��,��}���%tz^A��QDҭ��������im�e}��X ���&�-�h��:F�}���^mȝ��l�v����n�;��>͎����,�����T���Գl�F�!]jdN�j+�M�Ô\��cp�^��0���N��r[�l��͡�z��>�>����k?a��3�Zs�].gi��L���]�28~1"�� t���s"^.&8��E u�K�ײq@���T�%w�^�"�NkX_�ZD��=�l��8Z@�g�qҌ��G܏,݆%��pB�|�|e޾�<g�|B�t"}Y��';�M(��F0��H���r��d�+<xp�v-5rYzu� Bϳ��NX���;�.SN���,x4�-��>��?�o��?zk��W�̚\w�E�>����H:-�#e�!w����Iq4��`#t���,��5�'��H�G������Z�,�`Ef\����¹ځ����>Y�'Y�/������"�]ڒ���>J�J[} ]�W�d����9�Xy�tS���,R��	���}V=��g��2в��_�@�Y>�����	��
Z�au�{^e�x,��	�ܲy�+:��Ϥ��۾��O�z���2n�ZE�0��+�ʝ�4)��ڲ>˝�[:.�s��6Ǖ�9"w2� -0���"OY/'h�}PFnײH�+���dA��,D��,���9-:�j�����ӳ�P$ K����}�C(�!t������}�#_P���%I���y�,	&V/�r�2h��Z`�٣�'��%FGV�n�8/�a"�]j�=�m诫'��pϝ
)C�������E�e�'[�l��C�T:-N���/�m9��Ϯ�]#�:�bs�Na���6h6���0��r��LNIr�!Z��3\��5 �`�\B��4�a� m��ne��Z�ẘo_?k��,P�ꒀ&3�����d� ��]ݲ�{���')���Nn��V�Щ!�Z6ß����q�O��e��e��r[�e��~C��uI�J�f?��d�|������#t$i��e���>t�Cw�ܷl�y�a]�+�w~�s��=ƖW�̚#������<a�e��֭rwC"�z:����;�r�}���Iq��w=X��"t�5@�@G�HP\��4�[Ni��dPC��e�\�P��ǀ��(��� D{_��%�� Df>1�Mlb���|���s\���/,��2�/�b��UV]dbٍ�pB����~N\Tm�v���D��֬`Zӛ� Br��'8��̝�ޔm�Cw'��$%IKw�ɖ-�/;�Ѓ��%����G�m�j�[s��ַ�q��?��_ھs�����:pvC�}'��Г2�VY9]��&tw����h�u�Z��-g��JuY�&<���n9��Dl���8>P��ͼe� `B������5��b���j��"<��d/u����c�1Anl�f��%��ws���j̡�؍/h��d�"�^p��[����[����n4s�v��cȦd��78��;T�����;-N%���}��7[�n��C���uB�?Y��o~�_�җOڱs�?GD�y��*%41��������~t�@��92oV��UB�A'h��g"��c	��/ �E�1�ւ�XR�!tF�w9R �Z�50���W�3�Y��קe7\�2��E�i�c�5D8�`�G>��%t��.���c��Y�fdۺʄ�ʥpsǸ�Wr�|�;*[�l�&��De��|��4���t#m����n��������x\]��@>�6�pG�oݺe���rA:��k}Ƚ�wTe�пxҥ;v��x4~(�F�r<��t0�<���I1��_��$���a�Zc�x�+��u�{4d��f8��n<et�9 Z���mP]�9�`$��`!�#D"s�d����	>�sd�C`Ń+��>�0�d���9u%,1j�d�E�����	ɗ�\ɕ�Zy�-���0X�A}�"�F_pٔ�d�Y �"t 47��&tG��1��r��aH���Z�A�4|O�[K��|�pJڍįv{�uP$S�6��zw}sw����I�a�;�0CBǟ�ݶק�Iq����=䂤���N�s��#�|ҥ�\�����e�)C�W���,��0T����Bgt.c���g�{���
��ڕ�C�I�>-c�2����*zN����$t�Ƿ������s`�dHg���g�:'N\� �g��V8YP��y=�ڽԁO�>}i6n�]��yo3) ���5BV����ֈ�_o �
~J=����4�:�)N��yjz���2�;���&\�ƿ����{��^�j��GP�D��&�}�E}��~����������O|h}Q\WN��޳�g��v������a0������8 t.���0���K`1�\0��`P��^��cu�j���!!�.����]�D�9YkY�, �6H�҈=q�愮c�B�-똇�}��&��x��P4���+_)�X[�������[�h�,n�r3�u^}R��z��	jt�4f��q���%Dz��i�e GI��5�v����� ��)�,<��M�����Bwe��)$p�'���[w~��yo��c@C�9�Ӷ���O��+�>NG��p	�9��(2�Лa$��C퓠r�.���p�� Qs�P_�~��:|���'��C��6�2F��w    IDAT��3�(�e"�ݜX8���^�|��-�#�l���j�F��S�z�u�6���Y��С>N]힗��[L��&��Ydg\�O��,���%��i�	��N�!d���2)����h�w��k���N]��������Kҟ��ݻ�?�7 B'������w��}9��#?�r�>�>���u�Y[���'O��+�>�^L��2�����h��a�Z=����>o�WZ��F���M�H=���R]�9_f�sp	���ϥ��3F^6B�͗�@� �g+>y�pr� *��V}��>��F3�t�#�=��-����$���բ!�t(+�!t��2H�� ��wM���\"�f1��֑��?���`P:���X�k�.@���n��_!9$B'���z$�oݲ��#=?O�X�C��+w�i����O~�ĝ����YB�mk0�s�`A�g-B���Nr����πb"p��-2�+�Щ�ƨ���Ev1uǔ�B�|��n|�	���B<���-bv�ɾZ�n�/��C��Y�F\�/Đ��9N�!���#��/�8D���q�����+�8O���
v,���D�:`$̡�����p$J,��{:���+���H�lޒ�l?��5|���	�� �K�H�-[7_v�a�~"+�w��CU��O?w�G?����SG�ɑ���	d吡c���c	����a��Λo9{�� &7����K ��l����V_j��ydB������Z��R���#&C��L�t�
����"�Pp$���w�-j�`��rB��v�||����8-蔄̓�����w't�?�po���مva�:d�|�f��8��q'��w� �Px����'�fd���C�}�/:���>�O��}��n�]�f�5w����w�:O�����z8�ER���P�gv�HW���!���;%�j ��XW�й#��C@�U�1��!�9Jҏi��m,B���t��ec1���`BA�fg��.�ۅ(-�C�E,q�K;C�Y�����oi'�{�4��g�����z#�̝�1h⍕����sB���U�����׷��}6���˄륚�u}�Q	j{�p*�c
ܶ�'�m��G��Q�}���	����_q��SǣɑE����z�0
ssA)����ʝ������" n�1�h�F`2���~��/0�et���z|�y���鹚"� F�� -��@>��%wz7��\G$ŷ��gKR��~4�p��1�hjvF��]>r��˂���,�M��nb|�;��>a�3�G�h��f����nw�vQr������ʍs��uM�����-�����cU��9x�+�]:�]f�$t����{�Y�Ok����n�}��~�����s�	}/8�s�����	W^}�ic���	���m�Hq^H��Com[k�x��YB�nu��j�B�@�;�$����SO(z������B�]��U�T�o~�'y��%��p���Ђ������K�~�:�Q̳�B��IA��i6Hz�:�j!���b3� [k'ǈv G��P��uX�9�a��;XF�Co�F"�F�g�������O�|�A�~�Щ>�-��I�� vI��>ӑ���{$�� ����;��������X�o�#B���]�M�őp�LZ퓤ݙ+�z�:��U�.�(�O�(n �@%�45"ZmB�9V؇���H���x �Gi�#��E|�}z��W���r��y�e�f�99K[��?-Г$:��ҪmZ4�d�+e�>�#H��/�O�����S3.��Y�=OdG�p���7D�΃R
hyVs��9��E�V�,B����L��ɏjȳ��`�����}��D��e���Gq����*����#��+����	�zP필9tG�n��;T�:	��і�f��a<�*w	@��ŀ�^��y	]�w���?n�=c�/X�	p49h�a,�t�%�̩i�h͡K]P���'X)�
V�+��hZ5��ː.-B�z��$g�w4�j�m�a$�?I�Z���~.��'����8?�2Pro��!tm�;�		��Η�4�N�������G�!�s=Bۥ̡�d赿�	��'B9B߼ϥ�~�'�ir��*�-�2��z�^��{������5������r��i]�� ���*��o�,�C���^5&�Ѻ�.��9;wx�=��H`#֢�.�ե_�."��\���������3V��<�$c� ���/���h�p�7���"g��b�/��$d�����(�6[����<e�d#<`������\��ԑF*\V�/C��ET�z!�7v�����U��"+$[��6'�i6Br��lg!��������������$�N��>����
\g ���^�p�������|y��Ԑ�f�?��7�y������ϐ���9u�LJn�!w�#��y�b:0\�*��t,CXIB���G]	]�͐F��'t��j�{B�wQ0��CRK�6j�����>�HB���&^GH���V &�ɉ!D�+�o��|}���G�$g���5��L�lC6
���Rym��l��t�ۚC�]K�s�ڶ5���ko+]_K�@�ա2xYW5m��%Bww��}�{��%���'��/�����wU.��g���o���x-����a�{E�|:\�R,��8:$���о�G:Rl&g��!C�|8aq��l��bȎh0�oj�Yʃ��C��]�-��$h��@�/@������ʬ)FF!���%�Hys�!w�X5k�d28�ڣ�Rf������6�gx�bz����o[�����JUH���y_Pҝ���`9��~
w,e���v�Ы}�Pv����䠃���g�g�!m*�����:��������;:����%�y�����8U���z�< ��*w��WL$8� O����x{yv@�-Ɛ2:8B����]�Y�W���;e��Yn[�u���K�W���H'�sxJ�������lrŘY9qQ�gn#�]]�jA�e3�>�M�7�%�cr"�G�Ɵ�A��"o�k��P�m��a)�#O��0Ё�\0�iC�M{� ��	on:���*��!ˆ|ղA�O-l���፜�5v���QvpMw�l�g�uB)����瞻�g�︫v]w�x2}?X����0��OF�x<J�����pQ\�H�7��;$��m�$�	c#Q�!Hp�CYm^��G�3$�}2��ZA�A�{��\&1��Y�^9���5;��"�COL{C:�����"(��@5���l��kߑ�h�ϸL�-s2�K�����C�}����t��!��ۄS�3��,�}���NUsǭ�Ccڗ����T+'����ÊX;�ѳے�?��+a�s��%�3[�l���C�x��޻�(�:Te�=�{��=�t�5W]���x��9��}b�{y��2G��0)��na�Ӌ CCIt[� �޲k$sti�n�!`�F�9 �zD}dC�>������%��u�.�+E�1�wAŐ8���}����^L��2|8�k	�>�ʠF{���d�K6�WSk~a٫$t�>���o{�����t��ݶLhQ�~R����>۲mg�dw�_͍�<C��K��V�bqZ�C� ��a[���`(�}��-~����K��~�S�����,�i5[бnr��8������3�6�cv���)�p����j�Bu�>�\ ��j
��XC
u���"smȽ�d�iM2��uj۩d��%s):Z��HC ����\B_N�}D�YY���X�3�\��tו�y�Ii�,y�c`�܍-	��eg��y ����$[��9��Λ��ͭh��V���P<���;�na��?�3�o�0Շiuܘ�ܯ5�~i�	�����,[�n���~�ǲ${�:�w�D�$��~��s>���|�o�{<�%�����:,��ܧ0�&t�G�4#� ;� c]9'12D�9pg�2^�=s��u����O��`C�����{�,B�Aں�]\!ߵ��U.����+�[r��8|'�M��0$)_z�|N��$8.�P;�vF��(���fm���v�p6���W�7�hꌵQM�2{ֈ�W�f?��(�$�v�^���T$i�%a`�d�}�|�gr�G{e����Y����瞻��o�17|�3'��Sf��vq2t6܇s���8)noϡ����^d����$aj]e��%��;99kC�D�pP�m�%�9T4����)��:/#[JZ����u�
�be�%[�H��.�2J
�4R�v"AWʹK{|�-���btd� �_��@2�����
�,�s��*�X}�m�:����m�Л2�s�(�٣_�g���|�3�'�k.C�pC�0�������D����f �a.d�.�DB[ٶm�/=�!G|���?�����{���Z��ܐ{M�߸�L���H��7o�9e�&��ĝg��h:f��IqD�}�Qل.#�n5�e�`��Z�.A�2�!K�>r��'�j�5���йd��#�rX�#Z��0Y����Fh��i�d"3��"t�}D������m���O�2h�d#���a=�靯����~��U��\c{6��:<&tz���c�*#�
8��������Ӭއ� �+`�d�Y��w�o�}����>��~���y�u�r}a�ϯ9B?�/,�q�_��[n~�d\E�Љ��*U��G��Zhv�9?X�Ϣ��)�.�����S�f`�S� ����:% s����!���I��|�"z	��n�y%!J}��]	�n�[���H̳ڻ��8	�w��䴠��v�#PM�1����������C�`(C������?k�@��$m2��ȳ���i�b�{�G��,>��F�$�-jx����������Mj�D�H[I�e�;��з~��{���O���z��E���:k��|�co��MgM&��CR�}�8��2�4IF��UhH����wҵ2�$h�.ԍ�[� A��5?I���@.Ƒ@�#�P�BA���$	y[��?��>�л��J:'	ޮyH=��P�F@'�\�A+(��[ڞ6BYU�w6�<:�	Ȝ��F�ϒ�l0����\�<���rԂ�\�xLk"����R�r��Dn��2�����֐���V�-�
�m���n��ݝ�昝��z��怲J`�N���zɾ�n���q�zi���໾�7W�����Z|���o~�dZZ�U���S�dZ:[��b�V��f���sf	2Yh ({�N�r'��9�K�T�X���@�����ſ�!�J_`]ڶ�eC��}��קGI�Z�G�'I���W���k�I��}S*V{y;dP@�	\��=r��ǒ4��ϸ�x�Z}��~C��1�����}�#�m��a��!ɩN�$���
q���\>!�ڨ�Ϸ���y<7�-�ˠG����D!Cg�#�' tw��'e2�!��=���`6��_'�8ݷJA�~��s��7����(azY:."����h�Qx��>��5͗�I �����h k+?NZ�c=ԟ9Գ�G|Y�Vq�k$��%��t�:"h�!��4�堩���-�®����/yp�Ͼ5B�N���!�g���~��ޞ�Iw�2��h�$��d�0x?C~4�X���;
"tqz��ԧ��&0����ܷm���_���>8H�}��?XN�ĳk6C���o���G�elE�d�g9^��Ӳ9��uw�7?�C�! � P#}�h��	<�b=�1i$�Fg�q��QW���E��4���zdVj'>^V e����j}
�"�/�h����i�3<'�j:���䩿R�1�x�/k�q���hx��?��Cvb��jz���~5� �0T��qIuV?�C�;�`}�m�}�Q�~�ze��B#�{�C��[���zu�;E8�y�9����^B�[�J@�JA-�3���@%(Q�|x��;1��5��z�ٯy5V��B�/�]n��\B�y��]�^���Ԛ�id�J
�1��x�X�J?�g�q�'����q��/@yI2p��[����G��>���Y��ۦ��Y�r0B#t^�f������;����=�	]��ܶ��3�~�#ߟ'{>}��g�g�!А�ö��糎����=�G��r$y�Ž�0�ސ������a��h���C��A��24���Э�!D!�����2���w��F��Pa,��WH&1����5p����],�K���S�O�T,�qL�I}��&_�,'���`8�^c��
`|��G轚�p٬�C�������C�T�w���$�k�Ned�Fm!2GB�3M��3�:������3���)ߟ}�g7�y�ێ���ΘN��p
w[�`}���;���K�=�Mt�$͐{7B�ƴd.��r42<&���-g�\B��3F�V�l=���|�DV�B�ӏ�2>���g��hY|�3P+8О���F��I�����4�d�������A�
"$�s]iB��F���I���3���$tҋe��m�l�*s�����w��H]���8J�"��>��_x���	=�x�SO=w��}�]u�5����X��,$yV�'�p��L�;zC��+����n,�Ŕ� %�k^B���J�ΝI��|����dD.��s��W,Qw�$�_���M�\9��~xf!�ȁ�����QM'V �}��'�Fɇ���5��Km��TB�Ͽׂj��N��=�:��c|��5D�\F2�����~R��@��v��yX~aT��Z�}�:���K�\�8�����}ۧ�~�#߿���3ϼ{������ܢ�3�����������w��H8HF���^���I�+ݓdi:(�!¦�!��O��!�.
	9�4��|l���"�P���h������H2�G~/��"�P�]���%�B���dy�' N��V���|�
ผ�����ﴸ��Qj��4����=<�j�O�qߠ����O9�j�'���
ُ%I�To�>�VV��-=�ݘ>9����ۛ��-{��<��N�S�з}�Q�~��7�z�kʞ~���?����W����:̛Ð;d�H�i2�q�h�.T͡7��a��J�.-�CL]V�,@���ɑ,�� c��`#����c�e�^���,I��(���a(��s,��4B �k�=�kE:�m�;��t(�F�;-�p��mٕ�(N:����%d+qY$K���䁈�h�僖\�"@x^�;6X�y�F�>l�a��3A�Z[C�� I���>�m۶}��G��9���g�<�-�z��2@���N�q��:Bw'�A�7����a?z�&���,�W���݇.��iW,9�[���d`ܩe��3
-���gx�7p�I����B�ջ@|Di,_��[�Nb��M����V�.(r�$"�ED ����A�C.)����N�Z2O���,��X[�d��ǃL����
�@5D�2�A�A��ч0�o[���^d0����г4�zɶ��}��G=�ao���և�Cj���܏~�]���#@�c
!C�'���[}�/��!wI�ڐ;�Q�>�Y�p(���S��XB�ّF�T�d���7-�7���ڕЩ��8��<+��.ut�h,"�zr����W�Hb��9y����z��K�\#- �*e��U�`|juqp��s[�m�:�@�$���>���S#�H��$�I_�d���~�Ĺw��ݬ������0�k�&?#���C���������}�9K�҅�b/�{��w��U��2tX�>XtC{�DrGgùq��R�Q����c��|�1��Z��$�sǴ���!]�]�G�7F�Z�b䫑 '@��1m��ĴK+��}dΟ�l�@�2u��IW�8�Y)��K��W���S�Gm�%튓��I��'+8ЈR�C:'{�/��9qS|4���tL����/\W�}T��c)7K�>���':��S�K�  VIDATe��3͗�%ti��<�ة?�W.[�Erw�ܳ4��y����>��c�~ߤ?���x�C�]���ܢ��N{��.���]��ʷM&ӇOi�ֵ��bu�;�J,���n�#]8�V�0`���a&�\�P(n�>���T���D,�LЖ�h����A��\�EX������w��!���l}�/]�l�E �s	�R>��H � "en�-A��i߅dc����3I��5��l�j'�%���i�ɘ�;���-]��[�\#]�&҅�O�f�.��,{�x�)��',�=H�N�ҭ���j'<KA%�����LA(|1����<�ܐ����	'sv�\��w��o�	���wo���wᅟ~�%�w�u:�>�� �Ӎk��ceQU������	\G�g�E]�H�H_sv���Rsl��e�@��e�yp���{�5��_sz	1m����=Zb�ԕ��)�>��Z���e�x�{}����HE{�컯�����C���E#sM�̵�h~g���:�Y�C����ǲ���s����:�M720 B�6)e�A�N4[��D��kϚN���^B��I�x<vՁ�<�?�F��}<p~��`:;.��ܓ^r������;{����o}�[ԕ�V�����O?��.����׶��(����9��@��K��a:g��R@���8,έ|G��v7T*�q+	��m^³"Zh(j��8�$��@�gL8$(�"o���a�Ao85bE�XgHĎz�(����J+s��-�,B��$hjz��$�<M�\H���9�s���H��6-	Eh��4�sgk	�R�!��;d��h�E*	R��ydc�.�ׯ�6��͗��C���3�_��f�D�D�@�d��ƶ��`S����9>�H~.Gh�\��G��;N��ϓ���ܷm���'{ܿ�6N���uB�����'?��w����Ӣ|8߇�>uR��;�,���]]�2��#`���0p�����7�!$1p&�բd��^��5' ��ŵwőri�h�<����t�UhK3D�e��Q�H��:��	�>�qb�b�V�TXuY���-Vڈ$Hi{!��6��Hͦ%Yi���/�]�yw
 89�|�:���P� @�YD\�Z?e0!���k��_���~-h�țl�����:"~.k��V�B}��(˺6f�K��; t�!�<0�s�|X��p9K����V�#���ga��uB�bU�w����~��~���;�6�ww���zAyy2���_X��dM�7��jm��`ol�D�8�а�]0�r(�,�r"��AZ�!#`�W�'	�V�%��	\q'�r� ����9�f�t8��"�P�D��%'�|y�2��$L��\��I_Pj���OM�O��I�4��	C�m�'/M6D&�^��!ke�|dm�'���%�g��M�9�!�Rf!����D�m��Z*i���%~f�A}�6d��=��7ա#$G����E�85	�ܶv����w�pa��w��M�����߯�!w�C��~��;.�d
C�0l���S��G�).���ݐ;������q�(��Y���e�p��
W �t�X%�J��N�͹�g�9-���G�V$��!=�||��`l����.{j�$��h��l�s�����F��ۭ�>���@�`��F� [:�Ȃ��l��X�+�F#t�˖��A"B� LC��={hWK{��z/��7�С}VP*m����!\�_Ϳ%ii6"���le�<H�|Q���0��e�|��\6|���;���'�;���,�1ϸ��hG����	���p����g��<�)Oy�7-N�~�)��8�V�ܚ#���w���/|�qW^~�?M��j�;,C�@� �2��r��������u���p��VY���.���9wL͙|���k�I��Q-߇n������l�k�F�$o�_�~I��ء�6��8�k����1��l�
N��@j�-�^��W#t�{8�K�:��I
�
=/���2�	$O��	�
�\�_q���&�}�H���z��|*B��_�ݚ}KB灮��C�}P�W�!ץy�8��P;�ی\-z�6E�[XX���4'-Ry�-����y%0��aa!9���>����S�XZL.��׿�'18��e����g>s��v^��m�)l[����C�=����1�*ܶ�֢8 �z�{/n�ɔ��ZTW_j��!�!�݊R%���qNd�XL��C�"�W�,0��e�WY�!w��zf���׈G�)�I���.>�Ԉ�z/�Nb A%��v���j�e������K�V�K<H�g�.i�1�<� �o^�$h��;K_�74�>kv��������{�]S.oi+��@��ϲI9�aM9Қ�N�P�;7r�2�Bm�`pÆ5��9�����E�|8�Eq���%I�������?��Sߙ��8�S����,���9������N��‌Gc�A�8�JV���u\XUo[iNq���!CG���y����h�R��� �AZ�.�Wh݊|c@�G�|5�Ԇ�5����<2���>.��|�|ہSs���
�.��e)hm��� �$��@F�T�Z�$�e���@y-h%q�d����8�I�֦$42���}��Y��0�8�ig��n�kjF#s����C.[.w�����Y/�zp��(-���`���oӦM�q�D���=my�џ�h���x����������O}�SNޛ]�������ɕ|f���瞛��)o~�����y� ��	�`K�y�����!C%8�w��$�f�y�we`H���qb��|@�I�;9��H�9>����PaW#���L���de9���#j�)���;�5�k��>�Ω/�ǐ���,p�J����}�C���h@"��� ���܎|��~���һF@�/<��r��ur��th����Fp��9!r����M7�ܖ�@U��1mDQ�粔��t�e���%�v��q�.��a�sU)�3P�w��B���I�4�uBf:*�"��b�M�`���~�~��o���K]qw�˯9BrȑGM��{���c{yÞ��[:"v�.g�}�p�n^B0��̑9�ŎFc�0ؒ ��G�!���S:?d�ɝB���4�P��t~��`k$a9���n�9����-k͞�y��n_���rN��5�%���ʁT�C (�"\�^�[�U'�;D�ԿP��e�e��
�#���I�l�dN0�]���[������6Y?���C�[���N�������׋�[˾�3�s�Z��S
���������ǜݗ�̚3+f}�*�N
���&B߸q�K�h�-������r�ݽ��d����~�/mڴ�/y��o���;~t�)�4�����
�_��~��{h�d��~1M�������[�qA�6\�X�EO���$��1r��!B���p�GC������9Y�0���S��/�~��dS�M�ة]���Y�����AC �#]^VB�]dJ|KXu�n�mB�v���7�)Bo�y7����`�F�(��Hߔ�R�	�Ž��i������� NL�o�7<���G捽5���{c�$Oy�Os�ɳR;
錮+�{�}h��ށ�!�"{Gj���,6[Vf}��%jl��#��҆[$��.J>H�H�0��n��m��*�A�f�7��"�w���<ڸ�����V��QV���.��s'�}hm١��æ�T��YȔ�S:�� �~���ߔ�sR��=7�Ns��8N����b��a���� ���ɏrOrϏ~4.���ʤx�߾��!���_������rh>��{�<}���.�ݙHR�M-)���â�	��[��n�����Ɯ��9w�<9lc��>`\��=��5ʨ�2��ht�
:%�"ϗo E7��E_�e)��Q �09P�x�*Eܚ���v�@�vwH�.�����;�7��G�1էk��2U�j;�gj�A��$d�ʫ���NS>Oجe��o�T�5Q47'�͆�-�ڪN	��4k�b�͡BmYR���Eҿ�����i���MpG6:�Ȩہ��y�J~V�x���tb�5��P�5��=�1G�PxM/�]>R�1eD��A;Q���A#p������94�%��赩�m����t����j��j�,..&0<?���x�,�s[t���uY0��O6..${��Nv��}�ƍ�����o�x�{�|@>Z����'=i�q�p�=w��[{��Ϻ��{*�t �=�S��p	�;���o���E��6.�G�����ßŴвY>ćƎ�eq�<.��Q$��ʖ�:O��]7�P�W�
�b�L�g1��{n��I��/3lg!4�TmJ��57������	d�����������Q|��d��V%N��`�����IdP6���vQ�S}[��ϸ�	͘�TCT�w�>Ɇ��Hߐ��R,��	��l�My7�݌l�Ϻ�4�g>+�F�~h��� ˵%�49ʀ�˃�j8�ۨ�D���Sq�~((���4�Ə�� ���P��G�ڤ�a/d�ȍ���!w8����tm5�^:�F��o�Eq����{��y{-.���/|�?���j�]��N9��'<c8��x���"�?˲AQ���%��	$�S؎V�eEn%(2v�sZ��&9|^��J�H�r�Qb%�١�6�Cy:��G��-�ЛCO8���/��B��AT�ʲ�}Ca:�7w��5��b�P1u#�4+p��uX.1wQ�M�Y��["4�UIu������6��g��V��ڛ%%���:X�ڑ$л:�LRh�3�4MK�S�����qv&�*�s �T��˩�U�HMY�+YqB�	�jT�p�Ȇ��mdA�N��e�f0�ؼ��� �JgX1^�������V�pu$~={Q<-A�r(��]�x���B�N�@� �F�8�*��)`���[)r9�$�`��
Z+�l�L��#�If"�tv��ȅ�hdUfZ$eJb)�EJu���wt�)�q��G�h ��H�!V%
���(1i��$��-��L�!���zݑ�7�,�ʺ�d������#��O��H��8<���ʮs���=�N�����Nd�E؊J�BC�>���@ԋ�܂h�C�`��s�*	r���my��Av��0��t��`���<��7���G^�7��wV���Խ�	��㞺y:�}�,�s�O�=a8=�?X�8���d�gy�b�r�P"M��QY��L��L�$U��Y5q���y�$1`�F��~�	�k�m�}癙��(�Gp��!�)�r�� F����Tȁ㡮�5�R��������Wt�pq�>HiH��5u��-���:P1�C�0��%iQ�jD�w�WZ1����.���Z���M��ђGW\S`�*��Y:͒���%�HpNn�����y��^D�RY:���$��a�g�A�O܃���]�iY�.�A���.�)K�L�'I�egC0���DLlA|�U� E(�N��EQdeR�NRȔ�$�$����4c�gR�YB���}���#޲,�d�|���Fy���y�N��P�(rxR$iQ���fІIQ�E1�M��~Y���p���^ ���@HS ���_E�����(��t�Bd�d!�Ք,�p�r�T��Ρ��AGY� �$������e������z�d�bS�s�"U�o�#�]������G�2�+s����2PZd���](
� �gy��B��b�N�`K�#LWl�u���N��/� �"L9GF�C�4T�d�`g���1GZ��iw&L��-�Z���s%n���M�i�4�w�>���變��I��MCX�Yo]b��'I6X��rAf�|�iT��v6A�+B�>�\9�TO&ɞ��d�N��v�[w5�-�9f���d<N.ۺe�'ض�}�}���SNu!��,��	��w���}��G,--m[X�0�'�x\d�~�L ���j�J���qQ �W��i��$c��4D���ItE;�j+.�K�<���r\�!r���(p�����<�Kwϻ+�2���dyz��E��v�X»:8��j�d��S6�GU�]V�9���U�
m �!������w#�$Iګ2y���S���c�d:�:���hq��z��r',V���G�V�q=mD���~�K�"�{�|�O��f#�Cu��t��5(�^ j 8�1�K'�I�m:`v�kkPNh��r�t������#t�~98.s�1�C�j�_<\����|{y^� H�����B�O�~V��o����]����2��cׇb\d�d�N&�t2.��A0�Oa�V�vz�@���M࿓l2)�b:u�|��/`��e�-3v\cD�����>�9�
��w�ru5� �(� "<�d�t<�F3s�w��2P*�����ٴ0-����n$6�ƶ���:b���;�B�)B����Y���Y������A7.Pt���i?�Cu@bN8V�.�!��ZO� �U9'O(�C�8�Dq#nӂ�J0�G�t;�\�������Y@����A�!�Ǎh"��8�.�բ�M��f��@`�|BIYfER�@r:���*,�N]?]�ܳ� xR-���;N�.����S�]�w����^	A�x<YN�*��Al�^/ݰ�1���y����k��7�@�#��bqq��`pGQ�zyv�^7^�덮�����ܫ�<�K�X�{]�X���E�w�y���}��m����?�a�y��������h�ر����w׸�gO/]ZZ~�!�XZ�S�{���'=�\��N�ar�=l�0�@�,$��I2b`1�]�F��åi�Ӵȁ�9�@�(�	;�|:/L&I�=G�0���?IQ�3H���i>��aԴ?�N ڤ��h.(Ñ.0{�o��Ѥ|��E����Q�0bV}��� ���������S�b4��nԃ�AC 0vG� �laa!�����,�{��`4F�aq�b���s��e�d����s���\����?������^}׃���	�����6�K`]?�pSo|��3s�K��G>�<5���k�$��9|���wlM�G6_ïw�yg01�����$I����3��sO�$�'�m�q��!�{�7��^{��c�{�Mw�Ơ�<�6��3���t4j��Gi������֏�.x
��^	�#B8�i����F�ܿd�����f�8�@���.4�Tc�gO�g�� ]�"���L�,�%��K��k�tiX��p)�o�+��ϳ|Æl!���ݾ�0DA �\��^ W�+�
!U��J`�!�|�w�-t��{]�s��m[^�����/¿�0�E� ��K���,s��p��g��B�م$ @ P�1�A �#��{v!	�zLg� �(��]HB� b��$@� =
�g� @� �X@��t	 @�@��B�م$ @ P�1�A �#��{v!	�zLg� �(��]HB� b��$@� =
�g� @� �X@��t	 @�@��B�م$ @ � nd�G(S    IEND�B`�PK
     uK\�l��P� P� /   images/8a348e4e-00a9-420c-8c54-2da977db0968.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx��Y���u������Lwꙣ(3L��!v�<D�;H�<A��H�W���_�<0��D0���DH4�mǴI��nv�y�瞩NM���ƽw�=-��`�=�Ww�S�T���𭩆B�
*T��OE�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@/T�P�B�n�^�P�B�
�*�P�B�
�Tz�B�
*t��B�
*T�P�
*T��-�"�*T�P�[@E�*T�P�B���@��B�+_�J����Ǔ���Ӌ��j�X��x}߻�f�"�F��s� c���a:���}�c���/m��ӿx�����[�\�B�
*��"�ɀ<�;�|U�ۅ�f�]��럝���w�],������ɓ ��+�G���~�0�.o�d߷q0����x��sU�w�k[�>ԃ!�R���]�Q����]�ט��UU��&����{o~�ˏO�(T�P�B"�/~�×�<X<���������7��x�y|	d�nش�l��~;\�_��|�T���P/}�H��_�Փ���?�{���O&�϶M���ɝ����WS$�[���4��7O���A8<:
�� �]��|߭����gO��ן?}�՟�����կ��_�������B�
*�������g�O=��;?q��ٝ�j5�s|��o_}���j��s4�&��h8����m�v�����UX�7]�|:�m�]��w���w��˗_���g>�O��g?����]�-�"����7߬�v��������A۶ptx���Vk�U^Ut(��W�4[�ppx'''@�<A����װZ�-���8;���x����������/Wz�B�>��;_�b������|�n��wF��˳���S�f������s�j3��!C�j�A]#��6�+�+��BL��x4D��`>=z��p���Y�~�o�f���=z�����W^~�ѣG�|����,���pj\$��l6���c8<<��t�ȣ@o�s���������g�ެH����������'�
*T�#N$�?�����M�����������xZ9@��|t}�t�mpM��~����l�XW�P��f0��`4?D�ju�}���;~�����jx��w�����*ԋ@�#���ᤪ������z4ū�f+������`6��x2��B�$�I��m��!�h���m��:�z�������p�?�B�B�
}���w��:���e���M��$���L��L�S���
��S����eއ%:���m�Ѧ�_��W8�^�h���|�8:�W?駣O|���v��}����-�"��-i���S����0t>�pM�p}}(��j���C�n7l�w(��:�,ԣ��=Lq!��Ϛfs2��*T��G�֧�#�?�^^��]�
�-�Ϋ�r5@>;�!���xD�J0���z�<y4� ������B\���X]�ݟv�����]�h��`��s(��Am�zT���\����Xo��5Y�(��߮�:�l��wyyVH��U��:/�:Y�M�����h�h<*T��G��"G��|�6����!�P�,��P���<�g�T���2ȗ�f�����2�Н�������Z�=��z���Z�[�m6��m7-�D�c+��q�G�<�B#�C���v
����oi�A�zM�%.D:O��rG���,����ꋅ^�P�B����l\�P�2Ѐ�2P~o]S�G^�R��Xm�3OVZ�h8�[�٠�@8p5[���z�
h��
��///G�m���f(�}�(u�$�	>'a��6.2|ϋ��z@p{`���;�^�K�B�������Hq.L�������^�P��<-�.��z�l�'���7��>lQp�5��#�}���!;e��8~*�:�n����0�L�̦�,�m�u�����ȟ�[�{�@ߣ��j>V��f	�\���&"k�7� �h��?��v�蝣?��^[Ͷ^�_N�ȽP�ByjCpU�����(�+ y�R@�K"ʑ�&��9Z�p5/��X�_0�
-sBF��1lk�(���j?l��I7��Z�[�����#��_�*Z1\h�-o"�t:�d}�ޡ�˼��$?;	w��C�X���t}[o�����[��
*T�OCT���ܿUm/W��z�B��yg%:�،Ba^������P��N�)�A)\�җ��5�d�f�>���b�T�ٳ�ǫ��U�t��iyy.&�	��%�ݱ��(�3)�*
t\l���@9��I]�6��Z�<�B�
}��K_�Ώ��-�YlKnI&��:81�؈B>Z�`f�*���+��P	N��)D�����v�=tW�G�?~vtyu��i��7'�j�s�.6��-��k ��*W����z�w�y����g��v���ټ�B��*�Ѧo|#�^<	���֡��r�q|��&~�v6
t_�p0��Bc�b��?1��B�F�?@c�.<�uzJqk�����tE�d����h�Z�ܴm��C>�doς\��I�}�E.?%póz@$����۶n6�	�

*T�#Lo��W���?�����iCQ�(�kΜ����v�D�w9Pv,ȉg��	�'��0l�ۉ#����/��7��n���~���ߛV���f��LN�t:����p�?�a8�|�]����6l6k�ȃ�������z��6/um;0�8�M`	zS����6�5
o�k���1��x�v���%��s�#���P�B-z��������O�_%�S�[M�����b��Zg��.L�=�g=��s��2J\�΅��m;�.��a%�M�B��W?�}��0�P���|Y�p1�s��8נ �ZTߚ@	���t0 �n<�<��ԓg�/S�$U}����9��.>��gD���%@s"��1��x,
�;���㯽�`��/y�˿���W������/�B� *�P�B���~�t>9���COiD���g؝��P^z�B�-�^�v�ŐJl2��2G�+����6�`��m������`����_��W?��o~�?Y.�?��w���|Q�DX-�m=�^�e=�W�:�_j[���m��@�u���r�i?��RG5Ǖ�(�1� ��J�஁��z��%�]�FʫD��^�>9�O��/��������B*�L׶=����~��)tR�k�o���o.`@���ӄJjOLEϥ��~�ۂ���.�J�'-/�!' U���������w��!�u���������zT�t�8^m]���|�}��);���v���AG�G�1��uM�N�C��jR�T��Z�&x�^�5�E��9
xM>}��S�L&�~��}��PR�k���]��1���pqa�;<� �q�z����]8??��<88�������/?֞���Pg�CZ�i�~2�s���}<�hG���V?�܍ǡ�n������a7�L{�������ܓ�j�u�v��i���qgϰ����5�Z-�a�&/����~�w��sz<ñ;�ϫ�|gA_\xwr�~?;8:��qh�>��RGs�ǿ��|�����G��ؑ?�s��{��vo���Q�^}U>�����v�W�<t>T���s������>n�/}I��ʯ��.���������d��y�������OO�߿��SțG��$Z4Ν�r�$�z�����t5A>�?�Iθ(�ޡ1�|ZdX۾�f��~;9@����������}�}����j�gݤ
���BSm�ڹ��^.7���g���WS�y�m��������������)|��]���X�~�������z�	�I>� ��A$ 	2'?x�SGARԺ38�
�{�n���Y�!`y��B��5h0��99���3�#B�r�%���l�W���Y�\�����(�+��yCP��4W�!�?��NI�x�.8�3z*�H����|#x���:�� �����{�U��먔�ǿU,=��;�ߎ� ������o�(зn�u�7(�|Ʈ�$|�>�~ ����:+ܗ*^�rSX��=;:/IfO�����cI��K�k:F>�lTOx{A3��O��-Wx�Ջ@>9�{/���?���(89#��ad�����	*z=�z<�j���PR㈌��AU�a������G��mP��;�{g|4;��T�|�A��Y#�q~ӯ����ԯ��rI��-~�ɬ�53��C�2PF-Υk¦��5Txn�w�/��D�p�Mu��&����S�-+�m���=k���C�jZ�8�@�^����;4�-/�8��_�P�(aU��I�F��}����;�u|�O���N�z�&��m����w�H�|_�6mb?�W	+��7��?qrpE��~���[t���o~'ֆzw�+Qt�����U��G���P���W�C��
n�Wx���m�[��u��u_�ַ8�C>�ժ��:����M��j���i��������_�;�bq
~<��ڊ���p���j�s��a�vNUEKG��\�[��(T����c��7=����E~?�s�}��*܆��U�r�{��?��� ����$l+��<tKAdqw��F�s��s���Hy�l��݊�24���̻���d�����䝯����UuUƾrc��E�лn�F�4_^�Vwp#�W�����jyzv��f���/������G�o��懪&�-�����{�u�ɫ��d�Z�=�!xg=�K;��֖�?�Z\�2OK�&��n�pz�֛���cz��9.*�r~+�� ��I>!ϕ�<�ҩ�1����L���m�q��޿���k�u� �>�#�C����t�։���6�ڽ((�b���Ui��>]�����}�t8�W���Nc%D�E�F$
D�r�,v�=G�����XyN�|'h`?����|B�J*TA�x��{�dDz��}�4�79�g����8���9��<k���{���W_}�u^q�9�K�P�̇��X
����$�>~+I8����C�|��7Bu��� Q����	�"��,Yӭ��d=�
��_)ܑH�H��u��#哯!Q#<6�E��O>3d�Z^>�n�D�
��z.�,~�6Q�5i��]�?#Y[-mB�\(]�a�ǰ��W';�%��et)Ƴ���4i�s�_��a�q-[�E+hIk�#�����8�>(��j�RM�7������>*�08)[���n��q��Z���<>4*�@M'�,�53&z/@�w<���$��xԺC�2��80l'k8���+h�v��+lG!K7��:�7�g��B�&� {��yr8ʮ�9،&����h<�%�EOX�w۪F� �^�K��P��<���w=9����ǡ;�
kމbtуv��:�z��X�O�&�oH��Zf�\��ne5�-)����=�O�[^�{���M?���`�Q�E+�F�w�����ĉJ�O���=���϶�������탃��g����CD/�@��w�w���٧pBF�]�� M ��u�nv�k���<�6H�^�lY��h����M�>�V�S����y�)�vN#.�\��zO�*�粱��5�{L
B��1D��z���N��>Sj��vxv*�\YrA-�32��b7"�ٖ���jl>�:=s��� a":�v^}Hgᮆ�d=�/����E�R&B]/�L���ZD!���3����=x��7���^��`���G�d��F�9p�+6��0��FU���F���e5�a>�d<���l�k^�td�݈p	�d%M{Hօj�)�e�E�	��wZ��\I��.�y#�[�gQ��������u�D�sWYJ�(I��������
NY�$R��g�s�,#OT6ۆ�*�w��.R˒�!v�NUOV��h�\(�#7�U㱄Z����w�}��^,ȟ�
�&F�@R��9>����1� ɲr�^V��Y����sG>Ak�kc��}o<� G��j���0t�P������#�Y�q�~�V*�!r	���ѩ���68(h+*��C��&TϣЩ-�QiJ�Mq��iԫB�B�a{O��Z�iŞ4
T��n�O!�mHE����1�{��b����{)��+��A������u�ٿ���o��W/��_��%|H��?x���j�I|;�R�ф_di��d�B]2��
%m�s�֜!��뵳`���((�tQÍ��f�G$�7���f�׌��5��� ������q�R"����ЀdG������� j�1�}���!��q	c~Q9���yd��CT|���Pko��1a�Q������w����`���w�#*��P�V@���!o~���%Yk�Ǧ����W��7>��������/.P�w�@RH�(��v��>�k�A��iQ�p����w`2���v��BX�W�|c�K~.3��#��q~�֔./b�;ģ���#�o��
X4n��0)A��s�T����B��ŚD���>��$|;>_��X�(���~$Uҭ#7A��_���rv.���8�����OpkNjo\d+s�?�	�����x������Ǖ�64*�g�.��⊅�*;KXP>S8{��>��u�gk�� 0�,�u��C	����$c�F��LCH�3)9O��<YA�`�M �� ���l�*�9�u���W'h�Cim{y��"X�k��tэ�;�?E�(�U�0C��'���G�G���8=ιX\A� W�1�s�\O�3���ggg�y��j�������{�ᗊ@���O�i���V��6"BҤjbX��Yn�����Юo�\۲|���������� P���kD��7�ƨDX�;�1�],lf4d�8-�J���`H���ō����9��hd�"���� ) Q�C�jeֻ3�ߙv,��UI�9$��U�PT"���&/Աv����1����v�'�͙���`�gRvk	yI�=݃}Ϭ�
b��$;��<�A5��[����P na�!��X��i<��i�"����y5�-�`H�I�M�ԟB
qP�mk<'	sb���8��x�[�}�áZ�b�Qx�[�W�PH+�4�$�߬7��l�e0��6�ل��!)��`�y'�1���|��?b(�(	��%)���h�p�q���꒠�A�!�(F��E�V�Y�_� �枾'{/�G�F�2����H�ש���syO��_ 1/�~8ra�m�s�
)���5��J$Cx@�P�@i����^0+܌�*WH��P9��4+g���spK�)*�n�f�<�qV腝��
s/
��	�9_�V����m.��w���1���T�R��E�hqq��5��xc�7}��-^��v����N�XWv	�$Ax���7���c�s�ť��~��n?����-������r�ON>5����7�\]-�p�U������5�	bx��y�2�3�DY���=Z���V����v�e���hmU%��ί}�!i�f���X�&�Ͳkīm��-д�U35m�Hl ���h���w��9k�6$&�+B��V��꒠��ɬ�}F����OHw%P*������q.�WFnLm�S|��C����z:z�%ؽ/�A�j����di\G�!E�����%���D��|�zHhrvH���8���K��q����j��cZ�Ԫ�d<i�$�(��	�CT;��|�x0/ 4��%����i��������em�o�Sו��Q�k�c�U��4H}�f�Ț$Ę�z\�{"ί�Nm}�����h�'�?V�X����m}Rv ~����ޒkK� �λ]�W�(R2�D��]k;�+g�LR����P�/�(��}е���;߷�3t�>����~w[�C�1���}~;i�yQtU�3�p��0&��3M=�,|M�����1�L���q	mP�����\�{	p�2ݸf�V��E��X��z�#����A9X)�'ܳ8��i`x��F��=y�����������^H��������_ǉ}�ZoF�����ܿ��Gߊ�o�岀�ˢj�:y�����l�@l#2#��ׅ�9Ыb�X���aGK6}�m�>�O__�X%Q���VZ0!(�{:���~C�W,4S�r!��$�䙓1K�;����2������];j�-B�s��||��������,�=��G{����iɎ7K|�Q�������O$��Hf8��	�2wS�;Aڣ!�Q	���I��A���rr�t�!���˅�d"�pR8��殀Ԃ`��fzPkW!XW�T�SkTJ���A����YY Ky}=ЬY�-��P�g$��Y֑.V��]��Nr�<,s,>{qe����DD{�}��v���� �\a_~�h�O:?]�� �*A�|Ł��b麂ܹ����w�4���~�\�ʣ��	s)��(�q}B\� .
h������~<SDh��"ov�}��	��~��L�k��05Œ(O	��y�
�sj���F�-W���^֏ˌ$��uz-��+�I��<v'�c� H�e	3LqR��D����1�z�@
����;�L��
�u�L///�i�o|���7�'���)п��:����泃7�FװF�g�h~|"}�Y!O�c����
�HIA	)_#�]/٩�b0<mr�L��1!��ˋ��=��N���*	��6�t�ॕ���+Dk��Aa��:T?z�Gk܄Y��4�����$��nAM��4����PB
o�{UK�ϡM����(��������R��,�}���-e�)#����tAx���� ��8���c�ui�h�+� a�H��1$��`6�V��A����gg����!�ɝ���K/��	؊ ܭS���|>�Sw]����-�Y���W^�7^{U�+������2��&c?�)	���	�&��m��`v!�WkXmV|��'w�N���ސ��r��>Frȋ�C����9���xd�K��$Ks0k�D%���F>�ެ}��F�^K�-�/^�|�Jp�������K7Z'+����-��.�	���˚�:�-��-�r��3�1k�}�5#<Lݘ��Nֵ��g�>�!kɊ5a�*���2��N��U�Hb4����"�ƃ�^�k~Y[h+�Ӫ:��*
����P�v,EA�k6���B��6�N|���������>��*'���K;jH����w�:S�!��
`ݻ��۱�5�� �����9ʘ��1�M��y��:1�6����6��\+�[�
�<ŝ_����͇A���}�Y�a�^Z�����]��G���͚��d�Q ��W�4�X� z]�	|-�U8��N���$oF�xC��mR��炊��q�U��T@�i�↰U����m��]�|,��3������r���"j �GU��cn[�)x&��B�V�㜬���^�+:�7e+�%��׶X���a������ИeP�<�B��Y3��nV�#�1�hiI��W�%2� U;
���LH��8Wv4��.PS��huzn߈�AK�'K��US���$��^Hd1�0&x=��E<�g	�z�Q፶�5L?��� 0Jw[�V�����II`�Ms$V����ڠ ��x4b_f�{�-'U+ԓk4�;��q����� ��濍����X�r]�O�ҊAѹ�m��~b����1)"�"@�L1��bRm���d��\K���Q��c4�2$�Ý=E�d0H)�&4�Vsq�����d���A����E�@gx��j���y��.���\���E����#�������w�3�>�8�>�:Ⱦu�G.=�W�ٶ��p�9n��['��������J̉`X���m�[J��G��cd�[�C�����E`��d2���l���ûo�������=�?S��?_z!�bq�kbp�^o�+���G�I)(N![("�=H����P@����_Ù��U����>dڴ�O2�}����:�lZ2�+���j�&�:�K��f��� 6y��Kֽ��yX=g*9D�[��WKL[W�Vo���4�B�����I���A���[�݄�	.��[�4��*�����>5����o��Z���Η������}r�ɳ��#t��S���G�� ��c�a>�2�jA���&���	9<�n���H���Q�̧�:!J��Yx����:��LN�J�/!�(F�{	8#��NdJ�K���`"�$(I��q���~�Bz{���ڦ �	*-(DGj����2��]9����4=?�}���61t�7�q~~�>MR6�����{��X�	t"��gl���W�#T>�u~~��
�'�L�2o����O�u�x�S�����g��g�@4te�F�q�enA���|.|�_ݫ�/Ap���2�). G���� 9SF�������}Ze��i�����Q�����x�VW@��,Y����h������-�\���9:��r=	M�CgB���t�;7{!�/��k:�]墑���i�{Z���B���f���ݳ����nA��@��j�~ۮ稑����O�S�$J�TM9k@�r���n�XAY9~beb{������ٛ������)�O��Fa�V򕹨�Z�|�E��x.�e�{0�n[�-����rh�! Y��$+�T�$!�y$RT|��r��>���u�b�lP��1�=m�tO���:v/ce�A�&;b�9��^_�s����9ɵmc����P��9�ݵ�)]�0��ӽ�s@טL���	)�3�?�U-E��E��9���/C}.T���iT�� ����Z��hMJ ��+�e=��aE�����m��p��y*X��^k|��R`0��
0쌄����v]s�<�U�[�{������.	k�ݹ�`�>���(�/Pq���<6�&�b̄�|�^N�����V��QqgA�4�����目qtt��8�����"Q�:���KF�!�Q�u�B��SnsT�-�>����c��I�.
����r+lՔ��D{����-���2��D�]���^}*,C�]�wUts���ꂥ�d��78���p��$��T����������e�z2�"rU]���$���'�����j}����>�
Y�����P���������i'Gw`6�	BM�v�J�qZ/���s�Ь�����G������c�YM�6�<��o
D{�510Ñ4 bdr��LH�7)$�(��:=��������Vo>Ѹ7�0CU�Y�yH>h��ŏi
�n�a��+d��ݱJh��+�j�e�Lޢ��#����t��h��gS� )U��iF��@-F$U-%�<�y�ܱ�>=�A��U/2n����s���W>s�h5<U~Hh��Jx_S�P�{��U�n�� T ��R�!+�@���*��6��		-ET2��r6��i�jD�ݠ"���E09A��hHJ4�NU��5 .(�2�N�]�J0���0�����l�h�D�������XK��L�1H�r������^%��	V'A}|r,�8��j7�L�$����y�z{�q!��M�S�7R*C̷v����*���rq��=��(7Jb�	$�w��=w<�����+�;���1�(����z�As`�d� �춡����'�>rf�A
(�ڢT����\˅�{��AP��_��/f�ɐ��f�N1"���v�^m����C����E�<��n7u�;�'0'3��~p�TSY�j��U ��z{�.dU�4gU�`b�,HBâZ��Y�<P%i�)�-�%�������O�aLԇt]c9dΏ�!2�J-�}E"��..��~�ߜ�� ��� :V��ܴ��h�ʼ��|�ܬ@Ire$�N�ڶM�-�9��9���w��	�EQJ������qFq��2$���Xѯt\���.Z�t�O�>a��� 	��a�[�R���N�Q�u*�e! f��Ui��N,Q� 
s�%������^��3`EB:�.Y�,H}B�F{W�he]�?^ʁ��Ce��s:}�XQ�l[�AF�R
�� ���b��~zV��h���<n4������9I��\W��M���\�m��E@@��;r'x�?	o�x���^�o�Z��D��KV�h�//=�!I!
�!h�~&�9�~Ǉk�Q����t{
������nR�w���x:fw/|�s?II��E�85�:/�5^�@����}-�J�<e+���
��؂T{�@J�	��v�fX��`�ɜ�q�Pe�����+D9���3T@ONN����4w5�}诠�?+�u~��������9o���f[��h^j/A@�ЎT-g�$��ռ��B�o��"DI��^E_��!�5iCTG����	f��+�?��Z�S	N	z� �{�5�	w*G�Y�	r�o���j�U�+�R��*ʚt%5�[���������"w�
�GU+�*�מ����iە>
�"���M��P���Lc�;7�5ish���)>���g�+���2��>;;�?���g�gpl@��P1$����UHc!��A��\��eW�N�~m�zs�C�4�,���y@^�u���S���I�Uy%F<�Jj����d}�z>>>�X�����ݸ���kZ�%�(69�`�d�B�6S����g�
�o�#��N���VJ��jx�3�#�>M>�����^�[W8?;�ˋs���L�&�,��l��]H^��X��{��,@�n�Yַ��) ��zPu#W:��&��	�&�l�$��N(�"h�
rT��vC�(Q���s"�����k��2��vZ���;�� ��y�H��ظ�,(�V�]Գ��8j�R��{w� ��2�g�uspx���2|�ߢ�F��a

z!�ryM;b�W=ⲏ^�5�EK-(:(���BD���v�e�
*8��y-H ��sPV:����W�FI�W�y\<zo�֔a����۽q���+	�f5����ߛ"`.�|�k��ȫS<�bq�AM���"�{y�%� W$,��`�'������19[y ;�2=��˅G,�gU7���$�*��AF�N��+�:�.//�Z1�7�4�
fR�D�@�����!%���6=]�֎���Ӈ�""��#�rΚ��t:')cl�@�b+&�y��EРS�P��}���;�.�Ž��煨\�q6w����:4���J��1��$��撠qs���������\�K�E�K�T0����Hr��	:G�{Ӗ����@ښ��yEOL�5�r�ufߵ5oJ���L�
Ѿ@�hY'c%!�y~���Þ@�P�A]oʈ��d�{׭�AJ+C��)�b5��q��d�(ˌ q�������`y�t��o�E����4�M���(��;��v�],���=0��ˇ��(���v�����%�
�%��	�pJ��n4!u�%�0d=8�dA��%Vp�t5�!�xys�9��9��$���7F��	VXaŶ�J.�*D�ޝOp�u�z����*�i`������?O��煕0R��Mɾu�0)ژD$()�|}l6#e`CĲ�3,S"c.(�(9R�_61d���8c�t�����1�M�����b������1����g�؊S�DL_�[��s���}����+��Mmբ6XW�)Nk���������T8�^ɡTY�A����l�pv�>���=��+���~Az����W|�����n$J�\	���6iokF��>>�Z��K u#�'<�42�ȩ莭R��*��F���՜wY+�~���M�0+�c#�F:���ZUr���v�q�j8[���f7W�f}G!�em���
��%a͜BD'�f�7�-��!X�P*���}��}�Cz�^������w�"��!p sՉAB
(	ui�l��9z#�����qB9��v�M�f���pyWsC����Y��,}�H�;��>ơ�y�>*Ut[�=@����#�S}����
�z�Q���Gu����l��4��ݬ�j��i�&A6aPȊ�-Y��YKc<��� $?��Mp�Ң�f�u���2�0	]�.5C���yXS���Az �� C%�ƾR𜆽g��߉hG�p�V�j��K��������T''�1������Tp�-=��jc�ACS�@��d<a�[�\�Q�&eOw�����ک�wsPc�<����j�e���7Nn�,R�:��PKk޶�p0ƽs�v ����<U zX���u,A�� Z�T�\iͥ�p����C\->�Ql$�Jx#�L�<O�'A{0; )Q,���̢�� :�g��h�x:����;6@�כ5\��!X��)��ocO�e:�3�e4�А����E�Qt P���MO�[U��B��0�����vS�L�����Y���ږ�\�Ц����p|tR=/�(Y�dV;��
f�P�d��#$���|��τO*��6Н�5���R���*�ᑫ�7��.d^tu�������`R�!5�hO�d��N� q#�~�bt���q���J���A��H�}B�$%λ�#봂�_~f��G�p0
�b��(�����~U}�������~���[�^��`rt�ёnB��]�L]�B�Y���5.��ԝ
c��ԟ�A���獁�I+	I����T:�s���BB��e�P�$T9ˋ%���H�͡7���>0��
إ�
����7m�����R���(G��-t�T_����haGC�1�$DC`�>�W,���J��5��3��I��0�,�:�:�!*�X����͐��t�T�Ҭ����|8�KV��x���zڹ5�3;�}F�Rc�8b}f���9,�ߑ�z�6���������vcfU�9��>g1�aĒ��+ZO�:�I�Zc-(����(���2,���l�v�+S�����Trנ�]r�QTM�����2L<!"u�r]{�h���$G��,}�;��0�ԇ�!."��A���rki|�"%���{��ZPaZ�IyH�yA�}���k݌����R4�R��[6:�%A�b*S"EHnro�[N���9M�e�c�6�j��D�θ����j�Y?���8���j�T�{�@%`�ԑ7��3��orW4�Tx�W^A�u@��*�E��(�����u�/u��4��_F]RO��:�Խ��d�f�0��U8�6!��HZE�*D�T�� A@�ocJ���̟bu�o�f����>i���j%1�2)��,���r��P���Z�]l�j�ƈ+�w��g�5ߜd���n���?b,���Jv\����Ӳ�y�q�`�`6+B#�Ɩs��/Z��0®f�]__s�.Rh^�uV̷lPjP�85yIds�p�� V�����Vă�Mw�}�n�cSj?e�l>�fM��@�l�(	�����Yiъ6�A�g���������5|�Ztq`���M���iu3�J�$j]�E7m�,�IK�	t��!}�F�b3�TS��oS�^+�ݹNK�J���A���B����1S{F�U`s!��b`M�L �Zl�'v�3D�nm�Ǹ�
hˁ�wqqO�>��OJ��Vs>�S�I��(h�j'��b�VK�����x��R�V+I���,�'�iQ�״�E�����`�S�q:iqWq�zՠ+\�sp���Q��[	p�B/�Y�Z��X�ڦ��D�ZpmTf#Z Jg\8����r$��$�gwP�[�R�s�.��g([���;{s�뻮�lFqNM������{���g�/m.���d>��x
�h����M���X��&������s�>��ʫ0���}�?|�]خ��	-��k�$�$�E���վ��"��	�%��>�e4��bc&)��f	I��5�{����X�Ӧ}�����!m:��2r49��𽙰�b>�ux���i��?H��P��XB��Qi�5~�޽{��A�1Cq#X����L�d����De��g'���j���dc&�A�(w�ŝS!,~�C��
ȡ�L4����zV��������,\��`G�"-�o����|�w�1��D�`� ��S�>aAzFQx��B䓽C��3��@0E�9��G��:B��]HP�u���2�T�]˷�H�pe����+�JEu��H�<k�"���2��ɲ��?�|��I0iV�������������d����t�U���CJ&�����ײ��}�WNn�q5�K̄`��'�?D�^��h��v�@5�\���s:k����b��A��7t	��d
�?��rύ��o����J�$��&C��"~�`/�pԢB�X���Gt�K����>4��Th0���v� C;��X��}Lk�Q��r ��V��O����$<ڬ����G��A�C�m�*����u�T�u�&�Q�<�?�fu��pza:,6u����=u��k������chqQlqQ�7�y��K��G�(�����	�f0�N�}$i��<��{���c|�B|}��������h�^�\܀B�}Ҍ�3���jѴ�dA;��(2r8�����r��O�30��=�����!��t����
����VbsQ�2�@r<�,&��[L�|��g�@��h���5d�J6<��&���q�\��`&2�{�;�^�ҷ�bbl��k��kM[��)ǛA>>v?�����:7e�cQ�Y+�e(L�h�\�v]a�^!3��	������v���۽�X6�sH4bIt���g����!A�yJQ\A,j*�V� �Lg��+.(� 0�@_���9$������C�,�#�/�R7�ɮ����#d�q=�R�1+�k�t���u�7�	*`#���L��h��˔����Nc$re��C�b)݌�H�C�k\:5zX�R�kq���.�k��1Z���̇ݱ���������>_��'�����!��*E<�Ne��g��Br�2� �p*�Xt����%ֽbQ������J��%�����;��������x*g�?�/�,�k48�S�"������.p<���x��A�OtqI�"m�EJJ�ד��
������#�g��7��"p���ְ���5.�-5�wR��sҬ~�o�U}������W�BE���"����~�x������=A[�(8M�����+��ˁY P�MLZ����A�W ]�6�L<��>�����)��qt���C���0'K�	*l�����r��J���> :�����܂�g~���!B�V0G|�Ҵb$ֆ��W���Q�)]M�7�C&��u]*��y����TṬ�
ͧ�r���gH�H|��-�`.���W�\���r�mߟ��$�r+ǄTʿ߳� ����wM2ȶ�s��E�cnr��pxnn���>2��5�F8�[�1S6R��\��V�3P&�?��uVf�X���ۇvw����8��歿{�ȋ�,V���|�q��
�|U�}�veC�՛K"��Oh��m����Q���`}�;�j����탴�ew�?�ew]����|���@�iM�cb ��H�=f�z�zIH֮�n���k���C$�,��l2�C*���<Bz��o�Ͻx�mhА�q�����UCvP&�!֘c��)f�@�����$$�5W}3@K��_S[�ɘ�]��F�P�Z^0�q��3�-��]Bh�p0��������~�F�V��N44/3F(�t�z��������^����E��(������]�_|�ly}�����W`��+�j,�-lH����ɛp����S��f0�v�R���8���F���EF}}�v�m(��_)�Բh� ~�9�n.�<kIo !g/�����������ܽs�0y������AN�J��(��(�~kc>�u�+@w��M�����@�Ub4�g8R�o�VA]��8�yf�,�D�1�W�	E���-���..��K��x��)*ed����Ę��UC<�1���h>��U��Ӭ�u.�s�S�$�+L6�i�A�9ϛ� �Ϝ��cMyH����!wPxz��X��4F_C6�����+�9a��aێ�z��)c����{���4ʞS�j
.�x4H:O��ڕ)�9�a��,�u\���;
��>��a��	�|/�ř"�|�$'��D.�͊�5�������iQ��|��>*�t���%�@j��8
A'�n�h�мY�9jA�>���5n.�-���SønI!�׮����Ǫ��}�{��gH�=L@�N+.wNN��0F��E�8�5I�zsy	��߀����w�����dz���]��:�"w)�t���v�<r@�BF�il
���ھC����g�{
$����
����
����]�Sd�O�~��ȇ�a����+n���������(��N�;|��o�7�x��Z(>����a�N���␺)�6w:���8Y^49/��b������%<F�C���d��J���߁gO����1. ��&0����
i�Lk�hE+�w�m�;��l�s�j#�F��|�V-g^H����1�g�9Бx/��z�`_>Y���j�/�|/��A!!�|�k�qs���ٳ�o�'���L�>�����Sqx�X�f�H���ҋ�ʰ���:)�iAM�hh����A�����1	�g,�?��7�h�%!@����z|*S�����c��X��܅~g�v�1��h� e�����o(I􋛡z=��1ϣ2I8��2�ivh��\Tf�pm{�q4	��}�z�/ݧ�K���"��Ԃ�����-�� �%�
$�Q�E�s���kOs��(����7%���C;�՜���֐���B���@�9g��G�3 "T���z�<Q�5��9x�y�^��y�2��=��M�ʟ!�_�j���2I�����12����N/O!�>E�����?��Ω$0�9X�`�;.~�
�� �������~���FCb�0�N�,��u�pM��x.��R�\,��廬��%<�.�|�W]߃Y��F�h22�~����g?ː�Ƴ�����ΰo����c�F��//]��y:��#�jOP!=]-���lz�c.�O�pK��ׇ�N%a�{�]�!��ރ{pr|�ݱ�B-qF��6a��mj��y�(��hI��0
w�\��V�ìCcrVZ�FI�<m�A-�T
�)�Z��W�kx��)<z�>|�j����+#R盚QV���KK����C�+��<@+1��1'�r�RW&R.5}�r}��/����r�7�a� �v��r�ؠo4�<���ҹs玦��
y�P�B�璑qkH�) #U�$[
���M�5Y���׮��A�v�w]�7�d�����4��Q,���l��	/ê�}�=��%��!I�N��;6qQ���D�T�8�3h"#e+2��N������Y\���*��ߵ�4��`M��L�s��3� �����e q2�6��,J�YɹF���`4��qu�[AC�"�+�c�ȩ�Qj��7DO��۾L���Z"�^�I��u{pu2�*p;ֺ(ZB��/�@�Vu�g��o*��� �
�d���=�+�4�t��)Pe���߂����R��"�[^���6��z�/�c|�<N:��VQs"����2!�Иq#ᱝ�4>Tj�W�Ɲ�(�;�Ƹ�a��}R�x,��%<[]���
��
�3�P\4"��4}�C��K������4m�(2��1Pf�hD5��p@�|����?��|�������֟�jh���[D�mySv �\���B�;B����'���;�!.ܮ�Ț=6�k�-i�|e�ڷ	u��ƍd�������}�6���Cc���ݻ�>6	��ַ�	o���p�V�z����t�;w�qǸ��k*�/����Q�z.��Yw�T���Ƅ�[А��������׻+ЅaȆ���hvJ##�"����)��XC��q��2�d$A�WP�o�h�&tB����G��'i��a'�+���� >�������K�f�����i-��ܮf]E��&@E�殎 �"�ҺLɐ���>{x1#�)��B^3e���B�5��`��{MM��,��A���X7��Á����M*�C�@8��K��4]J�r�
e9�Y3g�=cr7Hn�� �(�|DA�_�pם����I.!V$7t��%�9G��#�.n")�3�򼍦���J�Ѓ���d����=Ӱ��dI��RO�U��k��)�D\T!�b-��i��{`�Q�[�.G^,�޹�>��CvbH@�$�������С�2;��@F�7��=h�u0��yWh���Ar��x�)>ㄔ��
�E�s�|��g3iYK�>?�轵�'��N�ߺ%����/j�A����ף��'�A�r������/���)	�W_y��]��@������:�E�����f7���D/�@�\]#{	ǣa7p#���=_�Ы?��%$����Q@?;=��P��s�WLG�:1@�k��7�3�(����P7���vڰ���ơ�&%�`7������q<}b�m:����'���n]d�B���F�a6���K�l�;���s`KX-4k��K���q)xk?�žkV�h�	�Y�bB�=��N�@�:��ᑸ'��!���W��%AG��@�	����+�4bPf��@�<xb&DV�D.ׂU�J�p����T(����֤��9`i�BT�B|6��e�U
̂��Mk�,��,SV�U�?A�0j�
��=�XO:�R�#�7ϩ����M��0lVPb��< *��?���wE�����״|�xOQ�[d�ܿ��|$mɐ�L	܇�Sc{���{���A�!I�%�M����I����\76���)��ǎi	J�7hO�~��s�;����)�<�ԩ���n0��+�u�>�;G;�Vwz�����?_ЉϏ{n��Y1<;?���%TC���}0EſF���7��
��.�c�@G��rz�I�v�:��������h(�	_��E�?]��ԣ�GC��C|��pL�=,�g_�W����gx~����*��R1���D�M��8P�	� ���E�lZ,��Z�(�Q�����е�NPE몓:��^�"��8��,�.`}�`_�J��NS@Z��I\R�d��/�n��[��K+�����	��ޙ�؋e�`kQI+��㌹�B�e!v!��boS�
��5E�����(p�4N�����g7,7K��|h�;m�ԥ����eHɂ�ғw���k�P�w�Z��2Q�2ulu��ȵ2M�;�L¼� �*c~�0��+]�ѣ���H���89�:2~kW)p�����$�*�����JaeUH"��Xa��u�C�&�s��q�@�ӎ���a��Kmxmlr
z>1�SJX�g0��_����X@����up��K�	䞒�b�kh]XK��lyT�[�?��
��~�I�f��(�uqg	�w.3�I,WH���K�׆5-��:�'��Gv,��:�trP�Zǹ�>W��w`.^�в�c���J뜔���W�27aK�El�vRlH,��c�]��~���ɯ.Ϻ����sg$����b,�yҊ�k����ax�a����B��z�W:�#��
�C4���s��TJ���� oܠp߶kv��Z횾�T2	�Q������L�O��=;G������<��)��ިHA;���5ϻ=� gbHP�:�⧸ꏝ�w�Y������	���P�52�p׸�7�(�T:�f�q<�!�3d�wa���GO`}��I�@�|9��Vz�����aضIZ'�\�`���Ah�q.���+��(½�&#N����:�𽵆$�Pz��nNg�
[�E�
f���@4o6h�(a.X���-L,V8d_��2D30e��Ʀ}���<�+1#Gbt��_{�5.���JV�L-���9?�l6aK�����ӱ�(w!Q�)�{ǾR�I��|���<=��������?<:��FBSP#S��H�DX�8�r� ,�#4m��`��5#�2bEC,,c0�����p�p��:��#v�X1iN�^m��dA�6�Mq`�m�kc�",][D:�Li����0;V �7NJ0�@���񊊞�n���5�`�Wzh�Ke^+���Q��F�ya�88��X��5I��z`��TF&h8��EI� @�]�e�[�vkiKksqu�ֲ iW�@��N�}j�<b���S�E��T�B4��|.��SJ*!}\�M���)���Ny/��-%�Uj���u�`%����.?�}�?Ҹ����`��(}RR����k�Ed��8B0�/��
�uB�W		cX��@#�2V�!�����[�p;���&;���ض��B�!�&@]Gns�
�a��|��\��|R�I���sĻ������,�S���\��ͭz�\_��[uza�
w
j^�h<s��V����Y	i���.M�R�5?�@7� ���LߡM���x��xH+���v-�/����`��4"x�^c.�1,��(o9u��I�����>��������	�f+�G���kN�r���
��ꌑ崫�k"�jj�Z�i��b�N�mA���-͐�EMu�ɂOF�O=�S�Y�S�!]�
z�Z����}��Wka��x)���RPA��0�(Cꀕϋ���}�vߍ���)T��g�p�e��q��(��X�>pfD��	,-�bk)q�ԩl�W���>��ٳJ ��31����>��[��>�!}�R�8ݥb,�b��8��`~g9bf�a%Xl�>u�=��|��g�s�\d��O��O\W�k9@ʣ�z��%ő�y)�ƹk�gHK��ཱི`EE�@�\^����2:��"ZBh�4�Ƀ�:$�V���5�%O��\2I@{���iO�+�{��E�⹜8�I<���R^L��� ��Pp�VF��
�6m`�d�y퀻��{�Ƙ\��~Z�,���ʭ���Ip���Eh4�]���Js���Ct�јS��͕����Ha�}���(<>����?�~�����ӯ~�;���#�xK]�h���A��q:�h�:���Z,� �6M&1��5 ����IN.-�J��ĺ�X�����yh��m
H�Δ�Ԋ�`_��*e��j�rE*�RFy��ٔ����P?��)�����e7aըe�n��<�ѪRQ�1-�LA��1�\�M!��eA�Akis���LG�A��n�8c�.YR��)���!W��F+֡�`�^�a��r�U���g�L��P��`�����G���3�- A�xޣ�.zcAP�֛Y��M�ύ�[��<� B��#Y/����BD��}4&�
6b V��r��^��?)�ꤶw
�SL���g�K��إ,�1H��İ�x�i�mk=�SIa�Jn�Q�R1q�,�l��u)J��B]k7��k�ǆ!�mb�dkfb�r}�����'����"�)Fc<�je7��p��@��^Ж��<)�����4^T_a�Z�6��"*�0Q �����<�Т}H)S��vA��	�3��>��Y�7��9;?���,B��Z��-A����=�7jSŅ �yTTw\"�C�͕0��!�Γ+�$���܂��V[]Ԋ}���^�K̩���Wy���=�YZ�lN��[r'p�[u��� ���T��n �۴�h�јǒ�F�F(�p�s��No|O�w��I�T)��КFѽ����N�9(�������X��^�>tg?�>9����7���}d8�Q ����*"Z��=/���tJ[����6|P�`6�qԣ�����(~p[�.����E�R�o����X����疎�mZA~�"�h�lT����5uLg�0Y�h=8���c��GC)��
F��v�[]�h�1,y/�$\��������h�#�A��*����F��ag0t����!
��G���8E���ܻ�����0�?������q�,$��*Eܚ��y��0��H��|v���՗_cF�R�ҊlPR%�!1����>�����	Y���~C��sTN��J^�T������9�R���#Ȍ�6\���RM��p �O9	D���+M�<�FS�hX	N�n�M�i5�GBI�3�80�]ip������wQ^5��G%�<�*\5M[�n�Fs�+^���Պ�H
'�^
Ό�3~>����&܉��C�[.��4����9�����p�x��P$���4�	q9Y�
��)z!ʜ(^$H�����%?�ݓ;܌c2�De�ζ���|�J��Ʋ���WaN�|oV�<H1�s\Wۃ�ܿw�?�5/x>U9"�S��éU���{]�]񸹘�ʛ�N*�\Od�D`���1[�F�6L���-�4o���=Geg�Z@{��f�Ǽ�m��'A�M��E9�0�, ��;
����lu�@��ތ�`([�񷊃6+1���� ��2�$����F^�sA��2�J��U�Zǅop�!T�NN�<|4�K�1�!���~�S���΀�Ϣ�7�b��9p���4̞R�̟�I���DTq��`��;�t˹� U�B�-+E��5P�*PiCK�	�^������%����:0K�؉X��B��ϩ�VU֭,L:A���07��B��^��9˧��%و=߳՛�Ԛ !c�K�֣���2�oQ��+����h<�8g
Rh�R�(2�����k��<;�V�d�D�Z>��!H�S��D�u0�9&姝����5�! ���w�G�Z
�	2?:M%5����xc�;ݾ�� \�Y��I(������3kp"�	�;�

a��,y���0>����&#!�Y:���aZ�V�%v/�[�YU�	P<�`'���V�T螬D���B�ݶ ��a�d�l���I����R�
`/��.+��o}�Y
8�9����b�J/��A��S�FjiL�I�i\X�VdK1,E�t�н[�2�)�ηMtm�3/�㾰�pD)1��x�/��Y8G�E./27���<0�;��P���5m?i��=�����Q):@%�˯.G����^w����ڞ'��G7)C�溰�}:"H᫠h�e��Z��d�TZT�n�E�� !��Hv���ϡ�/�0���K�%YzvNĽ73+���z��ٜ��4�4ðׂ�l��d��镡�v�b��x���,����B~����fk������ʼy�8�����N�ͪ�Y�OwVތq�<���<&��օ�f�<�7>�����G���'�o����ʯ������o����Knw����o�n��{v��������z>;�G9wחL܈��]��F��>��m��fB5:4$�m�۴� *ȶ6(AVIm��p�k�N��O���oO$#�Vv$ķ�z)W��ZT���91/Ԝ	��Yc}��Ɠ��2}Gj˫+0��k�s5&��x<A�p�Et�J�C���'�`.v6eX`�&F����˻ с!��%m�B"��C6�����%��B�ّH&��t��)����wr��ۅX�~2�C^����x�H|�Fh�Ε�AҧW߃zr4�'���SQ��a$!jm���;i����}��CkE��7�f��l�NS�O0	�Ca��,���#��G�f��U�JB"���%t�K�4ӠJ�p@��S�%�T��4�X�j�G�Q&U:Iɫ`*�src�)��32J��GMvU��3z�9U�J�D�PK�"��΁)�K�Y/h�8U2Ò���[�Ic��n
�Zˏ3��J�T�+��|'Ђ����)�bg��E����R�V5/����74P+�k��e��HR����%�i�DИ���:Iq�!��AU�~&�˲V�ʬ)��y88]2���7_x[�-�}��y�M���ZӺ��Iү��{|�9?A��.&G����Ua[���L��?���'}�?��n��v��������_��o=�������y����y���G_}�����_?��[��2� 13 ��������!�CC�WZENdT�l�ޣ�JM��M�� ��6*���MP�H�'��,���K�E:uޡ{8]l"M�'.ae�U��ݻ`3́8CJ��e���V�K��l�V���8�U� s���`ebI�LN?�t���'y]�ͦ��q�:��a}��nG�X��$6�ڈ�Mv!&8��M\q��;#q"��k>t��g�Yo,9M�_�^!�K�5pZ��&�2���~�TYW���Č�6H�_�f�V�G�X7�FP6kG��=�Ҿ7&�
#R��%,q0��SB��,�=<��ʒ�c%���|�N&H��ƺ?�1b�8q~E�� �x;ˀ�uS�F\�w�{�����[j��8�@�!2��2!��E�[��t�!ǲ��iWQ�W"C�lD?��?\�LW��+0�p�Le��v�{��Ӊi�a�љ��v��[m�yK	O�a�V���	���<&E 
�^`�9�f����\�Jg�2���/��~�_ⵦr�?��?�4˃�3<L�w=b�4e���8�*�FkF�-̐��}~=�>$$��)e/��p��m���̴jb.A�pؙ�(3��h����U�����3�Y�S��Ob���6��F�B�OSg��C4t�����u'�`F
p]Nc?}����]��������:���Kjw���������v��_�|C��{�CH�s��i��Z��
�q�N�ZE����ʒ���}D�c�I8�^]� >`�+&@U
�ի �M2ӓ����S�-��P9�#��_k?�2U�l�T���ZI�1p�m��0�*�INtY��ƲZI69��Z8kx�LBZZ�YC{X�0 -g2�5:d�k�W=T�q�A�A�X�
�9�G�Rr),�EӜ�|���a$�hQ�s��g�}nC���T��o;���Ҵ9�˽��4"�-0R���`��û���͂�^�r�wd0�hp��ؠ�wK��~����՚�wb��l	��!�M���V8�K�@f � %{�S�z�ï�����M�Y?s�b��>� �[�Q����i���r���z�E �c�G���3���ԖUJ:/���5g�E� |��0�'�Cě5P��<�y&�h;	�ݣ�a�U,��ۓT,kqPܠƖ�`b(�Ns�y���њ�7�� ������8���j�D/gj�ɹ����W��V��1��k&�E���'	�s͌��/zp���J��tvu���ŋ�������fs���Klw������!���;�/h�ɑ� NTjו}i��+�z�R���g����v�ic��>�>]wYG I
�S����]J8B:\�zC<^�k�H����D�ݳ���=w��$KR=#7�5�Y���U��9��'�|�uJJ �0:���̞�*�9���0�
;ס@��P�F�&�ΐ��߃;<1G�v*�U��尳S���S�3[5s"bD�ƙ��ώbee�<����l��|Wl�ܳcq肄L��JMJO��#d4 w��5{X��}>VDK�WնIײFPɦT�U�綫�Y�R����`��K���=����{1��:0�1��"��z�JNd"�z�s0efW�VtE���{�٬�R���
R<c�Z;f�v�H(&,h8�kI�t'ĕq�U��+)���Ņ��]G*�{�u�4c;N�|H�N�T�Q<�9�:M�[bj�3�)�eL�y�� ���ƚ�s��~Y��&��ga5I�_I&)����f+bJ�y>��[�3���E4����α��U�	�?}�$'���(�i_wʄi�U�á4��UF�I"�a�4�݁+�q��i�!��A���q�LfI�E�Qpf���
�I����'Gf*����w~���71:'�Klw������U�z~vz��b�~��ηNv���%��4�F� y�����=�=�&{�(Q���.&.��Kr���[����A��:�T�e��PdD��p�ȁCu&ΰU;>�-]%�"!v##�"dOP�6��=>X��T����R@��%Π�x�Hd]��T*){h����w����)��{�B%���g�ʘ��H!pqJK*ayL4�ߡ���^��kLs��VƯȞ4B,yc���h:FMN��^���T�}�!/�i�	���ptD�R�������L`�LSMl��}�5����{��n+���9':��j�ǡ�*�B���|FƘ�>%b�q_��9U�?� ʘxܴ׵����v��-�D�{Ee}n��<�g��'f���8
�ջRg�y59
o��� &��>�wlǇ�K����R��x�j�m�)��6ɿ�օ�[.z�=��W/�����,�N��ȀN(D�YH">Q�=��'K���N�LuD���3(w@k�a����w��h�D��_"�ѣw�XAMN�3S#�hLeMw'䋱Q��F��H�8'�w�N�b!�@0 �"���$9lr����5!�V#�y�l,|#�@+�	����Q	��;�6�"�:���1u�h)u]8)�%�dy��?K�_<��ŋoM�}�	g�,A����������o��?�÷_�|yJ6��C�2�\`��CNj$��E��(
3z�� ��?����ιXBƔ��)<��X�OF�t���ѡ��_�=��1T5��P��eHZ,�jG�л�"�� m��v}Ԛݳ�~���>HcHOTYC'�/��Dĝ����h58����RlU"uɁ�Z�&��z\�)���ͰVe�RP��Z}�d��C<d�Jch�~	�`�F�.8́��^@�-1�[�6j�Q���q�r/�(yaM�	�� �W�2�xE��Κ��I]��amH295+����!s���Xߘ8�b�O1vvO	����F<R���B�ux��{M���Ex"6�� 	�>�M �uP@jDp�yt�{��{ghw�.I�^�7{ᓃ������b��㞩�P�f)�!q�Z��8�p���^s��:�?��$��K&�C+	���� �/�Ta��)m�H�,"��,����H8�?�P�^P
hܳS�����B�hJ��}^���j��$?�h�!�G�?� � ���YQ<8^�&�����Yq>i�X�ʉ��p�^#PN�I�֑��ϟ�L��`u�]8�������w�J���Ę}��_��;����W|����R���,A�������>�����鬈pw��D�F�I��B��^z��KS��z��3.�A�^�u��AĜ��9~�=p��ٳ/��Q�d������~���_�IB��]'$v�`WCKJ��L�]n0��V�U������ա�V����OH�*�j��;P�*��!�E��ա��p]g~�����˕v�	̒Z-�M��.I�����7�!BD�fyr�lH?�|��$����ūc��NM@0R��5��T$�'�1��K��A�Ӄ1��6;f<I��p����A:RhN�X3cI� b��?�UH���ۭ�#u<�X�nN[��i9<��J4a�I�"g��3�Gߓ�LJ�ϊ8����
#�5���
l3t~�jG�48�1��� ��J:GA9Y��%-bipz�ph��8�}�R�Wv/	�4�*]v��3��byz)��f&�1U��P��hh�8�s�yc����:D����;1�f7{'���%$V�L����l��$;���ڴo"�G[_��_�0��3 	�$�k����8�Af'D�b�?�5�QO�w�~O��z�L���֜s
tb
`?�$1��ߝc��)�?�Z�?Dw�eX<!������Ge���6������s�������O� t��ά��ɴ����w����oҗ�~g	�G=��`�~��:#`$bMI�	>~��qVO�|�>��Sq�X�,�0m��|����A������O>L���*�����k���hH�M���O�S�~l�]I�D�x���w�L�82�'��$x����A�22�?�"{��p�s��%��:���$���-?����b9��`�-�ۙ�g[�^�cb+c_r� �rA΄�!c�y;��YԾ;�RI;d��t�)�?��G�Ѥ��<���&T��lN�U_����ټ#��SN�+��F�|&��Fj^"�}/^�ð�=㴸�L���<�I�+9+a�:NZ%�D��+����������R����h�������H���[T��O�:� ��l��l@��`�ɧ��2����ѻ�׀��$�hQ���S��i}7�|n�t��6R2��$������Ms�쀹-����z>�/1�!�p���z�7fp�J"�:S��`S�Ƌ;I���d��sG��ȏ�+&0�qr��BD��J���3�D�Ɔ�~v#L���$w9G�^�������L�vNE�R�}B�
��N���5�;�h$���7ߌ�$���[�z�^W�0�1	P�_�\L��'��o"�ߺ���\��,'�y6����l�&���K�g�<�jG�]v�dF8Ot�����'���?O��LĚ��/���dV�䓏':����G́��{������z���xs�x�җ��,A��'��y��~5II��+qA�����A5F�Pnoj����"QHΞ� ��[ B8I^��HHF҄�ᄳU�)%��P�^ǵ7j���E4�MjP�f��\F8��o�������;z�K�8���~�e'��E	eѱusB�yP�5�u\�?�JY� �� �tə�D����9��b�TdD)DU3��DT���L$���ԩ�^G��[������Z9L��K���:p��!'&��
.2�p3��؜��+_a�f�H�6�7=O}bBX������^:c�C����~r�Aq���~Dx�Ѣ�u���5����Y�vqf�K�����x����Jc.ӣG_IW���S�z�j/U�-&��*N9,�_W�3��G7�D�G�p;�	lB��	D�0KfC��.��ىW�p�B��  �!�G���%9�p 3Q7{��Γ8k8���@�E�O��^�e6l&�ꠉ$A�Na&jt�W6��euK�����P��M�c_}�C��ӹ�к��@{;���8�	(�ăI $"L�%�xԋ	~>��3�:K�A����//�~�M��?bG7b��c~�س��ku�s΄�+���>�����O��/���j��ڝ%�WW�nB>=9�\k�q:[��*(~ �T�H��Y��Dd&��	-��KN��+r�:�&�$`N��v�8?��SS�iB�j��'�?��`��wv6u9��~�����Sq��KL}+�C,���vD��H@��*�����>7ɸ�gT�E�����Ԕ�}�o��Cd��RXk��=�SE�����!��?^�g���z���G��*It?0z�6�p6BFDĠrGX������	:.�|�U����0�ڊ�r��o��XCB��:}���c3)0A�"Ҥf�>�o"��9��LwE�S�h��D����F�T���-YcҀA���
��֔D3iZ�{�d/�y��W��-�T\H<�8�Ǝ�,���A�2� ���zM�ٯ9�%h�6 L�����8���>��@y�b� ��x.\C�x p�M�'�z�wv�1����2��}��b��ʋ�$�'�1,x>:l"�dݯ*%_�����%i$NON��g����\|�k_����$-����0��6~Ҍ�GFz)%�Y�$̐RM?�`��D���c�詄̟���P��\]=g�Α��~y��i1� ��]��`����X7_|��[/V/�/��Y�>q=7�'��8�.�Ihq� �����B �EG,��pR��85�J*��ǬjJ `�3!�ˁ�� UR��Gd�����>9�x�N���J�ׂ�\��vck�0N�#�q�3��e,`~0&'�x�%����'��R�Ι*�!Nz�ݯ���y��4k��H���%�\#(8.�)6'�sG<y/�<
@�P�t����p5<�*M�O�q�}�!_G�W0������״et��o��Mz7�ML-d�3���5?��cc`ӎ?�<a5�6̹��55ʜ'@�ީϏ>�H5bo�y��=�1��O�����UƲg�5dٓ
a�22W�߄�	��1���Trt%�+~
7�&&ƼG��!ar�<�7�C g�l_�a�js��9��1<3
��]���Τ��w�Lk|�>_����낢��i���T�;�^��ұ�"Rޣ�`cIZ���n-:����^�'�T~8�����$>g�8L�:�T����)7ZPK2�uZ�"Q>��C5�G|0܁��K\J�`Z����'�ɉn �n1�-oL�^<M7����$J���e���W��:=;��v�P��}B�i�wE_� O٬��w�}R�$��N0#l��%7��Vzv#�è�䄱V���(=c���*�du�)Z�%V~^b9q�;2&9��|����r�?�Z�����(�h��i�����!%�e�U���p�{��8�̞��PϷ�K�x֑^i�B{0�rx�E/%��>���D�	�����5(��a���kN^ŝY��Y#��ܱfd��f$~Q	7!���9�ٛ���/�C��v��x���Fd$�"�f��u)#���zP$K��qu݉����E6v$�T�0(;�sXL��ڭ:b�X����;J�������CZj,?g$�L_�Wvl�7�w�\@�糃�b*Ue<BEϴ��r�}���_��	p�Z��+���>]�5�D�8s�`��y&�5;�:��z�c���6�0���a�n(*��X("ΠIp�Y�I�T	�E�ըN�BK6{ܐPT<��W7�u���>t5�y���tj9���Ԓg�Ǝ�����<���:!��l*�)37�6��J/P��1Bb8��B��*aDT';�<�@�WQ���"6M�z0�g���p��E��Y��ޥ�~:k�w�h,���-e��a�^$����a@N�f�ZҐ�B�~��h����å��z�0��"�6�j��&2�26k���! U�T�����sd1���S��s 6��$%	��+�ƞ%O>��W������AQ/�!R�g*���^47���e	tz�j����ך�d2a�~nkޗ3�Ǝ�4�G�� �F��/5o�(Ge�5`"&�Y�=��#�+�aF
�~n�{J=�����x�
 ~Uвs��6�i�S����g]`ïI�QgC%�>��9k�������GeJ�<s����&۸J�Q�}7�udo��e���V���ujo�%�smSE��L�
k��DC�Ʋ�x�w$X��͵�Wq��Vu�å��䇴%>Q���<a����^]��2,��VIՈy s%$|�E��y��0�]���F�u�& �E%yG�h^x�9:�+C�� ���ZN�r���nTr��%/�{���p�a���+&�!�����a�_�W�d
��<�u�I2`gG�T�."x���׷+�L�{Ep�o��3������d�5̚�yW1"���.V�T����h��_5/Q��K�(��z8R*�ʪ��5u��a�qP�Y�k0��<N>�G�Ĩ{:���b�Y�1��U��S���9��9#`���L�&-�Ou��b��؛�,�B� �x�J��s
/.J���x����`(
̊�0��5B��k5����5 �vgtFEs��NYr��Z�.I���.ء�������Djx75���x\�n4�	6��53�w���멂�
ڝ%��&ZQ$[1T�q���*��󒭏,�Ϧ���RB/�4Uo����tY�n�2����]W�*��}��X����v-�g>oqxWL
.3J�aޯ�����#4���بy��|�% մ��2�e��ַ�q)��OdI�^�e�,a�����j3�|��KDPֳ�<Fdi���x
6�Z�y�AsT2`���w�$�g�	�H\�f=�13�yũ15��������s��!`&b��72D��e�z�����T1 �j����RSDRx��4����o�v�U�Vp�y���������j�c482��`5��]	5F�j1�:�i���C��e�3oI��Z���>��p�L�S@41tţ��6)Nn
���x����������b:��Ta&�xU%Oc^8�%�;K�����������b�'G��Ć�� �$S�d�1�D��\j �J%��E ��Ѐ1� ,�o �A'c<�&g"�1��������c,��!���7.HRKk��}�^DM�/��A7D2�s0�gJ��p_=~ۧ�D̝���L]�d�ڦ�wa�N�[�X��l^H�Q�Q��/!C�dŤd�����N<��r���z����E��P�A������O���Z�1
���S��땗Ą�����W���*oa�8|��{]�h�b�vL��,���=��ꙣ܆�L�jT�[�h*��c��p����㮥V��j�e�\��%�f0�@<[�W��#0��|����=�Md�᳦�8S�R��ihԙ�@s$Cg*� �F���s����%�W����~�H�F+�;�v7]��	y���=P�1��o��a�Dh��g�>��FS�bs4`���!�Q�2�I�^�H�C�SQC�* ˮҔ�p�Q�S���/�ȼ�v��Au8��S�q�Ǐ���)i��bҺ#��}8k�J�b��0���� �Rj�?H�p�z�¼�
HPs.�$p(0!� %����/*|��eMΐ��ԟe�8���As��{�s�C��t���vi�`�C���$I@r(	y���f�������ݵL�l�"]����2]�p\������&�*��}�Z�-1��OK��k�܇1��`s��A�ap�:�usBRB�������O�Þ+ �i�8��sa��\��j����@�S�s��9I2���yQ�b�tY�Emè�G�uQ�M��V|��	 ���ok�C9��1��H�/��,A߾�>�mo.�����k Q@�lN�r��Ǥ��9���2?�!yƭG)Dc� ���x@Գ��nF㢙Y)�C7W@���c� k��M�Ls�%�-K���uڼG�?��9ש\܁��aMrӯ�͟��e�s��,�h5�xJ�`!��\[X�0\>�Kj��B-:va�K����b��(IC�^1Y:6K�Y!ِ��a&["�wD��ܴR�Kbu��
��0ќ���ϪQy�w�Ҭ~�Rka��?�Q�m�<�U��Rgؙ�}��b��@�`֎���o�,��C##��w�����m�����s��\3��q���V�<�O�4^y����n�sƎ}W�?Pv@p�(l����|�q����U�/^���l�������4.R	\aP�$�t�Iˈ:t�Q͌6�	z<�!)���7 f�I.B���A��z�ɮ�I9ơK���E
�����t�p��8��]Km��i�*w��x���dO�>V�i%g��cD}��UR�r�E�+2�N��~⼏���8�[=�H�Z&52I�;ģ�C����	�!3�ʵc=�]3sq"Z��_�3�`�2B�P"�s�W��7�N:��[j����.��|��]�`
}Zx���5����{�Sj�����9�.�����y�J	g�e*��v�ɅH���PB�a���Q��T�5�<��=~Q)	�ȝg�̎��Q�I{b���Z��g8'	}��:���vg	������f�*).�n]�����pճ^;#-q�MnC�\:��Jr�/��4na%�^�֍΃�$'/qZs�x�>���q@�Q�[���k?�l	�R�5g��1�֑ڬC$_�|���/�"��g��}y.3d���,�0>�J�qo�IqK�;jh`0:�-��X�#��ǳ���$�W��ýK��㢯V���%�K28��tT��{�-|��N|H�,5�)3'����{����^RlE�Ρ4��ǵ%��{W;ΙӈWZF����GޱDV�̈3�ɱ��> �C�0?�����vU�#���;k��J2n�8�kI�sԞ'6��x��ҰU�7J��OQ �ʔ(�ba���nz��̐u��bs�P\L�Z���<��^��vg	����z����R�@4��]X�2��p�\�3W�OՈ:A�� O����%���o�{��_�V�T+IE�!��Pf�g�j�f���Q��uN���Ӷ%�`� �fC���9���De�0�U���mt9���;���D�+\Ï�_%�� A,i5R�5t�����Ž|�?���o�q-W۷k���uۗ$���`�\�L��p*��"f/��S�
� f4�^H�L��W�j�b�i5;]H��"�,���u�+l���ˋE����iL��<���J�3i8ޕ���3n	�G��o���3?���G���0^�{{�)MոF�N�s{��F���y'�%��>F��g�;�!��5���̓G3I��*�X���;Kз�a��N�9ŕ��E��K�}f#��g�ׇ�	�'�;\����;�ȥ;�
c���M���!-��Г�� eX��Y��fL��֦��j��]����ꮺ�C�5����N�D��"�g�lfVHߥ@�_���禋J�bHv͠�+:#�c��K��cjG�d�4B����a����C�:_묳�L��������!s��nt�����U�p`��� ���'Z��;��xqG8��6!�9�I��a���0�CER2���=t]g�	��Z��ia]k���F_qPLO�(	�l$j�bHEߝ5Z�	��=��@s�V�QK��3�+6~����U!�Őq���G�>�Fԕ�d�܅#��5
c��f�E1��,���P�1�f�K��t�܇T�>����V)�fJ¿�vg	z�6QC��y���H�ȋ�)/���!g.}���l��~N�A�<�x���^�n;��H�������GkE.��3�uHN���'5��Yi�Q�1H���Rڜ��`G)�����lIEUg���d�S��IF$�r ��gk1:���.A\v��q�9!ю�Y���(/�`����)����q�uA���\S�����8���C�$ԧPqÞ+aZtҞ��V2z�C�*{<ڜ8�˼�k���c��2��Ì�pI�SjGL:;��^4�@�p9�� ��h�7i�c����Q�
�C�*\��_�<WBΘ��t��&G�S�@KM���+.r!�B��I	�E�!TGV�T�w��щ�s�z��Z*��,Y�_����R���F���i�&J0) �	�>8��H�7΃%e��J�J2&3[�u�~��B�㌄��@x* ��h=�"З�"�T1����E5S�]�B;�T4%v�yw��az����1����ts��E��m���PM/��?�'�CQ/>�I<�sA��;�PR���T���S�A�Z�v7��@�R �-g��j�z�H��	�L�J�?G��t ��@H��s�#'�P���I*@@���(KK����R�D*���	-p�4'N|�{��q��uէ�kGc�-yW|w-1�_�G7���4u�������0
D����֢�W����g�܋r����5y�ɺVA)� �,9ͅ�1h�u�!)[��ΐ��^`�+�*�s���U��J!�А|Q��a���o�Wƾ�qᤳ�a�A�r��u��Ƥ0L^;�H�C5vx��G9I��ߛ��.�[�%��{��a�oC��w��^c�cibMbC��j�����X�qZ�q?X
�18���MBP�wR����ZzL�L[��jm!�ׄ~�?�pW�R:�:?�������BLJ�@ �՚�sVLp�K����(�<6@m�x�R�R�S����u'��26&��φ�+{nI���wt���+nf���9����q��T:V�0jE=IS����C����o��Y�~}�r��Nȩ��v�]J~�	�ja+ F���x�v�3���SȈ$�D�щ��O��	�U�p�6KD��g��%J�Nf���0+[��ӁLKUBVc��o�C�tn����E0/J��Q�\�?�)xCE���=Y�R��X��Һ�{����:=�Y�h20��ǚ�B�U3uo��TeoԐE�h���(%"�XI�K�����'U�:0Q��!R���:� �e�LK����D&{IV��WpvZ)�|e'��AR�v�h�y��E�X�s���q���$^�;�:���MP<OcQ�7=o]VB&4��XG$P*"��x�|S�  �q�;�e�cx05~О%�5vFp�x͝a�
{�bX�1h|4�sjC���3��x\�C���oq͞�x�lt�!����0-�Z��?��A����axO ��8�_��!��@+Fr����Du���k�}c���̨�/yR#~� S=$=o�CQl(��N'\��_ǡA��&��G�� �V��Rb$�L%��Z�fЏs�H� M�z؏��Zi�� ��jvF��:�iv���;UC��9sHC@$y�;?�Y�k�@��p�!!j^jPs)����A6�{'УIZF1f҉���d���ɓ7p�����AƬ��7��L�~m��h��j��.]'�41�&_�\�HƂ�)z!8#��Ȯz�`�
�A��nwS��.����l�
L$���7������C����L�œ;O�r'�2�'5�Ԟ����Eh��w�=��_�6"�O��G��NOδ�N`�sed&���^��X�Mg{Js����$�"���م9�e�/2*K�u�i�X6�srr*�]˙����d�2�N�ׯ�G�ݒz�w��?8�<]?쇠���w��ǆ�y�۳��ڬ�u8uz'��{��O��jP�|	��+n-j���1b���/)�;PuN8�,�������@߲�ʖ�S���B?)0)��������3X���\���~��_�����j���Laa	�����8����@��A����s��@5B��.E��t"��|.F��ʍM7����@�u�8U�O8��({��F2	d��Β����K�^]q?` ���g���8�3�U�'��E�G*V����Qf:�TW��: x5}�ON�x2�����'d�\m���g
2ȿI�8J�;�{,- 2JN��������C�̔��Kc8l�G0������QSeyI.��Y��5"�؟���C�aXF�ʥ.=����1��"�7$�ڇ ��t�!��M�E2cIN�b�ZO{��;]ф?*Q�� ��l���'4Cf�h���rI(]�LU�=`{N��P�N�N�j��v�zy�N��^������o �b�	�XP�WB�{�>'�+:?+][Yb4�����Z]�����T&�2��L$�2ƝfcMD�F�j�"y��364w^�ڭ�LQ�|Wv���	�k@z���"If��}pb8��0j���In|Ȗ���*i��r,�HD�X���e����nkv�	p�G�ϒ�߃������ ESQ�c2'7029f
tBM�;L��{�6�s��.�����������j,mC�F�C/1ɮ
�@�5�ON��a�zӬ�7v���̱�����T����'�M�^�FIU��on�A�$Q���q2�3�o��KϞ�߫ �}DB�eLU@!kJ�
g��kd�J\`��~t�ϼ~c(�8��u't�;٪������ES�1�����9�GD{���c�����A��Չ(T\}PCJ��-C�kb�-���9ׄ_�u"F�K �O,�+����%p��xE�D�Y��IǺ�\�eG�l��F�9����U�f��.�Ü��ݚ�.8}���n�í��C���$��J��7y�8���6�Ҋ�g*H͞���	��a���>b��>/ڧ�� �Oݤߛ���� a�x �߅y��q�:/a�V�I��k7IB�$�%Rg�b�';_�{K�lB����� ���Pص��1�Uڞ��4^�x?�$d�ug����o���7�6�ECE�Y�|�i�rG�~a�mpB�>	"��4D�L�8B$ŭ`k���oq�&��p�J0W\�4������R��E�I0={>��8����D�_�����&襛�w���Iʄ��������ϟ?O��[v��Lv����M!�K�_���L���D̯�П�GH�$sl�˗׌ �o��6f_��D�����'dE}�	Qub�����pڋ��^0�3)�����*�>�7l�O �ja�ʖd�*���T�#v�!�C��݉^J��lȤ$z��bj`��:#!�C{���GT��*�HȽ�'\"b����3'8"�������~��"&A$g|ܿ�vۃνK���&���H���|�����/��I�E���ߵ;0S@�}zr�g��:i��I%��\M�� *��X��{zvOL\&T������Վ���"�1��p�#�/HQI�dVZ	�N�/��y]__1�bj�1�;��Es���~zi�h]�]�\'b��Wr�����O�w���;Iu21ݴn����6�P�J@+bΧ�O�����9�����{���MsCN�MD��L����æ �b�E�"�w���q���a����x� UX���g���j�x��������E)���,���_û�v 1���X��J �Q3���f�:�g�A@�{՞�L/�2<�i�M���	���g��z����i���)�T�x["�V�<}�Ϗq;�<0��H���o}c��Y���?�3���z_uӋ~����5ؿi�~�:q2�����������������q��$�A�����	A�O��r���0h hV�O�\L��f�HF���(!�O�*�����{	�C�/^��"8W��X �=x��OϺ�?�#�t�u	3���:�8S�>@νS[u5Q��@��cNm�|UK��~��E��ǁb�Nc8� ���r�/{�_��o�$LZO�A��̄��{QS�s�MX3&A2���#���g���D�	~>��3=�%]L�$�>x�c��p���a���~���l���~]\�gd{�i�܄@���N��`��x�=���ι�I���)D���ذ�a����o���0�%R=ڝ���P����M\�`���0Y��e<:��w*=��gәc�9�l���n���C��5�a���zk������՜�)#Ɔ�Eg����*��=�L�f	�SY50��)��ޥ5ذ�P����@�w2�K�1�_}�����?�C�g����P�^�w䬿�ٴ>�u$�0��Y�������g����k��A��q|���H����,��tt���Z>�,�)DGD�:
�8�����c*��?���{�/+f����i �="�pH��+mw��O-�i=!�ӛݰF��U� �蒤CH��Ղ�z�����8�0��4m9��ц�5��O�j�h�����8O�v)��|�Lw�8�텐��N��mz�Ȅ����U-}��-L�d����5� ���M�U�ቊ8F�5��AƟ�t�����E�k�A�9�������Y��%�T}��D�Ú؋&�ԃ&=�M����%Kz�4��~��R#�L^�gP�n���A�IF$ǝ1�{tH�`��Mש]��D��T$%IEkD}C�H��N�<`� j`Xp.����N����{�>jt�HSI�pf،����JM�����r��e4/a�N�	A��R_�m!~/�{V8�5!�� �I����[F\�al�>���	#��iM�J��s������h<���b���9���
���n�g>s��*�^�����}�� =qF�~d�����s�y�}"-{�㢒���e=]��pI=�b/�;�������	3���F�O��wt~������:�|��������͎��OjtH�'���=]'������}z��h��t�������x�1lw����?������Y���� 	���y�>��s#���Q<���E���n"H����g� ��Ñx}��%U�^�x���I�p��땲���>��'�~Hg��!tlQ��։���Sӭ� ���~MM����%h&�Ï�J�6�,�� �6@�!]����YA�+3�!���A-���q�	5��uI>J�^�:�/���;_�1Ƭf�X*��H٧���S%�0!�3�;@ءy�/��A�$�L'5�����D�&�-�����c"5!����}~~2�KV����[�6DLLO���6O����}�w�^��cd�J�K���=���C��o1�����㆙��˷�÷ߖ8`g��!�/�3񥹿��K�ty�0/�X����Q�qD���S1ov0�k���%����"��4 1�	g��כ#��~��H}U��$MQk�g�D,����5�[�GH�	��)yZ��~@�f>���5��7-=G��I�C�&6ƩL��s
���6v<F�~zv�T�EuvN=��X�����`�������nw��?z�(?y�����f�ݮ�~"�Q�+���NI�gz�:U���7)���D��S�����
����D�σ& �a�D�";6�AL�����
���ֆ���;��9�����<��8��R���MK��=,7�}GBc28y�d�9�YR��ҧ��M�	�;�{|Αy�#+���� -!�P�������?�L��q&1a�]�(�/Z�3YJPH*���J�[8�B� y^^��`M$M�F42'(�;�&FS������Wt/�a�y*܊����@���~9�wc�=e��Jג�eǄ8kr��A#=����f���c�e?Ek`!�%��S�_�8y!��\�*Z���8%Z2'B��;�4E��a�v��<W4�\Z����&kiN����>0����K�e��Z4h83���K�Ș��K�,_�U����d=�S��n{/��JD!E���O���MD���^�O��`0�3�8�v�/��q��^�z��>	��:����}���O?��rz���۝#��M��z�ڬ�&��d�ҐM����$�42R,k/R�A?C�% �"яp��F�0g��Bp�t�X=�D�Of��1�W5\_z�A	�;���d�U`�M/;�c�z��a��� 貦�w�8{=V��I��ڍ�0��O�]�s
ϋH`�e��t0{O�N��(i�D�ل�����~�'NQ����A �A2��@��V����Cz8t�@�jI'�lp�����B\qt]��R͋�&!�G�j��}���"��$^���lǭ���o��������7�5YBY�rG�J�=1�S�2�/xrF������@��ѽ�=2ّ3�2QEaM���E�h_��x��Y�f�ռ�0U4Nv^T_ffth<�*!?7�<�Q���m�Ln`ƜP����;�˴[��G�4����8�*Q.����e=NJ�*Y��H����[F�2���5.��72/����B��q!Z'�O)�fjXdp&%z��������X�2�8vBSG�a� � 9s�����ٓ'���n��x��;GЩ={�[�vێ�sZ�@k��m	ɒz)h�j�$l/����iL�80Ũp�0���4Bf������� 0�s�x��zp%�<ף�ӗ*'�|1B*ģ�ؑ��pɷ3(LS�߈~-��s�Z)��t?�2�I�fX��8��������ep��6�C񱡛�
����"ɉ���1���u���aX	Ed|`���)@�ݬ����� IR'���W`�`g�qJ��n�2FI��
,��2e��*��$va��v���Ȓ��T���8e�2�>h@O��x�Fa��鉙K��ɡ���
�k���|eH�«�UzW��W��Vle[@,�o���dQ�.�Kuu��/Ȩ�Aj��C/;��^����E8A�3�Oip�8+hW<Y�������\j�ܶ������,t�\�PΙ���"k�*���G�:Ŷ$�������D�j\�'0Q���`�^�W�/^|q��?��#��q���J?��8� ����8��ljv�^�elC��ĉVA��pG2�+�ߕ ����v��vO\$M�p���#s�y�&ԵQ���%�[1�I����1����I�G�;�䊏)�����R8�ɐ�vH��cЂk�$����ԋc��| qSŨ8c''�����_y���k���R�3���RP�kuȡ�3�-����m�lgQ g�I7�\����koo���z���
HH���aps�!�8�ic��7��V�%�"�hgLcgj�r��N��eW����u[2�4XU�|S3�j_J����>Gi����_1��B�f��>Y�>�.6���;�FQ�K�Q���i�ڢipឨ@��	����e����t�����޽�O0s�zJ�4-�g�z�άj�A8R�v
��FH�D�JXT�P���<��9ѷ�gA��szG��<�i�)"J����*K����$%4j��-.=���������8$�<��]�h�[�4 W�����P��4�R�%;%��WN'��)2$����97?����ҷ��_�jQB��E��a����1T���:���m���dy��%�_ű�:7�w�R�c֒np3z�T�9%�o g$%c<Z�.�U���sF5| ���U�'H��]���<�-�E�3+�֞��*3P�o	0Ue�aC@� y��`l��[|/��G��:�{S����L+��ۖ���9���O�"#=G����`��3��~kc:��zy��?���?��}G9p3�w��*�%LBH<y~԰�w�9������9!�x�Ε�!��s �(Í��kǛ$<�3C��r�K1-��ai >�:�������	�sF�$���$�,���v�r���D4jR�+`R��h�K?Us���L*�Qj"Z�Ə�kb_kq S��m�Ĝ��i����*�XB�*�\�50��@�N�-G~�5���z�xg�vc l��(�XIv��	�P�NƸ�� ��D��*���f���)CX`�ծ�����t[`l��'cʹ?���b���H�Cމ�>;�԰�[hc*a_���z�ϗ�D�ï�7���>`S� ȶ7��o����\��ZhD��w��v-�4��O�<�?��G	�=�3g�KI=V�JཝA�8`� ����L@��	z����)z�jB%ꆨb[ͨ�3a%v9Ed��驱�;\)RX�Sq.�p��
K�����Z��wF2mU��4�)� �v��"qFҥ(�ʼ�s��n��k���|�)�Lb�,�����e�{�G��<�x���tW��j����ޛ�O�EQn�{yEŵws�va,-�[�\��X�s������GdT�ۿ����>�\��8ǶEA��2�?��*���l)`������:��9&jr {Nn������r+���U*�V#��i�m}Qc����]�Сv׊�'ϯ^�����OBG��%"և�v�����c6�@��&�^�^*4��9�V���V�Z#�A�ߑ��yr|�<�(�!�3W x1��}!YB.�Z�#Lm�Q2줮�I��3�a�\�{[�7�,3"ND磌��|�2᝛o���*���Yr̉�n��a+�mX�R�����l����Rk�\:�8�M$�X�3$F�;��b�OJ�s�$��YIs�f���������ʷ�H)���uK<��ƭ�b<u�&������z��]�����n��ɪ1�W8��v������N����|o3��i���ه��\�-�sI�WFSA����'q��]ӷ�W�_ާ���۝#�￟���U�{M��u��D)E:T���j7)�M9��P��4?H�8����E�^sɑ���g�n�"��.a����א�h�+�W��Q�0z�PO�� �z�b�Ke�ؔ���g�%ے�Y_V1`>]#<!݆�È�o{v�b�Y�s�Ty����`"#�y�>ԌQJ���Z+��t��:�^D��x�s���s-1������K���k˄y�X.y��{]�q�ؘ�Tt�mG��e�����*`�o��?%Y�Ч3L��1���GN>_���/'7�u��@���!t���/�h|k<C~�b_.ġ�Nß��(�OI���뒮���W//���ϟ�~y�d"旔�5��XDO��pl#��7Ơ�}����	��<C�~��o�\���D�&W�Tj��*M9e��b��#�!��@3Ϩ��[��#D�Z;�$��8[�5d+���3���gQ�`����y���U��� k�å��zI��p�,iM�$�eiđ����]w��v)'z���v^�m�ǘ��E���`1:�ő�h�0;��l/�俊.�B��v�W1���澄,~J�~�ۿ�}YО��9��$)-���ϸ�m�%���
�g6��*��?-k�t4xs�w�+�{�WJ:d�#v}����˳\~��>|8��j�Z��'�������0]�p.�88��kN	,֝{�G��M��D�����xH�ߔ��� [�.��u�di�"�M��r8�#&������̣�"zC?����H������J
ud��W��'z�g]ñDǙ�jO���1r-K�l�5�q�/��F����G.=�U���w5�9N�d��?	z+)ȼ�}sr�P��R������7�_ge����}k�(��Y
�s���q�D������/%<'�Q�&���3�����*I8j�|��Z]����Q����d,�p=�#sZ���ˠdv^�y[zEm��f{�W/�����p[f��=�� ]��0�7�����<(�i�Z���8y���mR��t�_��9������������������_��?���hwu�������*��If��g���qg��c]rBH{P�{mcH���b���)%�����{��́H��'�gBJ�Z],��L]գ\�P�DU��F�UWe�F�|WKΉ_�� �f%��6 �u)�Y��lq���%���g����Xji+���(gJXGO��.!�V�KMk��;~�='���w8���e�@��[�f�#�j��	u���{,Gb�s�Ʈsǹ�74�7�ai���@�����w�7� �8S`�H�����S!�\8�ȻY��8��.��/�5g����$�,�T�BI�Z^��#>0]t��ɶ��Z&��8�3�r��?;a�yfJ�L��﫩}��5w�5��
�ؓTs��s��h�E:�p8�as����ڝ#�����iU����������o~����ܜ����5k)��N+@q�oM���8��>x�b���ȺE��us�A鏎҆*
��R�jf8#��˟��]be!DU�`"ca��T��A�bD��T�۪�P�J����b���[��E��F���E;�p�:r�>�K��0��|�)$���Θ���]yG�����-Ơ6R�2rw))NQO]k�$�A��yƤ�9�諭]����2m��^�4L���|�SLE��'φ���b�B�>��'^���ҿ/\�Jڏ�P:���0f����	��kǱp���.Iح��J^�4c��ļ}�G�f��s��!��3���|�U�M0�K�g'2����)�Tϣ�{�8�\���?��ֿ�l/��ӛlw���������������o�����ݛ�nM9����*m��N�$�S.l��4�}���z�w�G�Z�tGI;��X,���z�5&��5m��V�O�)�~ ��XF0[櫬߹�@��D.��b��Z�[��L�K��ABSK��Ħ͵��a,��pD�낅*���Qg��ҽ`e�H3�����U�G�k��T������vK���-kpWN�VB���������˜&�O���B��RLv�*Ȫz��<��#�0'Y΂�^���VIu!&>j|����w�������1I�LA	L��F�K�%�<�_�J�X`��'�*ә�~ɩ�$�GԌ���eT>�m2�p�����<��p�jf$�g7N�WD�v)�bȏ��9�b�2����ˑ7(l�iR�#\�s�]CM�-2���~y��v�����[���_��������Oo��Y�N�>�`�pX�׌鞿�JS7*��"�����Rq����DA���C��	 ��(�]W�s�~X��(<��kz��]��$ל1Ml9~����O��J}/�L|�H���w�[�j��~�����J�����}��0F�����S���F�g�kD�i�ֆ0�*��+"8.��n26.Yn�p��y�]����\���b/Y�����|��6��p��۹�UH՝V����T}7�gh�jV�L��}*��&-����iACT�n}$�L�갧�呾F3o�9����2��{`�+
+5�3'ǵ
je ��J�Y�bｅx
�*66��.��v9���&�f>�[Lt�.Vs\jcBEd~Ov��I�szB�/�`DQW��5�D�!=r2��k����Tfy�k��+����M��}2'�7��4A�>{���L�v��b����k"�S��V~rz�upY�����NW��\�u�+',mEUpEO:+�#�_�a�k\���;�k�"5IV�R� [��Gu~@[rH�.�XsꉏA *���^:V��%'�9.� 3&�B�]՚����锦l�i@���h?Z������X�͐g@Պ��W�֫�0���avK�����_l����J�@���R0*�٘7F�ya���J5^yE�7�ߔ<�|���6�����
�nafC���w��x�4�6�����c��TlI�p��Yfp�\�:������y7@�]j�=S�������>C�e��ZVƦbI`"�9U�>�oU�$_<v]�V���T�FyT&<�=}��l?	�����m�ڝ&�7e�ˮ���t��Դ%�?;��hi)h���?|�v:?������鋧O�ˉ�{����o�94g4�Gr�;0�Uh]����8����چ^�v�gGl5@���(��H��6~a:u��:���F���&u
W7hf�8�P�<����Bk�/�U�{j�T��G�uS��צ����ٸ�`�[ܞ����ZG;�!�X��X����mZ">�<�z����N .Տ��"��Fc>�;T�A`
�Uc�Fc(^a�j����L�
��Һ��iW������srÏEX�r���DQ�ldlB��#���N)R�v��8�c�1ӊ4��aKf�B�$�3n6col+��&�)���<sܯҎa�M�x�W۪���4DDJ&�P�r�{ ?4��:�,6J��n�}�@a8%h�x`��A�*i������i�ڤ�ɉ�&�I�J�>{�|�����}�:O_R����4�P)�a����ӴޜL����#��~?0���Q�:.�x��mnO�D�&萞X��^�3)y���bNc8��/�<���|T?F �t����i(
���F�
��I�SMlZ�X/���{���j�G�v���:�Q�1�xm<�;�M7$��,�d�W�{�}��ͳ�Ɖ���+�~�gsq����e��M� ���$Zd Zλn���v>�f�T�cr^qFE��>E~[3x����A��Rf����jmd6�I�Ϻ�&ԭY#5�+�_DM�FUm���^Huᳬ�*�؊QJ34$hЌ�(3B���=��P�6�H����6�Ț�,+Q�����-dT[�Վ��^�'��^�QsG]{ڿ�a�܉�с���E�K&J�X�0"5�s�7`;J��ǿ�4���%�,���|']�sW�g)��)<�b,��Yø��dT���x#��obܫ��]o����_⨙�������}���D����n�N��svJ�Wҷ��m��]�����ψ�竫��D�V�:L���o��i�>!<*J�YƗ �]_o�Nv�:����~�x���^mos�g?Q��+�@w8��>�g]���`��÷��"B�B�W�
�fT�i3�m@�yN�LG�i��(��"V �ˇ��(U�̉.uQ��~U:�����~��_Q�.SA���Z�����&�I�-��e8*)S��Ʒ͌�9�L�0oK�܈����s!7�`��d@�z[�\���s{3�Q'T�\��R"�iyM�FqKZU��!��PiHjq��z��Q����l&T���� m�� 76�l��L��jf[u5ϚKkB	��e,`�w��˶>��q��!B=�c��wN����0�8�C� �������������������Q/Q��w�|u^%/���#2��0��_�~�ęYW�bLW튮y�ȅ# mRE�gg'���x��lk����{��%Z`��sqq����5lzǾZ7�Ń��}��搄Nf`�����y��?�g�������^}�{�[���W��4A?==�N�����ݛ��Ŵț�wGN
�F�� ��,�$�����T����9����6�ը~�o���m^�|�L"��z�P���l�o������:Ta�(�fl�D��6�s��ʎ�9��n�ϳϸG�bxA�ѻ�]%E&��wi?����޿�b�E�ȁ4��l��aC؋1Y�����Ϧxn�qaO-7z0���5����s@����;�&_�d�f���E)cToB-�u�Y%�ܭ�v���>QsepPf��G�0�5��>Gg�ҫq������	�}NFl4y�
v��@�0����}�>���!��`]Ӓ��i��ov��OŖT������^��^�p�����N�r�qG���y��C���P|fM���䄓��V�K>A"���{1�	$8<�@�A܋r��I�^6<fk	�B��X��iH)h�<�D�������]M�'��k�&�}:�w/�����E��f�ĝ�}���J�G�j<��?�������G���;M��{�ן��l��?��ôF']^�w���\��B��y9�lr8H�-� ,Q�X^��R�I3�l*�b)ϨR6u�"d�=��2�%C�;���"�щ���7<_ 'R08�C��hÅ�m���J���:��?��C�E�e�F<WGc�RX�91�C�ܳ7�5H�5�f%�%�ڤU�|^�����?j; Dde8��Y`��>�'�;u��Z����"{_ аqP���s�S��RNpc|�X���b`ԋ[������ �'���s�0�s��f��������U�Vz��C0�ˉI���7Y���H�L�Gx�GI8�zU#�&g/@�"�QHg���$uF&��Z�u�~z�V��X���*Sx0��D�7}���*#�#�5���\v7nշV�%��A��9,ԣ�� =k
`єP%�2�<�8w\I4�?�R�$(�H�J7>���5��@y=v���Y�{O�i��I��w�����r��Ͽ�v�	�o��w�?����O��/�ǳ�ӧo]�����������nw����`�A�;��3�8eP�\��S�T��B�#@\+�&
�X���'��}`6�t t�J���W�"� �͘��H�~�ǃw8qý�\��c��������MAo��=�k�V����~M<�����~jFb�6�9���"u�U�dK����$�z��n����fX��n�\;6cU�
�u{�Ζղ�W�_`0��U--�w�w���{��a>��YϚ�/�!�O ������G�3�k��9��X�)ӊ+u��F:c�Rb3����j#�W:�Ν����s�9����4����|����M���u:�4Z�+�.�� ��5�#"f�O�yLR�ur3�������>==���g�����?�6t�7|1�����w��e����G_��~�k�E`���7/��� #�n�m��}o�3[�}�t[_q��0ňN�1��>:�H��l�%��d3�u��L�G�vɣ�r���9�������}��rڔY���oS	�J?K�X�\��=v_|'���w��u�
�(�1Jз��Dp�1  B-��������o�����0>�,��cm�c��\���m����i�s�\k�ߩ�WNx`�����0u[k���Am�#����{�C(]5����9e����G7oAY�}ݽv�H�3���o{ѵ��m	��a]c%Z,�:�����R)U	T�ı� k���z]L�����t�8=�����_}�_�������o��>}	�N���}�o�cܿ��G�wuu��gND�&�����slyv�8:��� _����=4��mpK�\#}����%-a֊s�Q�8����GD�~#����Z"~��h�'����J������1�]�q��w�k�,5C��x��Șk��D�Z�C@� ��~�o��:>��j��) 򴄌��=g{���Ao?��Œ����ь�+XM:�FsP��j����
��Fci\�A��X��m�ÉkKYg��Z/Vrl\XZ���s��^��&T�4��2@�J$}9�� Ayב*;�>�fo���g�Ξ������o?���������^�x�g9o?M_R��!�>�Vl��0�O��U8��dE�b�S��Y���ZO�$�x$���]�e���Eh�E�z�B����& �W��?���(��g���ҫ�-�k�Z�D��<C���Xj�|�+�1)�F"�qp�9�u�H�z��q�6�8�q��J[Dw�����.v)k5tk!WxJ\DG��+�B��;�!0��w=���f��Z���K�-l��R�ĥϚh�/RusiN!�ֶ��O��;b� #�z<���`�՗zWR�g�F^"��K����DD��	����Zʅ#U�'�0�:�Cr��ȒR�	� �q	�H�e^.������c����0W�9"�[�x�M�Z3�И�5z��n�N����j?ᗏNOO�������?���������C����A��������X�|g�,NZ#�ݣf�;E���:��gx��ku��T@�<�0[2��ոiy_�����q�p���c�%�Hj����H׵�suf$��	���9wF�8R�kK�D��~Us���w.5����!�R�k?\������\�����Q;qD�W�}�K�E4t�t����(�uz/W"����xq�qvYT�c��9P�̠'ZJ�)�}��J�t�5B��&�V̉^�u�w����w�{ 휪�<����z�=� ��]�^�7������#�N���{�J�0���ٗ��}U0�.W6����(5�d>H���}��J�I�k�Zֵ��GϬ@��Ɂ"
&!�>#U-�Ϭ#��]
)�u���Ԇ5������g��Nhyq@�����5rҺ3C�����I:'I�s~����O^�|��?��I����A��_�ve<8I�U��N �H�PaODI������ؔ>��ޓ���9A����G��Ƅ�t\�Z���G{�.j�=���}��m����;�*u�?r�w�~����`�s|�?/},�3�fv�C=�FD�}`}�loq���ϑ�om�(�!ر��XՀ���:+�%B�%+��L Ig�Ic��q�s���
t[������m�Y���w�\�E���&�+!FD7}��1EkG�ªqQ�^��*k�Z�^a��I��X��0�nl��(3�	� ����9�W��{�CQ��P������Σ���;��Uʑ3��pM�i�!�!	L�C��x�C;b�^�fO ��?�g�x��1Q1SF�I�kjs�z3�V6���5)UⰵC��F��"wdCO7}?|iRyl?3�'?I��ʨIu�8k:�<V�R��eW]՟�Q�U��#!tb��{��n���s��mu�*Ϳ��-U�]V���,���Χ^��V�c�ı�θ���x~����������3���{�k+pN�r�a���(�}m�z�,[�ې���G*	G����%͘|���<�)��:�/�ȃ�X�T���M	H�����?a���ބ����BK�0��Y�U�}���r���ٶ���/�xC@�6n��5i��U�[F�3x���j��ʐ\{�{GD��<ϿQGåql�����Cկ���������F/U̽�D_�}'�X�d�$�J��h�c�g��_\\�����fɽ�r� �`9+[�+$G�q��)h�q�}�ח�k ��Q�lnپH�ܬ�+:O�S��V{��=ǫP��;�Mdf�՜p��V��q�꾪�[lGF ��<�ɈP����[�%�1���!�������M�D�ֿ��<�8�̥������&�7'�7Ղ�'~�8+�
�?'�PQ*N��=�ʤS��Z��x��:̜]r����}X�gΘ
SS���6��UD���u·��a�x�_��e|�9�*wC;NIa��w�+|.�WZg��rJs��^�v� �	%0���q��+���J���5j���u"rr�-C�J�<���Q[j?3�Z���h����;�|w���þ>��~� ��$ZKn�P���p���>JC8pnrv[��9<�����\n��2b�&�Wa��^�j	��3z0�ߛ��������h�1)��XfF" ���W��*E5oi��ܸ��o�|l��������Et�|^���2@n@��y���\��}y��͹�낹"�sࣷ��c�M�49�;A�oɭ�*kE6��EQ����M�̴���I:�Y��&�6�9�O�}�t��=T�ݒ�)� ��P 
�%k��["|�������/kA1�ʁ�����|�����{�-��(�OH�V��ued�Dڧ0�#��[G	�{�)�T�Xm�T_Q:r`U@i�m�5�4��h���]�F�l:�5�:� >MI�oz��ba<�%.o��V�>�|�I��Vm���7U�e� ���t�ax_����L�D�	�O��?ۘp�$3��cBȵ@��[
�yi�@�)�����[֌m�;���3qF2����Y�\��J�E���[��,�0w������}y�^=ߙ��N���X%j
�deXFM�[Y������3D�� \���`Nqhl���,�i�c�<o ��<E�&P!&�?g�����=e�9p�L H�6���c;ä��}��+Ϣ�I�HX��(�i楜�eKTIy���z���-�[���/�K��ZZ���;���G��m�mI�P(k/j��zfr_������ċ١3*�-����S�)31J����9�̢K[�J�x{/�ע5�>� _��]M��
��~'<��x<�5k��nשo�� i��� 4�5�c�֣8ެMޓi0�)����B�U�&.ydUL������R?�d�d9#�C�]�F�}Y�Q �
PY�z�n��4�t8_JH��Ē���$B�1�vމ�BW=mz'��D�G�ToNh�g�����JzF�y)�,��x��YMcR�.�%B�r����2ߡ� ��y�p���<��@u]�y]�� }Q�����8� ��/�3{e�؄	S����9�4�IM�Ի9=���އ<򲭌��ji^�A�OJ-�?/+{�V}�t�%�8�,�&
`���m�w�3
�!���<["A�jOP̯�N�g|�`2m5}�E���Y��̀��\�Z�]�D����_z�SϨU߬����eS>}Z*}��Z]��[��]�	H��f?�D���V�>��;���"�(����󨓙�Y�I����\c�K��e������S�mJJl�d����[K�Y���:�NMp'2�� �6�P��R'8F��,��UL���5���24��ނ��~�v�0~�wSbi�<��5�7= R0�(�2J�8��g�[�&���>�]*���,`��U�Lt���Hi�;ڐ�3�Q򟪃d��Y�qW�?�Ӳ��X<H�Q���=ײ�� ��@�.�>g��M͘�q���bl&�<D�&����\��QiJ�+����G(�%���\\,}�%�IN���$: w"p<�6���r�.�^�aЪ��ٜ�����j;�"� @� �Ǜ��� ~���ԧ���p�Y6 w��1l�'����6L�{$�R]�6$�LiJ����e$]���>&3A{I�e�F-p����.��'�I��.[>
L�Ĥ���Z�L��������+��7n������8b;�)Ԓ Li@�%=jD���#­�{���,���/ט�~����VFQ��vZ�T��P{���2��"e`�����W�R���T���V���}_��&&�s���O}�=�t�~5��-a�I�6DL�v��Z��s81�������ﹱ�rL;��|�)G����L�c�l�
#�fxIgzw�k�2�d)י@N�B�I��_��E�Ar^I�81'Kkb��i.7au������@�A��J1��M���N/�*4���8��PYz��b L��~3�>�E�B�B��r���kW����,�m�[�J��"Fe�o�(W��!��4F�\��'Sq�\�)�8��V@��!��g��o�<"m�EqW	ǵ�-K�hy�kU����m��HZ���t��{�V��^]�l%���}떎\d�1��ؒ @s�$+|��U��`�l}q��m=�����j�@3QbF�<��A����R��N>�<{sH�(�G���\R-X�gի�g�2�OK8�:�jqȒ�DC�X(7BئS�q� �;V	�!�0�a%E�tH����ȰH�af��<���Q hҼ��	M-�]Z��JFe�Ο�g�M�&e&�-��PQ�͐�$e�O5����!��'p��>zU�GT�s�Y I-p��$����-�_[¤2< �3�']��2�L�KO	�|��*i��q�o����l�>�m�6@K�I����o����uc�m[[%V�s�L��m�4��l���f����dIޖ/1(�۴���R�	҆2��t%��cU�ny66EƀY�Ja�$�˙J}��?I�'��Z�a:� р�
�F�I'�D�oE7�p[tC.����ρ���/3G���̅�\�h�	E�
�y2�r�RZ��<��e��� fKCT�x�B:���v���]���X:��Z�(�N[��d�3m���wE�Mw�v�%IL1N�7А�
��]����OF�Mc�&nV����I��"E�����6�������������|�ph#`@Y��u������!v�Dg�jc��?s�[F#��&fx'��t�.���g&ǑO^��*ȡ�������P�f0F�t�,�:�a����/ی�0��<���6sLbf���Bh�>����IHIL*�����_���g���'�&�.�'4n+6�XR���y�IA���������i��X�f 
�)Mm��X��}F��50Y��A�����\5��`�K"e��PH����ٛ�l�8���
���mڒ܋z,EPh"����E�gMޗyD��M���|�8�i�J)_�C=�mZ�7Z��$���ƾ��kz������F&3�OXcR�Ϧ�r�9�	& o�n/����ɖ���@�э����'e�Z�� �\ܓ����D ��x�o𩮫v8N��gg�/
;;;��k`[�$���k�ɦ�-�{��H�;���֞��O���X͂I�bxԄ1u[t�\���d�}k�����t�s�t�li����uJ;YE�&z)$�.&�z*u h�V_��}��Q:m�@c���S�!����]zG��T)�Y�DB57���‖�:��ԅ>]eK�J���E`.�e�� ɻ��Ό�L�\��Y_
���Piz�*���']��y6naT�9��Y��w")�b;Ǿ0��S�¿�v�����Bp�����*<U�����(���	��*��*�5|�?���[6D!�
Sd��as�����?8��;���5�v*��>�'LQ���BB�b�3��#�!�s�W(fNƨ�E�8���2�eZ�lD�Ï��>�i�ү�ө�jՅ�N�	��z2il�X�aLV���ne�#�J��b�/����[Wa�K�����_�Z]��EU���Ҍ�ļ����Z%�Yj �4J���6��S�������ļ�=_~��Mڊ�2��g�)<���2��G��<1i��8�\Ú���[���q��j��uM���/���dA���\j�d-F磨�qI���dlJ<6qc��ꏬ�R^P�Ȫʂ_���)1�����X����ې�3[~�[�g��{.o81����m��i}��w����Ӻ��NF�g<I�����\�*}~��Y��ݫ��=�4��8&&��:�d$fpJg#�`�l0�٘��� )�iOΑ�ǂ	2��}B�����1@ʌ���V9b������2D��!hd���p�_�L��+d�k 4��E�.�M�5��O��S���q'tRZGZr���	t�9�R˔��l�t:����g�}��+��&X���Od4w�:tN;����i+�Ƅ�<i=�۔�˽ ��ʹ��2RE���jOcS�ss1߸k�ҚMQ��ƪUk�V��>��z6��2��W�Q q8��D�!A<�S�#r��M*���~�2���+��,�U	Az׍k��`�З�`��t6;B-\7(�[��tk�1QwA���������Rbe����d'T��T
�<I�zh�M��r
��	�韊־���ܩ1�d��:沋�H�t!R��
����,q��%��8�a*%��扝吤�9L�_%����D�����m��=��&֗��Sۺ����}�h�QK�ή���b��;~�5/�Ʉ���"dU���(��w$s���}-���0]V4����5��Z.����Y��|���d+�� ��T㙭��/�O�����2n{�ήzP��pۭI���kӵrH�ɏ�TMU=���'�������������|>��G��w�H����`~��X�Р�oR�CCk�k�}�4�:�� B)�'�F�xj���BB�P%C[<���`hJS>T�#�6)�6m�,��_�4�`�4�`�o�[�t`����jNt��0�FcԤ��L�k��A�0���]���i��#2�J'�?��ġ^Y�j�9f��1g�g��rW��\���.�Vґ� E�����:2>� ��Q`'K��PW���X�@j�l�&M`(-e���/�����Yg��L��z�I =�ɴ!6�6zGg���GB�`^Z~=�i������r�w�k�]����e�i�K�����������u6�������J;}��nj�*3)V�������G���0fm��h�	5NjmQO]��w?�O�xF�bF��-�6��d1���ig�Ӌ�pP�\�P-�Ĵ<q�LH��&'�Y?���s2�����i���M:��a�HN3�g\�~���2���GmL�K Dm��t#c	��U�5z���"���L�,i(���f %ƺ
��jifm?'gE�P�
(
\�,#u
�Y2���MWrZ�/�T� ۶�Kam��Bx�~,�m:B?���/D���T�Tًz"Y�a�c	+<��R�~E�i�������uU���q}���'T<�Ы�-)�xEԾ&�S�3@_&��
_��T�=��*��,]��ό#��#������|���.�����5���N�d�Zc�D��UϠ�,�b��VMG�l�ۄ�N�Ken�Y	��V=�-2��r�У����O6������ ��VѸHPP����p�Xhj����	�/;랶D�x8kO�t8u�M�ȸԓ}���̂�$t�\&&g�2rix��J`����L��07�򺻏!{h�Ր5m�,�iX�������yK8@����wG�_���S	-i���"�U����A��eYN��Ѥ�i�T������gIͪo�qG4�(^aMUM�g��V�1K5�����˷��AM`:�"s�����C'��`-�8	�5�3��a55��̙�����4�O2��B	�3�hjf�)f��LV� il�q�8��������)E:s	��!]��6G	�[�F#T�Rn�^<H�3�o�J���CHt}F�B�Ĥc'bv�"?�#�L�6�.+�)��ʨ~�4H�lҴ���y�bXnE��_S!V��a�k��Ӏ�zZ��K;�a���<s��RZsv�h����T%���
��V���V�1Kh��V	��s�#έ=<�'O��-՘�G+?���>z��K�}!_�]H�:�t%��������>�}�0T��y���W�;��,�k��ip�U�D�О���xĊT��	_a@���TE0��3�0���`^�O�U~N ��7��IK9��Yc=8uۄ����p'�kV�3 L$X����t�T[V�O�Ц~���	�K�AH#�LRi�Q�M��4B���N��Z�y�'h�t��?���~xtt��U�q?���[˫��� m­Kc��7if�U��m�A���Jxh�/a�������)"!��W��g�F	�jms�9T�6����Z�w�B�y��������Z��l��ha,��	��@�T>��u�n-s�[	�{4}��F�8�)T�6� }Q�pႹvm���f�ݢ���-�O�md��`f:i����䛂7m-�I��0i�$��N̓!�&J_���*�T���x��D"0��l�f���eeQKTi 0�b�)�&�U�@z��mkI��w���Ĕ'����mB#HHX�7!��[��+���84�Љ^�t0'	j&e�z}�-��a��-Q)��F`�q�=�,������c���0n���O�Wy�H��`�V�7�
!���l��(�vKږ�����mZ�J��(��������B�cR5�b A��p�s#^΋�R�22���r��^bˬ���lYk#U`JV��o�ƥ����t���z�\��r]U��I����D����zN�7�f��!�ɉ��������-�D�L���d��ĸ����) �mn����z"�kC�����˔t�NH�Ӆ��:9G 딣[�B�V�Ϫ&��(��AH�Ѐ��2��K8J褢�f�����|�J ��@ĬX5�[���,;Sh�zr[h1�ƌʐLȝqޭ"%��7�x�&,;i�L!�yd�)�`͠�#u3����/z,+�k��V��l>S:�OY��ABZ��Q�#�+����S�p�[^�d5��{P.������J�%��q@��GV�e��8��I-�5rq��%��2b��F���SA�� ߆�ݏF���t�;�%�|��
F�/���X@�ߦ��%L�1Q���;��.jA%�u9�6�-;?A*�dq�~�>��!�8]/�F�
k����硉�_�ȸexҔ*��
ɞ���-U��W)��x�J��d���Y� Dk��L�4Ѥ�7�/1) (;��=S,������} *�vB�VQI
KG��U��8��$�h�h���J�1�)Fr�+�%�*�;��T6�]WF��P������q�T� n��f��H�S�zj�HT��S��:���UK#Y����9ݐX81���IKm��E�[�	��?{�"�u�k�����>U�����K_D#�������ea3{ʧ��*��y�,U�xRZ�u�k"�`�З�����j֩�q��E���.�#3�34Ͱ�eB���ڐ�p�Dk�!)K�K5	���m�� X�Ц�T��E�f&�����|I��R$4��t�Ie��n&s�J�Zs�
��U�
s��0c���A��4��𚿗q����E�P�M?q��j�g�@Ɩ�ETt��T�X����V���i�<��PB�pݷ��n����/$���o��I�#�hǭl�!O��
��}�_#8U�ɒ�F�1j\�P����R{C:.;�4�L��j�(��2c�.wo�̃�ֱ�*[oMhA �9P�-x6����j��b[g��$��,2bS��1%<��f鮪d^#����r_~u}�uR�-���O �I�:�&�����\B,^��z�d*��d����1�Dk����DIܐ)/H̥�)	6���zL��u�hv�R̽��-hm�kB�֊&3���Q�i-M���r�D���+	D��7R��d����&JSJ�3����D�ۺV�:������7��� u��1ܶ,$�q�m���ދ���q(�Z�;�C;
ml3"��UlkZPAfOF6$ ��DP�[��60b�B��^)Zr ��(��+1�&Ʃ��s�V"��sl��Uq���S+	I6k!���Q*�>[�xX�J��&�3�AQk��Vrnl9D��8R�E����Г����۫q�O�1�b@B���Ȃ��畝ܖ���w��m�Nsc̳}��o�a�]۝5�mt�z�Ȏ����a������".�a� Q�6Z|�k<�Ma�v�YW$ٚ�Є�Xu2m�	N(t�c5|c�$T�X��	1������Oq*A���t��H(�b����WWV ��Z�y��`����b��'j"�) 7�^�&s2S��G>E���.�E-YJPC� �E0a=�^��������rb�8(Ju�)϶O�+�pX��Y�uо�G@�Һ>aR;�y�� ���2�Z�6��Ѵ�*Iڊ̯����-S�64�Vu�}m!�yn�Y�q>��۴-W,(h��� �s��v�iH�w�	#�9�%ּH�T��{�� O$M5�56���0�"��1�J<|%�� d�n���<oi�VU��[7���a�$�/	Ü����ڦ\�ԁ�Zi�D��A�%�j) .g��=��Xn���g���/7o޴����b�/��A��eM�>���͵+r�	bQ��z"�y��^�$ݴ���z鵩�O+	P��x6ı��3
Ayb(k��"\H[���2U:�R�*Fl���B�_�l��hB��+LƊ�� ����Z?_�V�_�~b��ԫ�uU3�47}NJ�kF*�!>%l���w!k����/���c�b�0��MN��Ǧ�yu0� h�Uܴ�6m$d�"��00C�F*�6[����@=����@'<��B~��O;o�iڪv�/�Z�;c��%��E���Jf�k��VޒA?U2�aq�n �{�{��R���ϋ�D��dyK#�"�GƓ�zh��"��ؖ�0P�����C�| ��AXS�1�&TX0����8V�7����#j�6����@v���ӭ����e���l�w���sF�e�U
��d�z����}��u�q4��at�	�@��VM�ژf���C�q�.8����#�f���ڢ��S�������aF5 c�]B<��Z��t�
kDZ
�4�H#; �L4�=��G)���meIb�ۺ
�_� �k��t�H�<�>���m�V��FM���/=MVLtAz�&�����ϙ�~$���h0���`G0w�����_"�>�`��b;h+Y�|l_��ح"X�߾��|���?m�ǭ^^u�#B1��g!5To�]P�:��,8�4��i�<:X�^�-�����9l�>�d�d,y��M����;���X,�W��Х=��qPf⠝��0�� }���i,���ޮ���S� ",�c�*������H��~��/�*GUc���eL딭�p�줸�a:�uz�I��\�%�5�"Y�/�7pC|�v��4���a}}�C6����B0�`8z��h
Df��W� ��\0mp���7�pa��U��.Lc���G�T�#���vQ#c-D�i��k��5YOo����.��`����<=�j�Q��@oUuE,#��`�����Pch&0�r�Y�dH��<�������&B�f"�{3�w>��@ #�L�4!�p�I�/AŌ��1�A�dM�0.�|��[|k訝W�Z�c)�u|�t�g�~ކ1�@97�/�p�P�M���d	�4����	�
� � H��6�o:��V���x�[�d
!(��-?� &�0�q��ƻ��q�M���"�DB�.�.E-4��C���PF4��|��4�H�*zhy��Cp��A������pp����.^�0���䠮c������W1��vr0����g��,�FC�5�Е��c�rP1�X� :���:�m^X?f��p俵������8�8q�����㍡�r2��0yMK��-4��H�J?9���DkQf9��dn24b�����X��F@o�64�X�"g��wM&�*����`i�yT�zR}��S���/qE�1^�l��C�~���O$4����D�m�vd�P��Ȑ�dv)�[f6�z�)D��-)K�?L�B+���f�:�N�9�<�t	�#���Mp k�)*�_�Q������77FU�v��-�N��j���6�9la �Fj�*n�����{��.=	^�g�������^L�����  ��IDAT�@�&�KM�D�:�f�q��c-i��F��� �������Z���ֱｷ��Cn�,Պ�����M%�J���S���������/8�(@���H��Ig���"�=];�r3\�����8f5�#+�ʽ�mL�DS:j/�����E�u4�3g����k�E�41�F��s��kf�]�[�t��X�j�6�_L��|��S`(�H�ð�æ�5X��mb~��&���w%�$���m��:#}�В����Y��U����K?�6��o6�����T"�����.�P��%6�C1c�׻��Ѫ6�@���
0�k�T.�7A�K�(L��6��Pd^���˗�p޶ۍ��{hb��'�(��>�[�C�"�eG`�h�t�`l\�B��bqѮ����yC5�������3 Qy��b����qx�s�d1����HH��U�#�&�^s�̏��.<�E�����z��i�^��$f�,X=�cXu��.�x˹�ʧ��i�hJ�5�A,9S�ZK�R�\�h�ZشJ��OK���)k4'XX�4'��n�v�8�{0��k���V�f��Ą�B�Q�*gA t`�H�J ��>Zܦ���t.���Y�$12�K�j���s�Ϳu�����6���a�RǁIZn#I/��U_E:�AZwM����}�O��62.�	���-�,�<b��lF�������4��?�< �;m'M\��%!+�az4YF�F +�U�/��,�g��@x#�#L���P�N�rZ�Py� ��ha��}3�2�;�i�B��?�),�0��'��>�0ksHy�2p_�~s�UKP�|T�ֶ�f:�>>���� �_��_ؿ��FS��M��=�sfC�f��Y��<$�De���;���Ld�l��:t�2t2�H"Ŭ����eF��2|��!-�H��R��$K�3�M.`"(j�8��p�R�Ĉ��6:�R��>�i����ʵ�cR�������*A1�$�R�R�^O�$�Y�3��C�Ng�S��~����z Z���CH�т[��P��8
ʘ1<n�s�E��#d�Ͻ����
�x|[�2TZ٥ouL�������2:���o�TG����Tiq~�[l҄��̲�)7K^��_V9�������0��ip|���5�ܬ@d�<3�4LB�C`*�<�}Q(�aj�_(q����ܴ���� }I��'�\���&.�=Z]�6���H��ffU_Q����0E�},j�&2k2o��^��=�c�k��
#!��d�W��"�,@�{Ao��T:O�-|h�ks�U�0�V�Wj"�*pI��K<?c��G.���dX�罰jO~�{5Y�I)p}�����1ic�d��d�H�)�ڗl��h�9
��EZ���ˣ�/���}�NF�i��'��2q���x4?lt�B"����� �Lz_���V��,��1d���4�5��M��g�ѠL^��*C����@^��M�'3�	]\���2yPr�� ���UZ7^K��;�|P��i��&��{�s{�x���Xb�z�ı�'CO��a�#m�(Z�|:] ;�{�g��Jh[ܺfےg��R�d�S�3
Ե� �G��	V�l2��!{@�XͰ�MG!��e�:Ϻ�#^9y�� �L��*AЩ�*A���B���� �l��m��:�Eɖ���8:�d��,�	���X�=�#~`�/���
��J��̂t��@?g8���T6y<]=����mF]t+���mI\黤\e���
%�_�{C�Eiʡ,,E��Ǘ",�����gȬ���$�ڴ�h������&)��FVjӊ�����d��v'�؊4�ˮ�4�����T4�� ��o�������`~U{$�d���"G`�K�'$cЄy%2���7��w+x?����M����n��z�'nTh�
�c8�����y�-��u�r?��l��^%9��8��s��1{aV��8��%�7g��:�{ڪ�:ctI�K4�N�B<��ܗw_�.��P�6����L���b&+u�]�{w��Djnt��r��y&�m���yq�o��_�Xl�������� G�r���v5ȴ;�Bu����i�ohY�NGE�Ba��9�����3�3:V��Cvdu4D�yrc"�AQ��a[cp��;�[����O��}��t:�y�泓�V	�H@=j��>�G̦���4c3� �Ict1�$i&XE���E_H/�x��:�� ��(�f����>����Y��l���>z�,^��>������n���?_�Yk�Τ��s���цÓz������t,	��2!ʖ_�k�lKsT���i�*5p���X���x��'�q�[n�i6y���g��z�+�G���4ou�<�`�G/|�ÎZ>���+}��^8<<j/\���W�M�;(�x�ZD<Ћ����g�k2Ƽz����RkX��y���L�䆭ek|��]!��L4w����=� ��qF��s!�j`�z�M�3Y��} �,Oˢ���Қ+��ɱ�ϯ_����1�m2���+��D�Գ�ʸ���L�S�T��D�R����iX�ܓ'�c�gV}�2nK+�R�� �mﰥ�Ub��qbD�31.�ڹ?��k!EB�2ơ�]�;̩S����z"=���u������N%P���k�R)]��M+c2�$�����a��d���Y��r�C��Κ͒�LT=yX�|ȟm����������7�$ ,&\�5�=�� +�U�0O���o�5�M�})�N�옚��
�g`�:�s�%A��wч*jZT�V�۴�Fd��ck+�63Ň��*�bV�U���&B�Q������'u������=�$zo0K%�r��I;���j��P�:Wc(� �[�e�r;��@��tVɣ<��e|�aI�P`W����6Q���8�u���L'N�~�s�о�Pr�=^::�l�4dVVq�vitE�^�ڕ����,�l�uK�x�/I�V�����X"˨-�T/�qn�����?�8^eg#苳^�
�ݶy�K�dt�;r"�:���������"ʓ��;G~����'��N,���(��&k�!G�������B���T�]@�
q��[�G�q��?�}�O�-�<��*��C=/h������N\�XHJ�Bz����r�f�5�c��j�%�ͱF��o�q�u,E7�|�In��.%����{��eqW
��S�y�ӒM�L/Kj�ht�e�P��-L���#�	��c�i�o�ggy<琙޺�Iƛ�i[�E.++ZOZ�n~�ƍɟ���������pb{f����h����w!n��v�ɉQɖ��rG�O��1��U�f�i�<�U�U��1����<����'׬Vͧ$�4�cі��i������</M[��?�}��l�XV���;kg�:��jPK$ܖ�Cڸ�<v�O�]�rme��1�kV�	������m���ĳlDf�9��x2������?�f�5t:]��c^P��Az�VɝC����K�|�i��hro��n�~8���	t����3�<e������ٴ�n��`�J�F�/zs�LUϼ�s�O>�Q�%��1��(���R���E���t[��蹘��o���S��d��(�Z�/��)�/eyP��L�3�c���Bv����J	��B`�0I�Ј�8Zy���X������� ɃIh])X�_�&]��*GG5 1X$
M<�3��#j�s�/[��7����dx�l�-<�Y;�M�E>0�x�j',���-ϱ���DERg��:�J��S
'��Lq} ��AoG3Q�4���qU�n�rI'$L5��l�tFe�t���<�PnE��Y�yܔ�*D[�,7J)�Y�\��R:>,��}�?�I e����{�"��B�<-Sf��?y��N��`���e�&��]�Ӫ���}Zi�cP��M�y#׶��<Q�V�PO�e 9,�+Xش_
����h]��lH�$�t~r��Qq,�8�Z�����p�*j�|'\�}���50��������l�X?��e�{�qI}���K�d����b�Yo~x��~� ]�;��|Ե�z��Į�2��2�_y{fd�Aky�1P�VfV�n8�M&�~fF�6�c\C��E�x�Ϡ�\}t��9py��.�3�Wk��o��C?d�m������%��U]N<d���-�{\�<Ĕu
�<�+��Y���?^X�ȶ�y�:��i>*��:�4/ФE�w�N:�tS��'�U&;YzN��}�zփ��Q��ځ������?_> ��Y��65�w���Mn�ݏ\�K�׶^C���l��e>��և&�c*����]EJ�ُ��@��N�c����ǩ�v�'�Jԣ݂rm��2��xGh�O�3� �K_VU��h�Ok�<D�8:���9��̤�y>�"�M��wp�<���b���L�;�ΘP���^v��@n������?G�ru|ҪH���%e���a^@���d�9ԥ���b߱�yW��m����H�%}Z�,���dD-��h�|�h��,�y�SC`U���A{4K��\�Ξ���xעB�b)i/=�R�i���Y�>8�Ɂ(��x�i����F��
!h|?Wx���eУc
��[��'�v�u�> oL�]q[,�E��#Y�k��	�K���f,'�.�'N�7-]�'g�����f�[�xX��N�7�r���X�:��m�0�ns�/a�u�8>9wߧ<��P��#7ɱ��W%��$a�Qϣ���0`����x=3L�ϕ�g����:Y9�����	�A���dcUu�.ȥAs+|�5����3J�t{je�������\�g��}��賋���MP�G�i=���*ل~���F�ќYEPR���� �z�b�U��l�A������OD�Hq;��t�� �B�����#z5��7&
=��"����Q�G�����5iB�+n[o6�_*G3~j��<���1}��
ۦ�����9�[U1/�A:�S��9���(M���Q����4:.�#�D�����ƣ!��HaZ��M�nh�'��
��d<%�Kn�J���q��	n|�>�?�����}��<9��rc���`�e���?�_���M=�E��x~�yfn��^����d� �F8q�CGC��KS+9Ih̋�(g�Q&�'�0�1�3�jX�x}�O�C3ô�n�ġ�L���`E�6��<�!N��A�oEu�{���Fz䴲 ���D�V�
]ݍH�*�=Θ,ۉ㙰I�S�hS��11��8ܟ�ɬ�8#������!mJ�A�����^A�UU{@gA�t!j<�WA=Y.�Ƈ�ml�Z���` ���(b��y�8�`(w�C䡄ݾ�t��C]U*�I<�u>���GԞ$$�<x���"���/�d
Ԩ,�S+hƣ���Fe����+f��-ӑ�P-��`+�&m[N��=��'��jB�%6p�3�x��~p�1�g���:S~�;��h[7�����z�΁��.����$�ȫ�#D��@�o�0=��nR@�ߕē������w�<�#_)�8@��,w\�i�m9h���A0?6�Ʀx��d�u��8����*J��o�8��sz���0�؁Y[Kٕ|�T6�*cF�e�UA��'iBW9X%�B��E"h���	i�9��L�gp�b.L��"���\��`8<��Z2�ɿY���w G�Y�;�@F+3{5 4`����1��Լ}]e��@3�p��K<r���o(R�W^;o�3��O��>2��A^sL�Ա��R*��[�uK������>Ʃ,D���>�Q)@�x�Ȼc�d�u��};sV+T��b�񷥴�w���/�^����0�l�_%�Ɵ�@�/�����<<d��e�Gh��K����ŧn���f�3[.#���*|�0*;��O�r�v���0���M�тֽ윒B��'�Xx���_�-�&V3<�p� ݱ/7
Z���u߹���|е���xF���!�O�̌k�
�>����w��/�<XOC���*2Boe��z��̌+¶5���B�c�Ya�TkzD���E�II��g�@^u�G �<�I���W�Giz*j>*�-7L�q%QѺ~=ϵ��X*�dG�D���Q��Ө��p%c ���|��2R<13���Wh�;������?��V�yQ�����W�7I8$:�� e]J��<�g?>�����$����$�㒋Ү*5YӭH&��H ��Y,/z�S:���W�$L�ry�v]摚@*�$kUx=4**-�Xʼvǋ'i%�R:&�k�h}�X��hY���i&��":�yw}�<E~$)%�ֵ��ߋL���v��$��҄9�[]�l����C��7u���O�/?�@�=�eRh��\��;p���g-�8D�ey�ҒR��<��wh?{�tQ9	�&���|(���x7�.b6k��jN^�·�M�� -C~��fM��"rzL�@:���,L2��>f����V�1'���6��DzHGc�D�<�G󪭢�UFL��?�
�Q��FWϤMA���@�+u�$�O�/)0���l�YnR�P�?�Ò`j�| ��4h|�,���I����ʤB�H4�O����'�EGy?��iqQh4\ye6Vmѩ�z&"��}�I���a��D���j��p��S���Y+�\�VX��W�,nb�ӕ�T��D�a-���2l�z:��:����"��� ��A���`3-J���I���T�8�Sϛ��&��QfO�k�:�r,9����������*��Y��i
X��E".y�-�M�s�{�דMe���O�x�ѕa���bֈ�_
�$ƪ�%�@�KL���v��������gM0���^s��|ބ�^t`�S�σ~ۄ�w3i11����y��=h�6�OC�!���-5`�q���UH� eKM�Z��vS��*
l��՘�ϙ���J":D�}�RP5	8#H�|�S�O���YF�ȳ���H~2�Ff����m&Xd�(^�$`t�Ys�Ҡ����*Wu�����ۅ�S�d;�t�H:_� g�eQXꥸ������/���q�q������t���upH�/�!רi����`x�0�F&��Q�U����`L4��pY�ln�	�0q
lc\�*X�k���l�~�V��Ȭ�5���,�@��z�U_h��H�%!ҟ䚙��7=��X$�#H([-��k�5�0<�3� z��0�	�v�0��`�~0Z㯚t�d4r�����ြ�	��zz���8���=�}�y����qL���w��խ00B�8>s�)�P��`��\7?��,h�?�<+�٨��h-Oֆ���� ��$`��}�~љ�W�fx��'�啄�k�F�V���.�K�ڃvDܭ*�*y��+�:����߱J���Z�FM�A[Y#0[:W��� �K�	}�ژ�����s�G�3<��T��A� ���փ�B8����B�/mRY�-��	:��̥\On+��K�Í�Q�����1'��0ҕ���`�
C�4gKy'(`����k�r�@�#/��}����l��"�g<��l)�� �L�d�e��;�v�;�L�`�j&x\�s;��l:u��*��K��B��"���ư6^c�?�c��-���QcW3դQ{�U��dٳx��v����LD�N�<�eΘ�8����ʼ�/6�M�GTb��2-F�ql:T[�ln8Oa&
Dc
v�J'*$�����;
9�'���e���c��i!"���Y������d��\mK�)��U�����j�d�0hD ��\<XFI�.e[���f��tf��*������w򣉛�f�q�?a�
+�TYOo�2�L�.�uX\?�iۑ6?H�S�6��\ʵd�HSB$չ+$4[���g̔lC�C���L�:=ÂD��p�!�陁%@�Z��w�Y������4<�߃��
�G0�a<l=�M'�g��m�m�x0��?p�������&�������9��;���fњ�5v��7�;Y��c>m��A �ێ)P��ǐ+�@�=,bAL&>�F�)+�T�~Z�����Qb%�k^z�M����QpˁVƱ�X���R��3���3��d�|rYH|o��ml'0b� �#����m��|�B�mS�'��˼�K|����d�b`���,�x6���Uɴ�q���E�	�Y���_Zc�iJ�,*����Cm�:i;��ۍЌ�.0���,$�	����jǃ~�,�ȬOv��ٝb��n�]���*r��몥�tN")�E�O���)O��{G6�ph�!A�Ƴ���(�KLس���M��[�s�hZG`G�G�p������}_��;
������o�=��7Q���r��� 6��d6�8�G�P;?�s667������	�=�̼��8g�vemV���\�f�Q����pQ^� ���,�;�uv~cyn�ijٸ�4Z�v��*Y*<��DE�+��to��s!o'��<.�i9��
�3M
���ė�$�.wK�P��Z�x��I$���xt�L�{��{�u��U�+�;�@�0�����"���W��9�h�}��U�)}ӝ��8u]�q���	��5>X%'GI���J$<�X!����֦�F��zW0�'�\C�.���Wi�ꞕ�Y]E�e��p$���\���ȡ�t�%ФG��@u:G �{h�pnݾ�}����g����;a<9!`�?N��C����|��*0��t{����g���iߧO��S�N���o���Y���(���i p����=���u�	ڗg�xw���w@���F�r6�;�[�#li)���N3{A��A�p���M6����E�����c#4�� 0y7�Ǘ���9�	�||Z��+�ı���d6mة�����A<@�Ev�3t4�W|����܏�*g V�c����hi�������Z��]�ߘv������j,c��Q�|�3a�#��]�3���2�N�l�G�,>�L�S\���*1�cdoNyz�z� �[�m�c��"�G�v�(Y�:�'�Zf*f 9��f�NR�H�I�OaԼ��P���H�;��oN�H��9h1��H�U�U��K�2gH��<��ڗ��}����	&�6*#m&����t:�?�]㎇�w���7>���{^}�U��s�����#
���f���14���=<�wn��Gׯ��ݻp�
]__w��	���h�G��̙���̧o"���E�����:6̔U�2�%���0pl~��a�~�f�����^'�IB�W�=4h���TC��7i{~�U�Z���g��2t��еc=�Aut-Z<(�0�=��N�1���&k��ws�n[��E�������g0=���X�Ӻ2��	�m���p<��	d��:̜ 6C�k������&#�z�]_�\���q��с���{4��Cd�������0q�?u�3ǭ����GN��5ڻ�iĖt�_`�V����<]�<�uv��cm:��ή��q|{!�867a����Xc�^����9Y��Ie�D�9�A����������<����xN�'��9���"cF8����	'�!*l&^m�_�x
Wؚ����M����$�Ͽ5����
�1�ĭD���<�����!��6���Rvn$�3�M�Ue'޳�ԥ��,RѴo�Ϻl�?�:BROL��D�Ioz�����ެ�c�B�2F�-���(�%�u�s�ZC�x4+��Mg��ޞ�j�c�k��7oz����G;g��p��1pmt�l��[C^a�ap0��mU����O��o���\��}ww��]x������{���������~���5y����!FYD y��ڋ���z�Y��O�O`���pz 09 ������!�0���C]�!�y�[3�o�]��^�[�&��͕�	mX"r�k'<��SX�-|d�;p�������[�`>�x ��m��;��ۯ���a:`ؘ5���N���&�Ooa͵�h�ս�0��:�����އ��o90�xc<�3W^���_�:ϟ�f}������"�l�n�4�6\��q}����Ý�ށ{��|ۢ��U���8}�%������_���s�WT�+'H8��r�؛7���!��?����!�چᗿ
�/�Ë}�6^а~���Y��w������`3�����ڂ�o|�}�p��� �xú�� �㒵4���IU!	Q)��e^$&|�D���?-'Ĥ���N&���c�^>	�y�҄�ڸ;���M�1e��	'�c�tFr�Y�*ӪL���<�A����eP�ҹ���%*K6J��$ ��(]����PJ�Ju\�ͬ��a�*y�=�M�&z�X�p��N6��ɼ���k�mD������$�{w�8M���Μ>���pz�:�|���pᢿ@�⛦L0ǆ�B�U؊����h�Le��eO\Y�����;���=w�\x�:G�:�o�m�U?��쫷����r�������o��ށ����"�Q�-Ն-r�_kj(8-�K���:@�N����E�y�*�.]�`SW��K3�Z-.3`�N�M�5$<��Cػv��tgg��y�1�_�򿿹{����`��0�|�.\���/�p�4̜:i��:p�������w��/��	W/{����̵�^;^�������{�:P]y	���;o|F[;`�n,��F��6hii��0D'�w?���ރ�����Ln|�mW��
��m��N��g��{�|����ڗ����v���y��L�ٽ�8@\�N���$��.��X;����6^��v���kϟ��~� ~�-B3�hd�,T;g�����7�p�Z1��t�T�Mgd��(�u@�J�T�X:�<)�����$:��^����~	�����`0h�F|���pe?'�[�@3�R��Iqi�������)�����}�,��	������V�w G~����?���rԬ�3Z����*��O�ҥK��s���Ύ_���E�Yo;m�;�E��\{RN��D	���q�:����C�1�O?��{�����׽������@sN��^"��+Z�����S{:�ut ��z>�o�>��`�9r�>�C�X����N���x�kjg�)ρ��N}�4l^|f_�&\��oÙ�1N��}W�W�Q+�v�l� ���p��{p��~�s�����r����b��kP{���9�~��_���NS�}嫰��
��`�5��?[����@�~�.�47�����#�X�C����L�]{�5�jv����a��~�+Wa������W�c'HM�̍g�'0��:|������'��©�k��l����G���a?�]N�x��.|��[0��/`�+_qq�����A�Z\{����;��-�p����y��8��h� N}}*'�,���q`N�������ъ���n4�\�z����p ���?.�E�m��[����4�K��=a���*q;VA�=��LǂG\��_���u;���ٟB8��^�ڼs��O��{:>��]����v��{R1�%�_B�u���J����/A7�����6���ƍp�4gtV{��|�}�[[[��M�Ғ������=A㻎��5|����5��_x���ս�=�z���>�W��G����;��;æXmY
N�ý~��2�MC������࢓֧.�_��̇�s�+g~4�B��Ʀ����s��6�@�4ߏ�� ����:�9���mh��0�?��o��p�6��/?����?���=��q��:0�N�E*��q�k��k����{N���޼�>��4X'x}���Қ�d������~�3��?�L~�3غ��śLa�?�����L�(@�=��]�޺	������.|������{hF��
�@�Nᓟ�����͛?���w�����L�e�ƥͭk;�~v�������Ҩ��p����{�p��N��?8f}��_`�\��j� ����Zn�[�ŷ��M<� �(�4�,�;���.����|2�c����5n�ف����!3,��C_l4����tC�?���2J!��0,��y*�9eG��}���'�Q:l㱜�a	�����Ǝۙ��|[ۢΓ�����XAKB0�&`N� ���s�f�{�P�_z�%?ܨV3�#�7j�8��-��JSƛ�QX�����|(D�;�����$X��&�WLqȣ^k�&å��H�@�Q�o�-�c�tO���9l��{��Z5n��^��u�""�|>�'���a����i�N�����>tt_��ַ`<{mu�K7?���_`���wap4�^݃�z���	��x����4�:mc�=8�C�f�h�������.n�������q��]���6����۰yx�y����G��/�quA �އ���0���(\̦���p��)g�,,��Z��ڇp��_���.��7a˥[�~�;�M�	�Zscg䷸'(U�܁q�{��ܽw�pT��W0��
l��6C<���k��?tm=h���Bb�҅�z�>>�/Kq�� a��.�c�[�~Z���A4H�<V�1�Tz2s���.����@���)�TX^PN��,�Z�|����8!�8J�Ѵު�����!�D�w��F�\��ZZ+� OZz;�V��V��<IKG�,tҠIcGM�o<��_����N�D�S�x�c4�c:Ң	�e|�?c<J����?���k��X
�����L���lj`�J&F �c��o Zf��ǁ��������*� ����S� k���`���5ؿ���
�k��}�!\s�O������%�p�,
9N?��>|��������=�0���`:C���ں����8��i����o�2�	;-�������c�g`��0:u�{�[>��������k���&c��?�sW`���`ֶP��ݻ{�^���>�Z<����+W�K��=�x��pԳ�1nAt���)��;�vk�8�h�Ol�y7���>��W�u�����|��=����3���o��/����'���e^�4g.�i[�ۯ2��ߺ��K:a=]*�ltp�@�Q�u8G������Z�r���֎��n �2I��IZs>)˴z�#��i{�:6�o�+��a���9�#x���k��@X	��s�������z�v���z9��_"�?Ͱ�=I�&P�Z�~��w�����)n��#�^�v̓��-^�F&Ly���eDU�%�䴓��Ûo�酅�_{>��o�ǵz(������;p���J�@�=��F��!�g�㒡?���x�G�*liJL�#��c�E
�u��p�g߁���������o���M��nx�l8��������`w?��	!J#�
N���wށ�;`k���7p��u����B��1��w`h��G��^s`;�;;��o�����s��[w`��� {o��>�P��j�`�0�-����r�?�������hn~��_3v"9�s
��_�/�����s����u���ӟ�~��?�W_���߃�W���8�G0^G��Ӕ�o�'��`��v&���?ru����K��w����	fk'HMN���g?����p�7�p��-�������wa�7���S�\��e��Mܦh!ު�6WotGV���n��!����­~3g��~S�Zoq��&�)�|�a�#:��&U��a�|� �缜oV�v����XʎFN����i����E�l��"C���-v�Xe�E��|�-��V���%��i�+�D�2��#0��g��D/s\W�����Mfpr��JGan�l@�1�.��Q�o��9�N�	�O��Ϩ����N�؄W^y��q�%~_� �5����L���,OU�V��2�9҈��8u��_}`�4�N��yVN��vZt=�;��`����6֯%O���L=���]�n}���~p�i�����6\�����믿�%l}����p�p��t�9m�����v���3����wwΟu�~G��@s��������b���N0�r���	C��4�m5��̚+���S�������/�t�<L�c�}������7az�SX�� 6�S�������58��U8��߅����^�
3'4��; �v�_�@�G�)צ�_~	��ο���W.z��v;k��� ��E��c���@{h����5\p?u��M�X1�[��m�Y�+xQݯ��\���*�������Z�sV��*��g˘M��(�T���éʟ��,'
�]#��_���q�!����e��,,1��_-���Xc�c E[���O;�:��?7=��iM����pxx� ��_;'�nݺ�Amm��qE�__�`P��~8m���9��|�Pwq��m<d�s{y���(@���K]ڸ��6�)=N)���~������KH��pF7j���4�.�R�� �w��CW��;0�{��7�C5�}��jך���'�͜�~�6|�lM`챦���O��ы/Ë��?�ګH]N�6<n�M�<�/�q@}t��o����{NPp �{��!
���P��+����okc������N@:�B�����Y�9�	���o��Ӕ�N�5�Ӎ?��>���H���Nrx z�s��m�m�; /���U��>0k���pэ��{�p��\��k W���x����>:��3^��3����������P�p���0lW��3G�?��K���`a  ��: :DkN4�%'��W�/ˢ�k}QǉC�� ���[[�I�T���m���������g&�e�������M����:�7q4Kb�=�-�L�A��,��MwXG�"�=)z�7�	[��t���E;'hM���q}�F���˗�������������н����yp�r�%x���)C�}�<HӦ�kEO$P�#_1������_�����������&y������XܞTp=������Ӳ�dRS<ji����	G��*�W5So�:�x@��k���; 9
�=p�~�>9Hr�%�&���C[��s�`���q >�u��܂����w�=��o�����
�^��{���&  ��q���5�'���/~��x@NN��|v�_s�i��v`c�4�sڱ������i{o��@x6�\���-^p���
Zsm>Z����[�#�U#��?���5��g7��ބu�����3 P�8�^�������W���?w���9�z�~
�7�\�/��#��?�`R�9�w����c]�'2q�/�5'@�E>�|z�W[���񼵧&��/�>���f�@3��tQC>�D��
?s\zq�ϼH�-ƭ�i�\��"��c��q%��ha9r��l��#~���nQ�~Z�� �_��_ǔ���y�=X",w����G����֊sܒ<~]4N
���_ǰ�����_�\Nt p��`V�xp��܈�u�X���9���qn�iQ������W�m�l���yG�g��v�[�vv�x�5�;N��sA@8��]�\W?�\�DQ%vܚ����8��x�_UG�?L\skӆe���º���w�y�-�8Ae6r
^��:���	<x�W`���<����5:sν�:�~����5���]��>p����pZ����7`p�e����a������1v��ڮ�*���9k/���/��Mۃ}��f6���;�u���l\}�/	�.�M'8���@�?��­��߾����9Ý-�x�l^:��M���[\��~��ݏ���d��	4vv<�-'�{�+�~�"�7�����9��v}�$dyG��G�.������p>lo�s���������Kc��ۣCx����w׵��-�����!^���Ҹt���i���/.��-j^���h��˵֟3�	�^�ŋ�=i���,�D�h�8�/�܍?�=l\��f�)�����7������&����[���t���k�~g��粒L�x�үix�k�����_Z�mk(���b�w8�5i������٥CM��� �#@cZi�g���	��fAx�oh~�t`�fuL�Z��s�a:9���5hZ�{�]��:�� Ν?��?i������&O�R\�� ��{�&��νv/�jP_����G�`}�F� �����������*~k��w��	[��
��-8���@�{� ww�:<t�� �f}ܟ��H��/ìv��.��b^��q�z��k����s�C����O���w�p����c\�/]���K�윇ٽ}��z���k��sʷv���	(�쳧at���zνzμrF;��܁ᦣu��hF��L�݅��7`s����(h��uظ�GӾ0�:Tи��8�ǆ�7��p2E��/G�V>��������aY��
���[݆�x�p���G������{���k�3�gpyc��Y&~�=�i��5T����v�0V��}�d�?�T}R�dM��l�:dq���Fc�*�>1����={8��_7��pi�����n�Na!��ܝ{�[yӷI�xn��掠tr������N�r�)�|w|�!X�8�v�2O_�X�v��ܗ���L<����`�����IϽf���װ/^|.�m�G�;@�����5�����u��|.����j<��9<8�� ���Q���5_�}��ۖ�Ik�GL�n�ņ~��/��&��n�o �{������I�'�9`�p9���������p0�l`�����lL��m�$wu��M8��7`�����v=�gA��:O��2s����B�
��;l`��pueF�V57��/��][���`�Ln}�5[<`� H6�yDN���7��o܁��ߡ=�9�����A;��?���N]�9��]���v ��לV�*����0:{��9�f�����Q�n���~s�G��S�����@�}�M85ݯ��6����ytD���S����;rqƮ}�s/��y�|<��ҏ�7�7�(�9M}����o��pkU�̱0���w����@�+N-#'�~Lz�Z��V�x�isg7m6ׁ���d�h�c�5�}f��d� 羛����xÉtpݷl�N�#�H���Ė�� ��S�4h��w�=���@��
O��Afij3Z�&-�����3#X��|4{@���>aKj���.�c?��:�qڶv�n�?]os�5L:ʑI^�D�8̫��I��O7GG(�W"����g��3y ���������s�|�	3�m���]�q����a�oJk|��.{��.�8�;����6�ۍۭ��I�� �eWy�MҁN,���j`��)跍���x+:���lu.��v����Z'l��\i\_�����n}�>�&3��~��E�M����k��ѡw����އ�������{>[rd�a'��}޿�����`f9;3˙�v7H)��"�O�s���~�7���XR��ٝ?���F�=����][�:&OfV�{�z�m�������Js~ǟ�,��mX>��hb��`V�T���"�=��{�_'Ot�D��:��͓�]��ց
	5�����6��u����� q�㘶�"�q�T���S.J"��܂Q�Y|#��c�|�r�z�A?r��c�𿥈�K��{U��F������u��n���h8�:��y&�4�>S��uР��_���(��'^�2��1	�^��l�1�����,^���G`�UqȚfd����<��q�GNRt�}^H.#�/ai*�[��ʞ&�	@����c�̃��s�SiϞ�[wjR%h���
�:��@'�$�b����3W].�b�E�� %�$"��-�Rך�S�F�h<(�j��ې]�*ǎ@m���$�h��`��_�ϊ/��<�(#�t�ĖJ�:�ƪ��������z2
�=f,���@}�4�`iz����:J͔O���0���i��R�T������}������{���
��8,S�ݯ��6!�����\��	������R%�1Q�����M�hQ��+ � �~U�9��'�9��z�\�?�q�W�+���%&�J��*k`p�ڛ`�K�����1V�<�W��R�֭�r{��1�O��U��}��n�����x_��m)�����ǜ
�=���ufm�_����ќ=4���#'zvu��k��W��v�t�_`a~��?�>��8(�v����w��3Ng���B�HXJ�ԭ\��R�����ڟ$�i��Di�T����PbH���ީ/�78��'�K���N q���&vZ%WSU��y��3)�H��U�T���"��3WR���6O'm�6�=U6�ل��5����7��)����6�Ai�D��.���Ԑ��xw����0��|F@L!hTF�s�WX"%�C%%SD�6a��8)4�l�52iPNs��J`��ʠ�j�����)�~�5X��2l\�	�oނ��w���	cx�n�2�U�V�g���)���c��oܾp�0*2;�{�!�gT���ȇV������ �1Y7�43��A��%�������H������l��P�W��׀���'��P���8��&!��^*�k���'u{{�o�ؔ�tq�y"��Mr�Y��+�5Ñ�&w�Hh�A�,:W��T��Ov�vuh���y���)���iW!�?qw&;p>6ք��xj ��tO�f8D	�'j��*���0
�G-�v�]��g�?��羦�l7�X��h������Υ��t^���k���`rr����mhl����//�7��`k�G^��=OD�B��3%��s�D+gI���.U�����{9��+c��G��.|�b�IZna�[(���?�/���t<�Q-���ۛPy� j�]x���64��m�AI���y�	����6��G�R�n.�Ϲ���#^S�C�����!pe�9�&���s��<�}��ƭ$a��� ��1�6��xʞt�'�s������Laaj
�O��֣��=q�j�W�q���݅��C�1S����_���{P=���Ih,.@s�t|���W��#X�z&Μ��u�W| �����5|�z7��>|�~�(��1dlQ`/@6:�6""���x.^ s��#G�٪C�9�6��Z-0wn��Շ(�o�u~�١�;�W�Us�����W\�^�aOU��K��4���g
�_�#�oe�x�|�W�6��x<5�Nq��w�����]Z��P3�z��m��@��
:�j<*��G6��vd�3�_�)P�5��Iy���n�Hr&I�B�H�^�_�r�TF���� s�Ǔ�>�tN�꟧�_�/�j5�U���k�
o��8I|�Dmp1Ew���Q=��jX��M� ��&�P�~�GI��<sg������e�	`��t��+�_�6��;(e�Ы��$%T��_~�=�=}��K c(�O"47+(ewP�&������C��]H�M��Pb�:����M���lmC��[�X[�h���@�Y�M��B>��_o���z�)n��	���:�\��'8���� �Cx������*��|��R�$>�+�ylaf�����v�Q�Lj��Cx��GP�U�6ǡ9!��R�Ro�4!�T�&G��	2h�ސ�2���"q�;'ġ ��j�h# ��ϟ;��	�sy�Z2]����Ǥ��`�g�v���/ўp�/�+��M����7;��1\z�}?G��	����E)\����������U�$I�6��� :KKK������0�2�e�����������۱_7w(p���n�uH�O������/��dߤ�`ʘM�q%�'	bRU�yox
S#�8�aN����i�ԍ�oS�bR6�&��T�u�`ס�-����@���f���M�D���`��^��-�����*8^�w��l�Ft+�
I�e]CR�1�J��n�<PC�քll2��`C��=�z����q�.��-���z�Q"�?xp���%��MB}~�Gm����Y��;J���0��K����R��Z��TR�uDl��>�7o�X�j�g����NԦ�#�O
R������&���}�9v�ϟa�y�l�5;�6�@>�$S���q��F'	�ۃy�SƿN�m�3K�пp�"�Wqܧ�Y�i������~��d��E��CB2����BFo�1���Ϡ�ka����^������|����B^�^�����p��� O�� 熊�f쿐B�0rlus.�:I)qVh��gx�	n�E�/���t�(�M����~��pz+�-.z4���ŕ܃�16�=���|��9<x@F�,a��z�HU=!� M�K�ub ������7�)�J�V����v���x��|?}���������&"�� 5:��}~Gj����U�Ⱦ}�Kʊ����(��jU��Qi��q�َ^��f���+�����l�ڇ�(�sp��9V��z6G�f`,I��u���+���a�j^��4��zߥk�_�!�\(+ 	R$5�:||��
ǚA���Gj�:9���4�O/�2�}��d�k����P|u���aż��	�D��9�5Q�'���=��w߇��~�����LU��E����Bm�T�'��(�?�����c�{�
���*�4�h:3��n�˘V�<���\׽��� �9�U�	��K]K��I�=9S�OC�*�J	򖯑��*<|����'�	�"Ә�d{z���(�o]����Xd&����&P�8vj�s�$p>7��.3&$��:$�<e���u)eͮB���O���{1P��D�q���d�9�@">�D��]3����LKkpH�eP��(|����^dC�]l.��O�U����__��S��)es���ɄPL;|F���pB�o8��zF��~����!��L n�"�b��k���$���C��dI}}}^{�5�Gj�3g� ����{��I��g,�SV9���:"a���I��d�V�7�1
t?��' !Fa��*���n�۽u�I�4�{c������x��zg)��©,i�j��y�Sl:��7O�v���E�@b��E�������g�@��}V��	t�#��R4�~�D	$ѣ�>���x�8�ܼ�@��ja��w�Q�����!S4u�$S.��mn���k���a�Ïa����1��������W!�1�V�oށ������o���Czsw>���סqx��$M�@��D���=����$�]֨�E���˽:5�=�CulƐ�9uZ+��Lc(�[V.�8�w4Vs�?�IkH��[_��7`�Ϡ}�*t�\�W��.�?~ Gq�/���j8=�K2�v�2��ȒC!�m���-�{�����s|.���	��L���T�Y�
��\}ρ����(�x:��F���
�`AݗG����9�y!��p���>T"WF�5X�}tdn�g��A�~��4v�����OT<a�	vw�g�P�權)pu{�P���_�1j޿���SPڪ�$DmA��l��R�|��S�UJyJ�:��Me���ŋa~~��ݻ���,"b�$mK&8)�J�s�ȹ�9�1s��0���s?vP*$Fbii�=��K����YD�Vi=q�FD�n\����B��)+(�Rbk��SFu*�Y��2�n�[ت�TO?F�m�V���>��V����9�u�T����`S���R��<P��' m����G���f�8�c�Nx��?�l�Ǟ����n�mR��e����H`�w�^w��G�� ���P_8�5��.߀��翃2V�k�h%�Y�֝;p����R3i
j�6��{�!�Gk0���L$�k��u|��y��O=����	�N$p���p��Ƿo��4vq��]����޻�8���g˒v�"�I}?����mdx�����[=XE&f�B��䣟6�����;��9f<��0d�Jl.t���9���g�/�{HC�R �[��o/ɘY�P��vͨ=e�:vki���5ߍ)������;�J{Y�f�zHc�B�Sq�N���W{<U��\�&����sӉP/ߑ���L�د�F9/���a�R�������څg���L^�L�WR[6U�><~��4��7a�OOO�	������7)�j܉��3���!�u�a%�C��m{5;��q����T�2�@�qRgϞDПwY��T��l���"��a�U]���%�����P�����Nu�)�+;�=\�.�;�%lx7�s�¤Z���̅\ȞK�\���|l���ѣ��X�TF=���'a��K��,�޹�*I�dO�C�+���)����)�,�I@�+��9����y�?�4Ξ�9�u;J���bg�F?�=�X���n<zp�۩
{�S-t��R?`���'{52Xե#P=v��e�7&�+�Vqn�?��W�߀���=CW��K��D棿����)k5u���4)���������CȔT��1TY�48���{	������9�;�&�LR�:��e�y	��U<�]��D���/ʏ��:E��`4������?˚3�,VVL��]������{3:������OA��0p��+��8��j�J�R�?���{X�< ^�F�<63zm���4��E/p}��lG���V,�X�G�P��[�!������WV�)�?����P� }�;A�r��>{�א��.n���!ٸ��ƍpA���!�v�:����9vl�\f7Z��">�ԟB�-�O簤�<S��f��Z��*T����{��7����`{{��tZ(�o�����V��L��Sڥ�N�D�ָė��� �S�q�7�NVg0Jz��l�����T]M]�B��B���J��E�]�Cg|`�0,��
L�=���JmUQ2^��o~��d�`��Q��5|�ľ5��Rmuz �6Ղ�9�R�;�c�_��ٗ^����A�Rt��pr���̞8�v���=�"D�t�^%����ف�V����3)�I�Zv��ٮנ��쥗a���#C�Aƍ��I�=~&�)�B����'����cD5��8�Ub���!�4�򶍷�&�\}d�*33p쥗��w��:J�md����9��t%�4�r7`�<�	��%�� +v(��e�C0�"�'f�VR���A�_b=Ċ�F�B^"�����9ɖ|�Ŕc�
����b{�.�����u�aZ�~P���������h�2���8��v�����L�g�#��By��m%8^�R�ڠ�&����=�I���.
�������SC�4G7�������9��Ea�j�]�.�"�®���av����[�#�h��$#,�S��I�o����o������.c8�`Yr�r�q�'Ǥ�qI��=I�=x�XO�>�!d�o]�S'O1������$�˒���� j)wJh.�a�kx>1��~��Ο�ٙiQ���	�u��۳P���`�Z�s��T�2�}-�VH�$5;��D�)�m�)��%a[�h\�p�1_���5�.�|5a����\��R�6J�k����s��_��o|��N@w��䬆m6�'a��߆��YH�o��>��8n��+�X9S2+U��F�1z��k�P;rf_|�~�O�q�,�+5���`�Y�s���o��kX��C���k'+����ȑ�O-=_���6Ҟm�Ec�H*�z�8��?���3� �I������\��^����,��~�{x|�2��8NR6K>	l�A���1�⳴S|�f�ƛ�����������ʌR7Oa���qF�&�C5#�N��hP�6*�J��H[�sU%&1�A��jLB�>�����E��tfHs�����:�Y�-�[����J�c�L�d�SݾUr1�8_�X$�*�(�[�"�
�[1ٗ�r�7�s������ő$���\�d3[��T8Kk�^�>������S���1��2�{�DR�x�g9�,��!�
Hg����>v:(���y�ڸ~��}ử:���ڪgZJ��8��,C�ǈ�)<�|���������=�����3�ލ��Fϝ�ء�T��𶳱��{�v�|�7a�JyV���z�*ܾ}���宖�r&��u����2d��>�����8�}vn�� 1�;�m����azf�=�I�B2J���Y)���5�h�r���>C	X�[&I�J��係�ukh�g��f�Q��I�����p8�}F�M�g`vyj(�N`��Zz�8��yv�{I������:T�_�����O/C�꧰~�:lo�B%'�:� &*�.=��"L>±���`��)?u:�;Y��Xc��y#/�_�dj�x����}~6<���K��̅`�4PZ�sg�~�$�N����3\ֵ?9mRq'��J�n�`�M�@��y�O��.,�̹�޺	��x��6�)i0��#�dr����3��r�,2>��=;�	 RNy
��iX|���%��qo �w�q����đ�P��$���G�6NN�k���FF*9z
&�UН
^;=�������ʥ\Ѕ���Lc��ƌ�-���I���sͻ�5F��Һ=(E��6#�y|�~�1��`�P�i�ߩr�5����~��=r-�*���K�ӿe�����1bvsR�o��qܭ��H�a�-��x� M'( �2p@�6�т�������m����l�m��������?�co0�}���S����*w�ED�	���ycc�A�"ٮwvz�ǜT�t���נ��q��?)��ϥ"	I��85��	�Ç��2��O�	,.-�fhuuMb�7����|hN!�h�w&��[޺��e.EXT^�)w> ^{�$l*��`^�~/B@��e9�G\$�����D�IY���HRJ�2�,_���^�A*CI�]��Ի�EI���I�Ҳ-C��@ �8y֏�Gs��#��q(�V��#}|�^7�4,]zf^}*x]�@Nj��#1�OfSJ�j*Ԏ�����`��`�a��`�<��6��ېS�p�OAr��	X8{&dd��3��I��CƆSUs� d�Hݍ�b|A}l�O����a�]�ǵ+�}�l�?fP�!cBI�����<,�M��2TΞ�\#�ʷ�J�fb*3�p�oB��M���5�#�ns�P��þT�T%M��ф2T'��&Tw�0��T��.�:��-L#S4���E�C� =W�s��pJ@k���y,����9π	Cl�y�t����0Z/����]������n_����{y.S����Ib0�뒊r�\�UΤ��C�=�3'(���[�
q];��u_�P�	������{�s���~������E����~?��
E�='3�|�A&Nf�amP��9�����7P��2�=|��3����7������uJc]EKj�D��a�<�ur�;��7%�!'��o�ׅ�+������@���?�p�Vk�o�|�n�Q52�9���c@w�Q��]?�T�N6ӥ�r�n��N6	G��723�m���c��N�vn�I�����t�+��nj�d���"y�ǒ�Ɠ�ʌ�cي�p��ej/\�#����S�(A��-�s��H�[p�(�V�m%�A6% or
U
�KɃ�Hu��Y��^�Y35h��
B ]��`���=\��U�c�ž�Op�ZbD:ĸQ
\����d�c'2�	G����U�#*�E�yo�K}�#�{��i{h�q|d��� d�	h%5��8��v�˩�}|�K�b?�-�Z�P����P,|Jq�x�*�#1�> m��R۾�2r���~������r�4TĿCw�rT��/w�D����F57�S����{,f���r�'*h�h$�+ب����^��}�^�?���{$\ؑ��cuI_��8�Ť�u�Jo֖�7YJ�@�U�&:
�K�n�+��-W��s��)���|����6~����'ר�tŀ�e��n�)���I�QR}���� SX���l��ae��O`L�^	l�:[�R>k6]�L&��f�Y�S�r�Z�ףca�������B�����^eg('o[��u�Q���1�<v�?b/d�Ώ[�0���j�u���2�P�&��Ȼ�R����;%@'�1*�B���`���/]�
��$+�M�|�9W���M�=����
�LOB:9�&ДS��]{-y��7ք��ƞ���PLv����
����8�*%�����PG�vl���a`6�/.��U�ø�E�c��9���)�JF�X����D�\i�kr�~�ȹl�c��/�V9�[ǠG��h�W�,-��F��&�ͅX�q���Q:W*�nu�ޙ���z�Td�>;��-����0�4���(Eq���p�#�rf�y O���e�[��8 �=�8��%Z!$Q!o��@+w?�P�qb�z�χ�{�)ΫU�,���"��c��+#.P�J�د}عe�<�S7jYr_W��T���/���C��� x�����p+!�x����`�T�.x��½{�0<��r߆�J�gI�n�	��Ҩ���C��Ij^[[�n�n��Y�H�4J�d���$�<zZ�" ��� �V5\��m�JmT������#�@0'�z�H'�n�r�C��T@���)k�h�cf������ܤVo��H���nG���;�$��H���$,̭�?k"\2d���;{m#�?��āy�Sb�tGPIfҔT��"�>S� ��uE5L�a�;I2M-K��,�I� ��	����	�X[��%ϝB"�(:�O�^#��'2�dl�;�Z/�Jz)ǀ��R��T�47���MK%�Ds��c����5QxSO��J�1�eFe���?C���Z���bщ��P;`�����8�Z~X� �26�1- �Q
��KĄ�i�W.N<獺�j,�$⋀�����U?��at�{X�f�J홄~�cp�A�Ɉ�ep6�_�ab�e#�7ޠN�)v(]<��l���	K�K��_|-I<����z�}�����J��
���~�_���
�_ SP:g�{��u6E��5���R��3�=���I8}�4�����;�Ã��Y��S��w��L�c�"�ת\
������]�R��>1�`����3�C��ٳgarb�K�P/%u�H��&K|�4W�a�6�93�J\�٭;���+\B�(2H�8r��P/�_Nnֹx@�$�@WJ��� ��p8���
ny�ʺ0+�E0��[����z���ʨJr}'ë�m��N�'�V����2*f��BeYi�(�i	R��뜴N[+�񺝶H�8��/����^rg?&�z���I�s(}��wԉ�����p���<���H����&P�?%��OL&ezs5�Y�M0[)�˚�$�C̼���I���O�(��Ԣg��2� 9k�|,L��6l�h���S���%�s|�dY��߿��1�{�̀�d0s�7*�~���rX���G�X&L��H�by]	�G����:ۑ�-b	�wI�Ĝ��k���L廌|�]�܋]������i���(
m��s<�����vH;��#8Ii�\J���4I��K��ȉ	���ѱ���y?z̒;��i��e�#u:]��x�Ն��mx�M�S��v��a���u΢�`����=}�p���'�1�ޚ�s�Jx�Νle��P�g��e1��O,I�y¡vԀd)�dn���w����/2ax�g#�pF3���s�(_:�pe�̘;�%:F��15}Y/F��˼�8�)���0Nka�' q��.���qU�8L�f�*-j��$�26:3G��Ĉ�<��t�&��1�g��F�$���C�T���_�y�e����������.���km�U]y^����'7������Gͱu&H)��e��z;4{�c���pk�!��+�wR2�Iil?I�Vk���ńA�-ƃ��'�|/��@t��= H�z��G����R�cn���
��^��s���Fz�����s���4�x�>����#�ߛ0^ʆ��v���!��a����s�vv�K8�`�I^�I�����p�&Y���&�����2�Qq�6e	�b�)�����>)�S^�ԩ}��K;��ϻ]g�tP0�rL�u���+�qs��-Lxb�تI�C̈_��\� �߃���_��'�۪�U�-a@�Sn�޲�ڙ0<�_2�O�PH*f���Cǳn�
ˬ�s1�X���x�§<�DQW�������}�晝�2�g	����,�;�W���?q`nX
�p�5	e�8���O9?f�+?q/�M�Åe�Asf�S�Cz�ع�Y*�]&̌xa�F,wcbYm��L�W��6i�zv黯��6��ˣ�k3H�z��]�3r���Xa1���wL��"��x���C�G�?K�Ӄ�r˞M�d�z��$�� ����W�:�Ns�����4��0u|����E�6��TU�-��M�q|�@��TZ�c�
�*gms��������d�3�ot,b>�}o��7:����@l����hӸ6
��m;_ϥ�_���ꑋ����U�u�RK�0�f�'�c��:��Ty������H5+)_�	���G�p:���i 8Z;$��LdqP��ڭ)��^�+q�F4	�u�>��
0����>��zNQ�%{�2I{՚�p��%�!u0jA������I�ͪr�.e���.H]�;ݞS�r9��Ʈ:�mt_R�S8��J����O�M�l�OҠ���]����" �Pҧ^��,^�uh��?.��c�2�GrD���]�J.Dec���3È�I�0�b�g�7śӘ[	���*�'b[��C�
}v�˙1N�1Ԫ.NĉM��Tږ�'�01�,�H�?aډָ�H�4��|d;���Z�%�8љL%h��ԫ�}�]��\�=!&�r>���v����K��p�SB_l�]�e&M�ڎ�Ѝ�)��c$5E�r!�� �{���P���Pb�]�9@?�	�>T�#���8�RAG[�d2������9���×{o�_-��t���x^�)�Ulٖ��{q26���]t~�s��V���}.�^DNi�ٲ�>��>1SS\� ��/&�v�W'�:y���}���2�t���}�zvFs�j6J:P&����c��.?�3)�j$�Ӕ	�w�7�c���^4ʰY��vsg������Nb���	���H'����΀�
��f��7f/v����۬Ar��(�� �+���� ��γ����Dº�V�-$v��+���5A�9�h�.1��*iJH�A�qI��]i ����3��ԍ�0��e�Wu�`�yh�~g2=~sϽOw����tf��>�znť�Յ!�Ft�_�)1~�����9QG�IBk�4�ϼ�r���D�G���>#I<���s<���v�@��r�N��=w�*z�p�W�֒bdb[V��ϣ�5n~8�r�C�y֨���+�G���{�c%�]��D&fduvq���F��yIZΫ�y=&��K������q��:��θ_2Bd�G�g�y��g}�ק�����c�׼��,y����L��Yr|˝4��K\zH8�Al�t��fM���(��E����N���n�]�IІ�4#S��A~�����*��O��,y���᳷4I��\9}.I��+Wa�4$='e/Q�'Nq�e��|V�������b|�3M����$,m3�!�uS7�p�8Ɯ��9	����T�����ݼ'�-M<Ca�sf.�D���.�*�;�0�D���p��-�V�1���0�7ru̓\�J�7��gE8�|pϔ��U�͙��b%��}^P�&E�h�N�lYH�k��lrr� \�=�:@�c���$��*���g��:�Q��9z�����=~���o����5|�����R�%{�Z�7�k��(6!&X�j�H9�(n����0���0|���d� l�}2��]��q�"�y
�<�aSis�fTc1)A��06L�҈�
#�j�0���ޗ���9�=Kї�m-��[�*��p-'!�>??��6H$/���~��֊��Q��K�~@��H�2gC%��,�<x��dl��0-�Ť�Z�#�!�{|%.]-L�Sq�Ң ��b�T�T��CVCkF;�;r�%m�xV^J�#[]w���f��fk~�W���6�3�n���Sn<��b6�z��1��	W"�M~��p /��*4Nb�����<c�����sյEߑR��Pf<g����w&K2�4�)cf�*���u}�ê��N�����/�s.�?}�u�s&	��YI<ḤŎv�	2	�������+�O���U����$����iw�����k��b��\"4$���Q���x� ��b�~��/wE�<}?8�P�'X�ٯ!jxe.�m�ҤϜ�!����YMgՁ���gP�Ǡ ���[l���W:&�ʸ���`���Ȗn�T, Tᣎ�w���s
�Û��t��`'����i}�f Pu]X�x��m
���+z��WE@��o����L�6T�6������lp&�'�#e�X�e���sM��#gm�Oz1��U�"���5r.#I��ӑ�>���H���_euK��kJC�֔�=_	�4q�p��t�C��j=��f�%�F��f�<�xiW��w��ǹ.7����˝Tj�z���X7֠��W�Vq�9�P]��lVc�0���Z�~�E����i.8L���e�K��s�<��%N*��'��S�_�kӏg� �G$߻�<��\�O�Iܥ�{��6�7%{����.��m1�d\���iyO��p�g���_��
�b��$֚	�+��B��ޅ��x� �[�M�;'ǀ��"(so*��o�R��fC�c�7N�@�ka����ʝ$��NB%IG�p]��x�I�@�'��i�<����~�8�4q�HO؃w�H��9�J�
�%�L��w��S`r@�C���1�y�q�lM�ϼ
��W��Qbc�D�1w����!sw�Bta�>ĒB�n�������UrG�����'>Gol��t(|BmC_�s�I�ƿ�N��k��y������O�x��0}^�ڦ��
�j7�g�3y�GA'�\���y�U�HMm%�嗳����=��q`N�u�J�6�ˮa��ɻ|{s�^�Ȓ��՗�P����P�̅��d�ʽt,E_������xm�6�yP'ƯJ��������{pt+@���][�N��ERt�J��a�J�|~9���c����p/���{d���i7a�ԩ7�ݦϠ{-w�ǈ]@2��c�6!����U��i`<�6�i{��D��ҮXP��z�K�FRD�ZS�瑱4��˧���}<��t�8<�9����=����/��|3��h�wpcݼ����0��	&AcN����Y�gk#�$��:��MV�d@`Е舍���5/�/6����2�dRbo�!�m���]hR"U��� ź�%BXl�z�[����@I���{-���{.S_I{��UѶ
P^:?V�;�N���;P�6��c}v^����(33V��Lt�S�>0^ђ� "��f��^xv+�[�㚬��U�9	�]pn���Y2�&C���I$�C�S����F/,l%�����?��M�Y�T#��I�T����W��:?}�f��	|���%�gMlŭ� ]_�����Y��������w.ܔ�L���H���~������}�wΠ�� iGjY�s�s�<Z�F}I���5�:?y��At�����gJyx]b"eʼ@b]�9�W����<��Ud�\���б�=l��e����(�]s1��|�tNA��+bi���{��H�S�����~e�-�R���nǨI��{��ml����;x��#hL�8{��jv;���&����{��ɿ//y%��wh)�m��<H����jO��V	c���IC�QO� ��IB$��/�P����
������x�b��b���#��F;���뤼N�=�q�����|G�>��s=iȪ.�� 'ͳT�8h�>:�F�$��q�a�tN%8b{�.��9�<��_�)ּ��@��S�U�� ªQF�E�Uʝ+ zξNB��v�y ��ǀ�C��.�W&<e,���I#$j��I�&zV�^�b�q�^BN�.�i�~��p�r�Oжt�c���3�}`͈d~7�~��QU�V�,�*{�d�3R��W�tA�=�w��?(���(��5�&|��']vE+�G%�c*��ib���x� �f�$��`;̉-v����H�Ü톪�ql�:�w>�t�>TS(�;��-h�9w^����r�F;�*�t�#8�h4�g� �i^;�s�������F���\��'�l�=)Hձ�;V�������q1�]`z���b��b�7�/�!�mx��p�sx�y��p5ah��g���;�t$�yj�:�k��_ܽ�rq�o�8������ 'Aj�p&�]������M%���[0KQj`�"�ǌ�jxq��\���f����V;Z���n�;gc0�Ԗ�s�N��M}�7@���3
cL������Z�02�&v�5Ə��G���F���-����f2�ʼSq��HM����t�T��mc�E�c�� D�	Q�E�n�9Z$?Է�f��:�>@w��� ���·�׋�2㻩�Gqx�4�s)�P�Ә��6�\j�z�6��z�QK�7����m���8IǏKa; ��yDJ`
���CA~�C�$�?���=�\��#�>e�NLt[��M�H����ItN5t�MLA@C�<��mڨOJ���b,m�h��e�(�rߌ	e/�?fpb�[�¿5�i�n�y���X�b�1�8)�sϯС^^��f0�T9��ߜ����HT�2&�C�`뺦�a��P8X���Q�Ж��7?��g�^c̾��3<�K�\���)  8F(Lb%ݪ��s�]�D1c�ʝR��t�H�a��!O���ctl0+�&.^���
�6J��5��B�U�� �|]�U��H�zC���Hz��(��R�������]=��/�4�h�>�:V����x*����l"��m��GlC�&vS�奄����	��ⲇ�:�ڪ#/Z����u�WLznD�yt͐~���A|��W�s�a�1�(tӠ�p'x~\��hq��ȟ��ѭ˧�B �p�� lܦڠ�+=.{19�+v�y�S��F�B��Q��0�����D E�噩#���80�q����{���Y�ϡ/0b\+��2E D����5�R�u�ȭ��uV���GUg��t��\���m��Y0�*�C/E{�V��1"j�ְVs-4jW�8i�ށ����*i7������c�hl�z�c�|����13Z/@}mL�&HZ���rƺ$��	�Gб�J���_h��4�����kd�d��XD]ࣗbv�*�f������t�|4�:��ri#=�K�|��1��%�Y�}��g'0G.�
�ZкE^�*�(w�?�OY�9�" �Q>��D
������̨��g��L�&�NY�%6��{:�N�X�������-^Υy���%�}rf�խ�:�>=v�9�<�[p6a�NwJ����̌��a�9҉P�+�G���W�‾���zۙUL��#�Y���Yw�`�	jbpL�>����@�}��ο	?[�����ɻ�9���]��`���Ǹ4�ƪS�cH������g�: ���Xq"�]|�	N�a��e����מY���̂�;�m,<��*D���JP-H�ZN�kձ���A�+�!�f���Aχ�Bχ}�<�.���\ ��#�N$_Sn���_��x"�S����%$R6L�R����G|��1ʶ^n;��[����e���Á��"o���!� ��B��� ��*Y�
��C����9�y���'?G4$�&�u���@"	Ƀ������i��ď+�x����~�����e`]C��<�j�
�[�C���Gy��Ii<���8�[�]Rpwߙh�D�dh�����[����|\>��Ú�L檙):�w�2h�8V�s|&0��/�8�q��'��
�fь'
P:�.�_3\��>��?�M\��8� �&l�)�6XWV�'Q�$̝��gn�W\�Z��#F�j ~.� cc�����H��=�?����i���\D�P�3���k���0 ��A-A@�b�}�;��ɳǪx�K��@���I���V�#"��7I�^�}�:,#m$
��9����}���{�}���[m ��U��a�Ӽj�?��A2�Z_�*p�T�M�T�J��]��\��Y#��9pOĸ����{/"�Z���G�:�w��:V����Tt�ϰ.S9�!���Dݦ��y'���p�	oR���������ה��ܔ-��Pf Bq��,��T�+�c���7)�(~@��/������_�ݏ9Lp�J�%AP}@�`7��������(S�x�i?�W����R��3}A���>�$ė�->���@^������ѹ�INN�u� &��z�R!�/ T?��u�#q��LW��0������m ��|���\���߂�H���-�^�d��_���!�����7�$7���]1�Z*5�#�/4�.�Ͳ�ks:�:@G�C�y���ܡ&�P� >\����W�z����T���^-=�t����qq��+��kɗ5�j�
}H)I�-�_G)��^8���q�:S݄�F�W�D��*�5�<"��lwr�+�¡�Z^��Jg�mh`��5h��y	�iw���~1�.KP샆����:^׬��o��%'�d������v�'�1* IJ�0ެ��x�	-l+�+������ǯ�����6������\V	x<���e@7��/?� J��%�9gb���HƏ�(,� ��_?�������sڏ�Q�E;Z��ț���-@�����_��~K�¯��WǴ�)��Č�/̇~������,�Q�F���p̈���ك$2��]��8/���˗��cY������d"$Z2�� ��I�7�KCRL�d#�����@���,��K;e���{�)��vy�$���V�>�����uB{%c4t"��g��E�Vnǩ������fc/��0'�a�A�R��h�;��ٌT�O����2��$ЪXD�~A��3p��8th	����������݇����t�
�!���gl��n����S���� ��т[wV���F+Oh<��PתT�
���� ��T�r�>��p�;~�j��چ��� .߸w�b[U����oօ:�������sN���,����:|����^�����V��ݝ<�9��w_���0�� �l;T�;�� [����ɵ[�������m��H����^ש'���4���N	:�ӑ�����(�Y���m���v�o�-p	)a��9kW��{��Ե���B^]� �G��?Z}|��U�)]
N��.��3�Skw�1B鹶^���� ċ��o<`��wCv��G������<D&�Kq�/�̥����[|���N�q�k���!Ϡ��Q-�s��tm��ǝ�8��x��DK�(6��R�M����U�^��g���<zN�o~
�r������&Y���SRb(���3���e��%#ht �$	��5QIV�n�����\��H���#H�Y���d���_�?��~�s��X�SX bЗ:�&��h/�fL�P�j�g�l3��vq�&M�BT��XB��l���Ⅳ��Ԁ�����bx{kVW7�Ν5�q�1\��||�1�ri'g�Z��Ff�����&���i8s�z�l»߆�܂�N;���ڭ�*H`��("/.�·^^<w�;�f桎Rz�?uj������l�:� ���&z8q��x�4���	8s���h�ǡB��zplyN_�3܂��}ֶz��K��8ql������c2�}���3a���]�[����C�b@�Usc�u1�H{
~�ds1�j����iL=�JI3�-$C����'}X��+���7A�T���@�6x�P��̥�,/U3f#A�>gB���p9֍�ބ�G�58������K���L��j����]���lt��C�&&�0d;'���`+Ob�~�Ѧ����*��K-�<�q�^�+���z�*�����30���[[��M��@.S@�g ������F�&V��C���at7����lm�������qsa�.U12
92�}�r����4%;���'������){��Zܔ�;
�Ww��Эr�kK�!�*�mY��K���X�59h�����=�ӧÏ��;���3���Bk��j�F���U�յ>�|~�����{(�v�Ϭp���*1)L�U�,����WN-�x���ͩu�f�P���)�f&6n��M`SI�|g����4���I�W�����C����p����p���p��1�[ZB�>�� :�T�^z�8���Sx��C�rk�++����<3݀W_9�/����Ã���?��ȸ��b���'����kml���&�3- �����F�(�K�pk*M%�!.�%�<�H��'u'䕐צ�K=R�i�8a��i�2�NR��p9�>-n|/�)�ǀ��#��0-�*ߺ<�6����b�T')��������wZ+�j� �I	ܾ�A�������v�8ŇN��� �Qr����B
�h۸iwG�A&6i�X�/Y��i"0���ImR�"#1j��X�@;p~`Z�*�'H�C�S�{��_����$�rf%MK<`�4�];�P'L_	mx���T�
!j��qK����,�U�<�Kō�j�?}�Г�O�ӑ���3<>�lړ99�-�c����yk��T*S�`�g&����O�����@��k>�z>��:��n�s��K���j#�W�8��pse~��5��W��*��n{�;��W`y�	ׄ�� ��:�m�B���~���bJSjY�}��������,̌sI˕G�7��D ������?�>2ߩ����6����?��./�+�/�/��x�}���g��[��&��K��_��?���i8z~���p������"�Ӂ������q����[���'PMƘ�������N�v����{��!cS�gh���,TsM��!����*��!���e� Mŗ�6?9 ��T��H� ��RG�� ��~�׵�~��U���R�ˣ��D�u��)�\��<wt���F���aR�%M��@_�"v؇a>�f��n����DD�h{/��m���c�x� �m����РUM�X��(D�Љ�&�GP�V�V�o�ORtӳ`�ILkoS�� Ŋ�=b`���q�s�2r���s��k�?X���G�S`�B�����7�h���O�{jt��C����î _�����Q��6��3r);;䶴��v5Z���N#=޿�t~��r�YDr�w���l�bX�'z|M�R��}�T-9:�K�H�{p��#��ށ_��]�x�^�7n܇7��"�t��O?��w�C���rAS��>����.�=1�z�,�Oա�ڂ��LMϲcPZI@�b(�(!հV�rcL�z�߁�1x���n֠��7nޅ�pVo���+p���p�|-M÷^�v>��@^ǏW��O�pH�/~�!�����ȑ���|�f'�Q0�47(��>9�%Ь'(�����?�罎�5Egr�Q��*��`N1��uţ�𤈡U���J�qL\ز��
J�K�r2[�w�xM����$�ML �Tc���
2}aX2v��؄��P� �dF�+�!�Ʒ�(J
QX��ӳ�=��Q��I�N��k�]����@Ć`gXá'#~����Ь�HL�|;�*�o��9���
'��0A��$͘᷁��
D�	�D}6r��@ݬO`����=���1�h��}l�{vW��h�ݘՈ8���/�s7�L{r����w$(���oi �1L�C�O�<�G�0-�qU��Z^:�xz,{O~�W����3����q��QV��������w{�oT�P&`v>��)�ъ�ڮ"�O+ݭ �4Uh�N����+p������xjn^��]�ݷ�ރ߼�.�|�(�2�U�{(�[X:</��g���k�WP��B�9!k�
;���
xME����U�\CTY�����	Cܼ~w>�>�F �{���r���CX:4��3��٣p��
���;���۰�q����G��g�a�Y��ׇ��=;l���C�Ղ~��*�F���^E�h���@�waq
��n2 ��j���Y�"�mw��#W�닣4i�}���a2.���S�':b8�	��d2�<�cY��-.����4���P�ϱ��^�	�NNj����:>#14��>2��$�ЌU��TMD�$;���$�hd�}^(�O�Fu�M��8U��u���z=��+���%щe�o9{��N�"A�o
�zG �a`��1D���t�����>�{�2��h2���";S�qx^+z?���+¿̨0�֥�5%��!qKpڌ��lUĚ����2Qn�ƛ@;G�P��wϣ��$M�G���iy�9N���P4��Xi)�-�P[�#_No��O�9F�o�I����7>F--N$r�J�����Z�!��)�V!hH)C��	H�M�c�'n�玟�o\zvV�������ނw>���?�/� ���PlՅ�I�L§��)�W��_�w�uv����� c�q���s�'⽞T�ܿ���F8�<�!��7�M��k�83	�)p��d$>��
�r��$���V�`}m�f��Y30=9��4�lg���mx��
��膀�0=�}1p��	x�sphn
�kUx���{���AcbjubOj�ur赻p��I��_�Ξ;�z����ـ�����o?�^�*T��{D�
�q��	D�C��(��D��B��$2)��K��j�!�U@�xe(�W�:LN�-�(Y>Ī�G�߆:'��]�UZ8�	yj��ߓ�?v����~���.���KmAr������H/�Hؿ:i5��tҳ��*�P"�#%�<4c^P�k1��S�#�VI��J�d��} �#���� �&�`c�P&�L�g��f��-�X�ώ�
B/��`��No��h�����З!���o��6��F6���AZW#�����&��_Dm��}�����]̥���6=�%���pE/�Q�0����7�2�HWM����x<}�ΙRG�7{9�=�c��RA�V9�����,�l���I���[��3eor2��[ܺ���I8vx��8���s������ ������r�sXۢ$�"ŉC[/�x��O^�7^���t��*���Gp��)8w�yq��D,�e,�Pq6orP1Ul�Ǜ`vj
��P�y��m�(��n ��$��4�����>����8�Z�9[J|z���������g��	8�4� 95�������'?���uXE��B����&���1�&Π���4LLUally�;ֆ��L������X�걳\/N:n�ņ�묂@��kf����S�� ���W�^�7o�ւ��h�,2 Tt��Ds��c���܉Ç ��<x����g*���ӆ���d$?	b������O�&�rd3�T�;�L���'.Ԏ[�}�J�^�TSO~]��G�!k��]���A�a��7�ky�#�%��w�����Q7��󽔥1�%�bW�ۈ.$l`��E�Y�.���t_E=����8����3&�����	��jc/FQx%Àcca��������-3%� t��t=~?��V�����yz1	��f��ζd��Rz)��W{<}�#���a��P��͐��I�	�f��F%V	<��
2GIb�r��V>x�
,�V`j�(�V�#���G�Z5�Z_Y���݂_��H��|��[;]�;�@��&2 ��_� ���>����]�q�.�al�*��eg#{13�l��E�a[���l4��4K�44��n�z.%�w�Q��BO y��Z�)���xIevn.]z	��ݣ07��*S������׿�5��Ԡ�'领`>�����A7��8�V���;03;����(�����|�0\�y�7`4}yO�P�D�QJ�5�01��=_��Μ�{w�!��7o\GI>���Q�1b�z=��k�@g{��g'&��>AF�OR:>�i6�d�ooA���Nok�N�%c*i��=Q�ك���ݥF�@�7C��>ŭ'�� {"Y@��pD×ny��TQi�޲��"V�G�EJ]1й(��vt�Ψ�6�����>���ѝFt��V�-�-��MG�����B�>���%�LL\C׷�ـ���lm��Д�"��e凋%��/Eq?�z� ��՚��l�04N���K���X�{)����&���{�uO!�SfJ�>�����(1���A{�������X�k��HZ2����ݜ=+��Iq#����O��Ûp��p��qX>��^�s�	
s�f�p饣p�����������Ç(��������.��1�ݮ�O�������`����N���64�G��;'� �{5q�c$�L��G�x�c�H��M��Tޡ�9�e#z��1(M��������-O��l%�&�����^z��?�~���G!q�\�݆���B���M�|���ؗ�<�o��<��������G����Ga���Ǹ&��MfTr�H����M]��`G;�盧y"��2.5d��S�,-߻}�x��f<�t���*����Q ��J�U��)����k����.v�nOT����I|$����+������OC��s�k���'@��Z����	e�Cަ�����n���9r$���@�S(8�J@\~2>�M���ﭐ�%h������>�m&�r�6�zx�Mg��Ҷ�a���8��� }4�o~/{��yp��5.���R܆I���(U�뚈A6s�J#�%|aĮE�*0�qW���v�>�i=�-���Q`W���/��1-���R���iR�V+�>(�<��t�&�Bvs=v�'y�5��a�'}C��#��3��D�@SVZh�[�ɧW�1�¡E�����LOT���E8s�(�����4�^~�<�=\���=��w_��Q�OL��{�m�;{N�H๋�ajz���U����,��W }�'���+��w9�-���#�J�]	�	3j�:���㙏Q��9�I�Vˣ�ݺK��
���Y��欭=�?�>�M�`>��/��O�s�����X٢,v��������2�|�2
9��6>�C�vv�P����~}���p�jxwd2X�Ჹ�~F�J�j*It��;mhuZ����V����4, s�����j��LåK�`kg��ir��s0T���[;ې�d�W������F�_E@���g�Bp�2=Y �d�R/{p&� �V�*���#Ĥ������"4��
z�D;	؃�"*����ʇ@����;�2���~h�0bK��"
0�z4�o	�U
/�5��?^�>�9;K�	�p�~7���3F���B�^'���z)�������_|!���-�#b�
�<�a�l���0s��if�	u���MP�}m>JN揂#=�:@g��ˠ>4Q@�3�I���b�a��R0O��Ӱ�(Oy.i
%���^�@(�ѬB/��������>�A�r_�p
���+pti��u�9?{�8|��eho>��^:G�-@�tc{�������,-.���8���R�9���;��r�jI�c\v8Rr�Q*]Yk��N�c�iߏ�O x�#0]Ù뱊}�l��-�����ن��*T�M�o��Pz߆�7W�����k���+ga��)�o��"����"#����i���}�.�6;�l$x��-���!2?=�6�|���Ol��l�8�K.9�+i IEN���z��f���MMM���!G�}b|�]8[[��@lC�{A�ل��N���7aeuvZ;|���2��`a~���7n�6{�'��2�B�؉�r�ԉ�l��Nqn9咹���בƄ�j-�M~&��(\ذ*!�:�58��&=_z�Ёt*]����!E�J�z�� 6|q�b ��Hb�t��;M���G�
@[�o����l�&����5��\��+@�h��f|�1����hĠ���^ .:��c�j���?�2�^�-1eJ�|�d�
Q�R��
x�o�-ܬ��@�-kE9a�Pg�A`���O�5��cG�,w���bC�p�Y�ځ�QE���-��cs������F1}s��r��M\����BݔVsC��r;��H�K�}�	�� 9Vx�����%����?�������
7�܁:��?����8����C�ZGZ�J�k|���jg�?'��b�4~\���!c/���|��#��v(IC�㺹����Ƨ�h�`���c�qu-,-�����O~�;X]� �m���<�NWv���d����߃K/�ȱ�o��1��7��?����ާ�#Ot�e��~�q���
�8~�]���\�r(=\����d�%sJKK㸽���SH^j�`%������vp��0�0�F�%�*����w���v�������}�G�>txVWWX317;����`�����?�Ϯ^��2�܅u<g��QX8�����㻟�q@,�y��׎�I �F���Id��e�n�Ÿ�ui��diW�j�Um����%o�7�����=W��~v�q���c)�)����M ��SO{�B�0X�N~x>G���q���ޡ0�΍�Wl�Z�@㠅�T50��X��K����Y*w9~2��K�� ʾ+�)�(���xԡ<c�b�ر*�-"Ӕ8�7uci���z��{:+�����}W����1�A�u�3 60���Wއ
'ޑI���Š�z�y�0�>9{�̱�*��p���I���A'Vq��9�=Ν9���@�cGI�-��f���&d��*��}��3ج�א5�6dr���ޛIr]gb_D�K��^���� ��(������s��6��#{l�����ociFG5�D H"v4z类}_�*�-"|�}�EFfe7���>��HTUfd,/޻�]�k�y����~�/m{a������6����I`n~�d8}L#���-(솆�=���g�2�HHI�da��o�qϟ$�7-Bmqa��ԋ�����b���o9�*O�˝�r�:n�[��,w?�#�*`!D���H���?�����:6ַ$.��e��	:{�8�;Yܝ]��c�Hw�q��8�^!�ch��ك�c���K��[��;�XXٖ�yT�'ON��'B����x9�.�q��ѱaR������A��X4���N�ڥ38urgN�ct(���~�ʋ�#E�8R�.�*�A����M����%`�d�m5�R��@V���-�%%a{kKnugs���F''%���"G/���Z��Ã��=95M�ҋ��a��xG
�d�o���Px�jO"I
��ԤV8��==�U(r��bE���W�LM������^�Aб�5�i�5��2V��H�<m9;~�nߢ�vW�눠�T��.��4+4�?&LS�pط�E����nk�-7�`�5B����ג���
���.r�P��
�ʕ��
~� eGl��4��\�m7y�ܢ�z�2"`�yR%�RD�x�;��kE�3I�_	�JQ��ǌ�s��C"G<���AVx��$8Q�K1�8���}��d"�F�C94��JUz��x\��cg�9R�y�$$I����\��r,^��X��#2A�+�����R�j��K�[���m�� ;����ԓ�Qb�-��tw��=��G�#~ꭝ!�Xc��O'ki]�jz�����5ǎ[�E�9~�7�So�̜���߿1��惹e�LN�����e�״�ZCʺ�:i����+8u|T,���^<�?��G�(�0�ӍS'&�&��������&������tt����ٜ�]W1lB�������$ H�pLzg� o��1fg���ْ����h�3f�Ǳ���>}���N�k|b �x����H`��i��]��?����t��;��%l �uw�����ˠ#����0��G�H#sP +~+��t)1t��L�0�ہ�\�փ�'����1E
ĉSS�am3�{�1;�N�^�廮�s�L�Վ���F8�*���HX�Pm4EWG'N��鳝���EP.�	�7�A@�!P焷�c��^:18<���N�H �no�H�������q$�ω���[%aΥ~�\��<}_e�{ښ���W[4�s��]g��y��� U�����nH7��c�^`�*�S��eC/�(D�O?�����n���QS�U�A�8]m��*���;`��ߍ%�j��+KN ��)]9q��R���C.�+�CY�Y��KY�̘��<�[�=�H%r���1R��Q�HY[Y��Uw:B�h=�2����CqR��4��$���ׇ�R	�0N�A���N9�H:Fs�C��H$*����̏��C:f���>��q2{aR������0 �:Irb?���Z��knE\W}�-��,���n
Uʠ'�����>+/��q�RIs��\��ظ�=U"fy/�qw��6S���x#V����.�nY���A��kȽ��a�[�,���q����7��,���n�ٯ+���51hS/�wCd�U�X���lD�)q�.-��g?�E؊���Lwa��^�$"P�w�z<E�X/⽛7�h}��(��lUZ�^��_U�\"kǧ\��!��K�:ܛ���.Yq� p�5�,�0时Ȣ���/]Bww':���ʫ�E���;ՙ�����o��7���n	�w>�O
� �'���'0�#�D�P7_�,�4	˕���x������먖=��߽M��"�¹3�R�?؝���M���~��O>����-�m��zg 
!����'��u=-�HP��zN�y��kr�9�1&�@_Og���r�i�C�u���bu}�� �>����&&&��7 g�W��\�P��7�{ۛpã#8qld�3rN +[��X][��a5sI�cR���F���E�p�WӅ#OB,����E�hnpI��z]^��F�;�8��e�yBq� (qVOB�2�kK[Nls����x����V�(��DL������o��с�_�Y,m�I��de���4>!nxr����C�!e�
`W��~�� �ּ��icw������h�y�h���������������O� ,]'�bx��������N�%����ϐ"E��o��ᓛ��w����b{7����)�fp��u���oX�adx��5��Z?ocm�.-���8���DO�e�O���Ņy�I�N]8NJ�Y�<x8��?�X\ΡXRfK���H*O�c���?p4���a=�dH�V3�M0�B����B����.�o����,�#�MxZ� ��y�R[W��RT_�hx5����@�����9���t�ʲ9��.[�]����n7��c��[��|��4��Z��{�U����x,��u�����V.`}q�=x1$�6�xXb���!����&�|nu������I�%Qʚ[G��-�0'}96�6
��`��4O�����v�r,*��Zm{������,~^��|��6�W�&N��`�:{�#���r��`	��Y�~�NjD\⇹R6�J��YRPzz�d������x��E��3��hs����bE�sU|�����&e�����$;U��-ְ�]ć7�ca倄RL:���XHuH�LY[��&��hcc��$��� z2Չ)6�dDz��\JV@o�T�6�6��fQ`W9�g!�GWg�Į�MM�9�]��}��g*g�������j�_@WO7���=$��H�q�����#�"׬� h�D ��:��X�m���w
5Y���{v�:�����+� 3��-C,�9����>����u�.e��c�X���c��M��S�= �,tT_�5��0�bYՉ�g	�:�����T��	�Rqt]��̛ y.j�r�k&=����ɇ�aJ&"���emc�#�wљ����r!�T| ���ѳ��H����9H��z;S���F
#�ofvI���p��)�Ɯ�����E18�O�v)�u�',U(	Z�I��+Y�j�"޶k���0�G��X4DV~��=��b\���W�H翐��7�L��X��^������)��������a�d2�'DH�s9��7��mr���ޟZ|�7 ƭ�^kƻy���sY>��:+���73�%�� }@�����ٟ������o�`0����h��yp3��2CM�va�0�)�gi�c��*�(D�]��:>\����]��㤝���s�z�`�
X[]ţ�U,���B�j�$yJ��L@� �-lq��9�v�d-<��Y�d��e	<]��=vQ��*���MMlE㒀��+��~�3�wajl��'a�BK+�X!Ks'�C4�I�&�H@���G�XXXŭ�Cb)�:b�H'eݔ
�g�>}?_A���ETr\<��5����nv�M�#'��B�+[(���P�t-)���b�Z��X���ǂ�R+�e�A�ƒi!��p�67OVY7|1���'�ɧ	�`���_���ȢΓu�LG#�>.����FGF�RK��%T�`�����}������R���1���G��׏����pu}?{d�0����~����4�Ṭ��BWT�5�&�y�`����hW�������;��!�pKY���YΖ��2�9���/���#V�����{��$�nyh�ެg4bW0	r>{��$����Vt$���4ӡ
�h�A�����t��Wv�<�A�Z��3�`֫'��7/
y8��R���j���J�8 E������={��#	�%��.8Wp�=g�y!a�ysǎ��и�L`����."�<r�2͛2����mfJ��D�"��(r�)=�S�.�[]���"2ɬ(�R��$F���8&�b���C���gd�y:�xc$��C���/3�AY��M�D){&�� c����?˄��E��"y\�� v4 ��<��?ثl��W�b���o8�e=;�|Aۋ
�~�Xk���Z��8xޭ5����sU��y�E��� ����P��SC���t���(��v���[�_�W�)�na�"�/��^''A�'���$���*�I�Ϡ���K �O�RS�g��bU���u�d��)F�#L���qi�y�g�(�W���!�L~$��,sC$�z�$�lU��W.�՝26s[�{J��W�27����jIj���
g�G�B���+b�TU����z����	��|V1QS�.��X@����L�<3;�xz�=���$`�Ѝdh�z���!��t��('AMNL#K�{gk�ZQƋ-Nb�ZY���p�OбΝ;����������UT�E��@�.Y�{��8�qz�'N
���l�`W���2 y�i��[���	Ӡb�c&~�b)q�٪�'Bb�l͆<�\�m.�;�-��={���U���qU�(qkϰ�慴���S�a�JP�c�X�0i���q��⮛5�-w�{P	���&U@�����w�"��_��-�:�DBIt�������4�G�<{��.G��E�g*�$И�lm�Z����HA��ￅ��~�J�h~d7vi��q��Y,�f�uqW� 
�CX+9TiMfKt�;UDS�n2(�5��;H�����;Hb{f��ƅ� O�z��/�1�8̻��"�6�wK\۝��抷1�h+��_��ml���Q2=fY����D8v�s��<+Uʙ��3`
�5�O�`���z��
�;�mG�UXI�9�L�UF���~y+�L2���?k��n,sV�"��Z�T	ٶ��_&����:��q=�Z�����)����p�f��Zb�Z��;SBY��F:�ՕE"B�����l����丨N|b�հ��5�t8�>]�#�_5��lm}U5Q� L��,^�\2�0����H�R�Vն�RN*L�Jח����ʔ#�ch��T����Ե�����.�x���N��/"�B%$[����Ss-��m;�F�q��s)�U[��ډ��m�3�uT�����O(�=���t�����O@�3��jQ�n'Y��e���2	�ޞ~,�,c� <GrrR �{�/��`{w]۽8U?�$׿��ӑ�s:�%M���`@)\�xu�~��uL����/��S3�NA�d�oH;�=�ֹ�j���,��dNoqS�ntBX�K�����bU� K�@ƍ�^���(��qB^Mu��K^�-QG�oݺ��-;�JT'S1]nLW�{&����b��œ"%b�d�6���*�=l���#/nx����*���Gݺ�/:W�x%d���8�&)�W�U03��˴�lKi����Ǯ�D�h���}�<oݩ ���0�S�,�l�������G��X���ڪ���J��r�	ubO��aV�빼qs}M���]�GN�d0ڣ9ơ��{w�A��k�[��$��E9��� )/�6�E?�1��kJ�Ҟ?��q��ih��8~r%�'���?�KE���X� 	�`I��	�����ኡ�5?U�d��<C���t�=S0��fkt��.uC�!�bʍ�J�T<K���J���'Va�^U8$)�Y��"�C�2��#��Ֆ���4��<e�[��q����:���19N���Y�C-6K{����h�H�g��-���S�<�0�#1U�X�Z���`�1O�9��zjK�s�
^�l���,(�pL��g���=V�/@$�QG�Z��C���Ġt��	q�/..#��K�nM@��#�|��j�&�i)����\"u����c'�hv�b7����s�ϣ��Wj�kt�$h7v��s���2	n>.'5q	��%?�.��`o�K�/�ı)��"�	u;����Ъ��m�7͝�Ľ��v_��LeK��9l1�&��)+2��ɇ��D�S���	�.~���j����9q�{�'h�Ɣ��ԹrL�1� V���X�S]����/{���*��c'�q�����9��Z��LlN��?^au��t*s��r�r���'��;Z�PE�a�W��(p4"��nI��Ƈ{U��@�po�Б P&�憄�!�Q-P���@w���g��<���N��nMYa����cY���p����wQ+�3,��C�a������Xzn���H߸�O���C�=G+�����3g�T���!�JҌ��_�(��SĠ��J�|�}*<]�-���>X��U
����z6Hoͫ�z[��R���8�QS�.�R͕X>y������	��d4���r�MY���& �t|����I��Y���!,���D�Z�KE�� ٝi�c�Hf/$�
���g�VhljPQ�r�!�`KL�l���<q���bb�y
l5����ZU���G��D���P��a�8��/E��mjump�t"�b�t��U=���Xr�2_+/,�b$���Y`UR�Bح::Wy9��j\/�Ԗ�Vj,������ݮ�Ss�/���Սs��	@77��D�7}���##C��ȑ�]")Bכ�'	`b���BOO
��XW�XLy�� �VW�T�H�$F�W%�Y��@�����ɪ��䒸�$�1�F�-�Ԅζ��gO�"A<���\��@,Ĵ��V�M��eaULU{�Ͼ&ʁ�1�T����c4���g�����k!nFzш���rū��$?qbYMB�dC}]�H����� �IYYXb��[��yb]�
�k�k�&C�s�lTus�plzΝı�	���)��-���U��\��^��+�J+܇3s�{�!�Ò8�����_X�L���9͂�~��B͆~�\��c���_���ax�O�h��WVi*���J2]-L�ɚ��-�����rc&7Q>���q�ʽ��Z�H�S˄�I1�8K���&B���*9�~�� UA�Q�Ui��E���{P���+x�O��(s��v���b�:v�;�T	�V�(�o]0�n~3AO����<��b�O���t7� v�7j����ϲۖ0�ʷ��z�&��װt̓�8[��N�����,���jH�����mh�f�r�>��fE�᪚_�|�����:~��*U�LN=t,�If�ᮑ&M�u4 �t$�Хb�"D��ĕji�N~��.{�]�f]x�k��UX��C�tF��_;6=E;��\���-�DB���D�k�2��u.�Ay�$3�cYp�>��\+��#�w5Y�0�o2�B1�A�����
�н���H/tn�s�"*�&	xRd8�Q-�<�wO_�bMc[X� �ɭN<���F�Q)H�X��ΖX�ʅI�cתIڑ�4=~�Z�gbI"��� F���ד�<�7w��l|N�b7�G���U�v��̘�-��~q�Jz{MVT/]<��O��x��c���+_q������y��b,����󰔒�_�1��8�4}Zí�>�����chO�냎+����e?6���|��Q���5�������$�fn�~�!��V\�,�l��IY�N%pjj�C�m�or�B���JѨrݯ���
h2�AfOȏ��'bR?���a���T:A���W]H��\��l.+G	���	w�ʤ�2�L7WDМ�k�V��J�T�P/��a``}�}4�P�s�B89=�ٙY�'p��	Q�*���O �H�����R1[H��V\W��%���9�Wc��
��Ma,߳�֢�N����*?��������tK�����o���ݠ�6Vz���6<tV��p�~���� ��jr�<)�L�9&����ӥB*�'C�IϛK�N���c���$V��d�{�U�����y��j��Ԓ�f�!KYq�xqt{T��QZ������Ŷ`X}�MN�DݦʌW��iFL���`>1q�:l�T�B�
PU�U�:�Kх��$"aۚw��җ��Q���*F7vq�-�Z��c�*��3�_���d�{漞�X�Iք$��XA����#A�3�H��axl��m,��b}y�����>:2�Y�\d�p̜�U�2l��E��(�=�kX�J�}!�R>G��C�X���'p��1a��en�L_<�����4!�.�"�I*�uy������L'1��-��ǦG�:���% )|����s��s��V��Y�4��j��V�N]��c+�z���Nt�(�(	���k_��enW+lw��c�Y�?�)!B�v��g]EE ���ezU��NT_��Ѹ�q����������S�Ǌ_�xl�*��X�ܺ�q+����K/M`~�.�_���|�"��dm��P�q���mDw���y x1U2?�8�G�($��\������Ρ�#!��o~�	R�4z|a��+M�C���z(��˘��*������$��ɩal��᳛7	�{��h��{r���1M��>u����0#�u����^ܻ�1.]����=�L��St���X���7��`���\����҃�w(���%����<aqnDķ�U�A�Ơ?���L,]In�LrQɭjЌɣtC��kV��SK]��[-o��7F�yO�C���^���M�`\�V�b�K�^8@�Y��}�K�����[I�㪃?݁��'3��V]Nj����[�V�������'K���܈x_]Yh��Ik
ԅ��e�+� �H�)0��ڻ/ֆ�����^UdR�CH�h�-��0E9b�qy[В5-��TB�[35��
��y9^�P�eM}/��alѱX��cI�R�)�%W���*E�Aݩ�(��1݉D	`-ծI��{��V����zm*b�۞��M�{�"����D��������"�7�1{�>�׶04<�!��~�}�2�7����,�n|V��9���v�6IX��B�Ι��n�lK�6M��KWo`dr
;{���T*W������0��(W�'ϟ�8�����\</�2���ӷ�`b�屵�rgŨ��W\����ߣq(`���յez�
c]�R�1a/ATB<5Ǔ)Nv���˗�ʍKt���ɏ��g�!���,��ם�{��7�I�\8q�Y����˿�r�)7�Y�d������m��U��lo����Jp����t��2��|x����]�*�y*��AwG�\�NVv�������[��?���%�v�u+�k�8p(���\i�������`�)^Qx�*gIBJ��\͕RQ9IT+dE�ܪҽ�i?C�
\.����"���RS���&ST�C�ŝ��>e�*/��*�Uނm�=C�Q��4g�-�/��z��I)�$��%����<�2�����N(��1bl�j���2\�}`���/I��"�i?�-j��Ψ3�BC��c4��y��� �Cs8��>��~v����н��n����%j��
~�_n�"��tjjMV)�z�y�%�Ǚ��,U����B*slj\�Y�����;D�0G�\���0�'G��Q.�Ľ�E�_��0S�?Z!aI +N�12>�4YI���A�@F��(kW����k��3$|ϝ>&�{�p33�ҁlzr��=&��Xȓ������
��>=<HV� Y	�y�����:sϻqy�H�������p("C�h@V�G��gBj�\K[F�Q��x���5Gl��Z-�L����g��p�1���G̯����Lw!�V]�:H8v� ���m��77��
B��S?Y<ɔ�A�i<Y���{dA��g�l����%E�CV:[�ӎؖ�ަ��8A�i���]���ĝ��25h'��I���3,,.�\�G�c2Oqz���K\8� ������Q#ƙ���,�dd]ܽ?��3����F�p�µ�N����w�}�ܿM�q�BR:��غ=U�*5D�l��P��c�����"@Ə;M���)�99����6[P�M��T�Uy �ֹ��T[�J�Q\m�g7�V~L
�b�e�2���H_?��w~���hak[��ªI�J�ӊ���$��p%���9��^��>i��4�����U�4�Y�.����T�h��<T���2]u�M��3�ߌ�Z�� �^?^�޺�@]��7�ǲu���V��a�-����1:\W�?kU�b�@+�ሄ���W���4n����r��o�>�7�#��+�p��0�a�k��8�?�S����y:���9o�|�������j4�5<��a��w�"�B�V��d�6��L�Sq�t�n�|�~6��w�5jV���S��k/�;A1����E|��\y�,Ν����ۘ�]B�����+��;4���9ȪR��D,��2d���Ep��s�/��mtv��˿����If�k_���o\G�P$���Nf�6HP��$+��c��o]��t?�����/����[W/N�_����.�ynU&K�Q@�.{�օ n��>���L`��С(f�=��<�����t����k��J���g�u��S�!+=BVy�����{� k}eyU,���Iq��uS�2���թ�H�����Po����K����5��e���4�a�Dy�(�X����Pd	{����@v�q˅f��vH!�3���0���ƅ�W'!�$(��,����)�ǧ'�?ԁT'�ՃH��ol���F���i^F02܅�qT���*}�Y����r��2B Ȟ����v4wܚ02����8NLOatb�x�p�sҜ	���J�[��4�{�sE1��w'dD�#����y���z�t����Lcy~.^��+g126*�asg�g��I*���E=���l�^&�T,˟w��^O��}h��U$Z�4���WS/v3�q��`�{M����6�<�v<mP��]��U	~��
�p�(H�*kS�pg�D�����q͕��[��V3 ��'����L���fXƣ�5�����q���}�IE�	��b9�A��f|�C}�g�W��.�i�mX�:���6�сh�D�o����Fvq|�w���_;C�3�����5���9{��z���`~v��w��{��k8u,I�ى�{���ޠc�q��I�$��#]U��r�,$�8����Ξ��S�Un��4w��������޾E�h�,t�|��"���A�����x�װ�nꇟ���Ūd�oW�S�d�緄�۾Vku�.�ሦq�����W����̃����SB� �|�VE�j	Z�\�/mW(����
"d�sw,i+	Z��JubnnV�ח7p�w���NLOM�kw�"pN�K�Ktb|\Hf81jkg&w����V<� ��i,8�]�۩�q�2���te��H������k}i�RN%/Y��h��'�݅a�*��.t���nc��a3��'o�X�&���?�W�"����Ӹu�)�E��m�$�Ù�uW����U���ZbEsQ%'����0�]M<?�R�M�#�V�y��4�bH%�Б� ˭��t곸���]��z� ��Y���t�����d^X��������P)5R�U$)���_�歏�o������y�B�����,}��Dxj�q�=?+�d1Xz�=����ϰ�2)��4k\,[74{�j�H(,DJ�\���x�{�0G.�3�D��ҰzRz�~ڝ�[�h(���7گ���jha_�����Y�����|I��nAm�Ȏ?�d�@��R5�j۷�� ���O����w���ή��eWu*!!�893��xp��6�����+��H@�B!_��VǏMX.��;d�������E)��S�t��x�Tf}����D@��={f��@����`:�|�@_ɚ-dQ/�`q�<N�6я��.�l/�$��X�{������R�8�_�H�%0���s�/aqeFRւ�R �oG�Wܕ��,��k�����><�
�C�9���Q������2���T�,�8R���{�$�OHg�=�vs�C��f���X��d��AzqV{��#��`��a:�~�@,)!J�\��FC�b��5�����¶�%%quz��_��<�Q1���^�&)%�Iɚ[\��S��u�����n1Y�ŧ���9��FskmsCZ��r�F$��ir�P8$����>��������0�]��T��./�|�&n�"31��<&JaJ޸̃T"�g�Ș��u�CU��O�����&���W��kk�r�ku����S�=�i�}8���	9�Ă��5̀7��Sg���:�,g���tv�%Ǆ��d"L
��C� ^,dR@6YV�a�d���9�"�K6�U6�<3�-}�fâ��lw}~�ҹ/�D5�Q��!)cUV�4���,c�3��u|kX{���6��� �?�V:��v+���0MX�B�"Y,]��r��2��f��X���P�S)�G��xʓx�[o=N;PV.���}���FSfs<^`���
�jl� �0w�t��aqq;�C���E���IбF������D"t�����p�a_X�#������bd����0N��ǃG����A�\���gET-+[J�� ��ӹ�plz��nn,�ıA:g��j��f���<��o�� �YZ$h�2��I`��=�>z�s'02܁���}q�r]��������&&(U�ƣ�%!
�#~ş7�������ބ9<��� ��آ���s�CvoQ����xR���t�b!GJQ9a��DOg�@����@����~mЋ�wg���$��Bvt���2{/��)��	�c-�yz�2�A�됪���x���J.�0���R�8����||n����@����9������2قP�`��E�'-�Y��/����g�=>���͝RZR��J�<�|�ỳ�������{�4���9��|��>���y���霖ъ�*��2�)�}=������X̻[;t�.���+(^yO��9�*[��J%$�q��t����OJ����������gh�E�{Q�}���I	�Zu|��7���K�ɏ��!��V#����U��z��f iO3?�{�j�#��$��Kyh`���=���V�(x��%4iͺԔ�zTGL�H�������EU�T9�R���X�z������tN���tVy�����k; ��Vy����׽/����С��t�i���툆
���}�q����D���D��[�J�����li�`f_h4��[w������Y�ܙU�,�z� �,�j	�}1|�_|�\A�R�֦k���=�+�����l"�A�x������!�"��1,6"�)�x�+���zKK���"m��)�g:Ed2۸Cy!ǥW���o��7޸������t=����������5TA���n�Bh�u�?��	Gp�����wHXƸ���к�vh��?��\ӏ6��A3<�޷��y���פ�	Y�r昭S����@<݉8���#���)��S(b���}!��;I�p��;vˋ�X\���ֺ���B&p|��W�))�Z����m:	���-.��`��S�6g�mSF�JȔEĠ�[����?� _�%�>��ҳ���w�u��?������S��:�5�twİ����?�P������o��-Tja��0�����9!餕=��޽U����[��W���6�������I\��2���7Ⱥ�{��/�9�]�2��a]��}��G�}� ���(�c�_�F�)�R/���R���E�e~n_{���?�:�z��[`����8�����x���bUVk�"1�գ�+K�#�L�Q,�i=�{���&�B8����ر�g ���n]߭�7&c�#� /�q��z��`�>��K��$�e-�;���мt*�U�$H�ܧ&T�a��h>�DA;����B+�M�6K�S�2�:��{k�G�6���J�%��(���e�Gt�1p_���:��9u�f#��E�|��'[�f�؁�� (���nކ;LMp.+���'t!R�RsI��,Z����M�Xzqi�����t�Y�cX^����:�6����Ȥq��М@�,�l�&��b?��c�D83;����	מ���op��������*�aph ��O��qQ��;�ݾ��j�z�'OLJ����iD��-�E�'N�­;�$���+��B�U�F�5VW���ɭ�kjOG�m��������П��_MP�׌����et��@@�����h��0)��`�w��LZ� �?��,�;CY�	�њX޽}����%+yO qaiE���DR�lW�p�d!W��ыA�k��ܬN�[sTsN�s]U����T	8RIp���I����ֻz���>�#��B�Q�`���|κjؒ��$�?��F�&]Y��@�o�`}s��k���(jt�W�����5��8qbCct)���K	Z�\S����܇zE~M%��[�&:{���w��W£�]d�8�C���۷X����/���5�inf�s2�7oޡ畧9~�0=�*7�y�AN��vi�W���X���?���8ȕpf�w�������l�]�G�3�|�zB81����B��~�C�Z��V��٨#o,e����G1�߇t:!������a����P�V��Z@�A4�dp���y`[ô픁Ǎ���4�ő���еNwd�ysu�ٞ7���%oO�P�c~�kXZ�� ��Q9�X�t[:������f�X��}i�cdd�p��/_�7^�BB�����y!�`˛c�++��|u��xwo�/����	����յ����b�.^Z�&e�Fgw?��I�"�Ճ��q�0:::��3 ?��.Z�E���Y=��� ���|ai}&�g�����x	�8���E���ފ�1`��6�hv���g��T�ԥF^M��_�yf�p�tFI[�f@g�f�Y���(�'�ǈ-9�Xd�9a�bo���0�;�0I�2L�hia^\���}z�4^]%嫦)����,pϒ�xΔh,
���ձ��^�(OK1g���"�ت�M�P�������Ʒ^���}�֛?���J���[W�nĺ�|�/suÍk�Ȳ�*.�[��rp�R��-B�dZ�#F����;(��f�x��+Ҩ���G���OhN��M/m^B���Z.���]�K+8v�)����?���Ծ��R�B�E�i�,W7������v�וSǥ��;���ܣYR"�E����]E,��/��S_Y�#����2�N�aEJ@��>!"�M�i��牙����,� ����e�B�3�ߟ �^ӏ'��9���H�bt����uk���t4IP��y��f��^Cu�b��~�7�u,�b?j�7�D0=2x3�rf[˄�7A_=���t@��j;۹ڟ��Op�����oh�G��x�r��C����Y%�Y��Y�@����+�t�t�r���E��aG\��0L��Ӊ���;}?��>��.vvwI0���p�S���[]ޣs%	T���y]Y��R'����7?�T�����\:C�<|���>�G,�����:^����������������2	���?��ε&�\���o����N���E `cn��r=���,��&Y�d�E�Z���:��2z}� �~�3�z��H4�+�{��j��ekH'`�{Һ�,�j� ��v<)9 ��$5�z��K >�ׇ��~�5���8u�,��Ymm������ (�UE6���8��PS7�'��ѫL��%�	�
�����(_��|i�TTc=�7�������$y�JY�I=��U��^��w�:i����[��Җ�M��<�%.Q�+nt�� T�Ǚ��(�<������z��;��Ր$C8!�6�x�R����0�V�+����g��Z��evj>�b'��P��.�A�1ȕC�uw��-˽V�qz&��n�87�4Q�Y�	�p��By9K��C¦]�K�Lȳ�����_MVZ���dó���1mO��&��7P��l����j���qm�iL���	�:�)Q�8g$�i���ܽHX��h�s���R����^<�?x;3v���QOH{%Iy?�Q�zG�aZr7�����:ۗ��x�.���]���F�y����5z�Z��N�O_��H����`����*�j��{X�_��#��ݽ��\����9���5{.<[j�g��q@VG���;w�K�POw>�d�;��i�z�v�Oo��%�2�C��su��ʤp�5l��������
�c~��QB���L�@|kۛ����K�Gz�0/�Y���޿���u�gʸ}wk9d˰$��>�ϖ�E
3��$+Z��ab��t���v��W�/��xS�kA���k��K����+��A�V���y�t�]�I�;� b�L�Dv�g�E�K�b	]]���D:GWw�$��x2|��q���N�\�g���Tj��1;[�ꁆ�L��L�׶Ē�z��-N�a>#7�)�6��ݬ".�y!,{ʕ,#Ru�����g�J�*J4i/c�j7-S����4y9c��?W���5����h�T~��ܘ6�{����އ���Z��c����;����,��%��fU��C�����c%��V]W�� 3�1c�Y�/��7*���Fx����H��[���*����N�|`a�W ���y�s�L��PӘתe���A��m���9B���woP�jy�A[x�aJG�F�BDKϓ��5s�i������w;�A�Ya��-|S�.�����X#�W��p��x�	�?vO���gv�{�H��"l��E)t��f�+r
�+�����r�~�����D�%�b�ES�2�2T�i��d�)g�:^D�`�(.,���ܢ�}�H��q���#ݽX�JKQ��d�Y���
�h�g�b�/���>v������?�L�Y�����VV���7K�� �R+������"�
�k�^�E4��c��N�긆5����~�N��ߞ����[ߊx��
���{A�b���ݒ�
5�m,z~GН�N�@��!���j�"	Փ����0��~%wimKVz��7�э�]��A^��bU����1�.�y�0�Ƅ4RjȖk��c]��U�'��l	����ъ�#��6��ݸ_�Ӗ9�3�#��]��%�\J���h�&�"e۪y
��̆�����ԥ5��y�U���?:O[�R�˴�t}պ�w�,�pH�S��JGQs^��g(�+0\���sm?[�B1+��E�#!�����B�sY�v�E-�-��xO0Ώ|d5����l'[ځ�ӗ�>U�n�<�p�o7夨7�\�����������T{�b1/���T����W�G	Z���F�0ny�vs�T�6������=1D3��V�=�x�|�RF����sl\ hN?[�$O��?���4�=�7����R�cOA�\OQ%D���-aa
	�:�����PV�PPF�r�6^8&B()�E(+[&������qD�ŉ�" �f�f���%x�Ȥ�a�&�2t�4��)]#o�{�k|�۝	6 ����b!���_��k����X5��BwS-^�yڤD�|?Q��q1/�S8�l�4Q�<�B������ݷ�Z��� x���@}Œ�����NT�DpIa� Y�.Yz�r6S�F����ý�sd�p�\�zg")	s<<���7x�R���μ��Կ���f��ɒ�T}�k��v܀uN�Z�"�4���|!��Ǐ�Z���6�U�V�j�fb�4�6w�cϤ���������y���&�������߻�&sO��PϯN�����FW��y���u,�QS�=i�7����K�� K����Cڎ��C���tf껺/��f����(ƞTWXVP��)3�<���0�y������A�0r�m���ā�/����t|C�b)O�!Q��:�e�������k�t�O/"���n/�������3�u�/���Q���a���D,�(��c�������k�Р�l���qmMhk'���ԭ�\�>߷j�ɲM�z�g�ي�o���"�¿����
��@o�ځ�/�����Ԭ���ut-]L�q$
� Ǌ ��q��jQj�y��S��V������,I�G\�w����L#%�X+9B^�
Q��JC��R�Q1t���f.2ٙZS\��K.�N╗^�������Bu7,�c�{V�Z�=BBd)�9M&�ɖ~�Q���$z��G�d�V%��=��m7\�x:o���%��(�<u�3���{���	���7L��f�q��,��Hoq�*YءXDb�쩨�~L\±�C�d��$Rјp�Ǣ�E�WT�U�%pg79���*J�
��ľ9>�:�^�<s�6��f|�Lz0����{f����q���.Q=֦�u���_6��3�[��CW$���D���r��w��	R�t3#�Qk �ה�f�T����'�L�q���ϖp�[�)�۲��F_q�蟷�[�;0͂
�u��lA+���v�:��ɽ����M/������{���ӠV/cU%��|�,z{{�9O�Q��I�t�[�	�);�q~�ڌ\�#_(?���{h?�����@�ũ�L�Zs^C����A�:Jh�+�^@@�.�u<����R�g:?̜Unw?��^������F�Z]w���' L�#�!� �@�0_�>-n&k]�� ;%s�;��g��r��.!B�H&P)�5xP��W�zuV�fx8NwH2�WV�t\τ�Es@��bq�����*�ܽ�lfӣ=��u�.acJB|mm�|#�#�MX[����.�;��Egg
�|7��Ù�g��[�̣u��K�ͫ-K7����h�H�R��0��0{�[�pA��V �0��V��$�O�ut��0���j!	�8[���B��4~�$Y걸oII	\�3�i�L��C�H�qk��wς�}//��7�WFl��ɖ�ԛ��H�1nĵ/��c�'1��/�y�צky�TV�]�Hɫѽ��;Q1{��p7���/\�l�"rHv�[�m�r!��DP��g�R@w$��c"��HA��)O�-boH��\���( ��YB@�:�y���[S^���jo�LG�g�5�lM����������^�Ї����" ��,�:�-W=�U���,�h��u3�;�R"�R֬�D��7d���@ݸ���8j�?�'��t��jM+(y#��aj�G����,����K>x��#Z�?�l���L��fX�%E���)�u�5Z4)��?�NL�wX�?3+��?��W_���~�w"���ł����;��>�{��W�ŷq|z]������<�?�s��7��p����߾���.,����������TO��WU��ZW.\�W�rCZ@֫ELM�����"Jbs�,
[:{�{���^���8����+�W��w��>���Q�<~�����?�%֗�p��%\<wZ?�?���<iNi��c����FV'�XMB�kļ�g�if����5��*q�d���2����b���hY�YL��a��a�f�0~� �L`� �ݡ�bK�%`+e�m&�[�z����c��J��}8��*����QT[*�����wv�{=�q������O�j���K	\�e�.���ek����L�����`)��I�;�氿�����T�ʊӞ['6ʝ� ����y��+��0�G�n�*��	Z7=}��s<�� ��&�Y��\Iu$I$,)<�̇��"zxt��Q�[�G�z���X�����1�R�݃��Q�
x��ϓ'AE"�o�z��.{�l�3���V�� �5/{��6���Qw��U�m\����k���XYm�NOuu]������Y�p�ӱ�dJ��2�-��7-T�HӶB.s��K�^8@�LO����r��ߚ�q���J��qJj�R2�JC���
ݿ�jig.M��;���O��{(�3�\Y���"&�Z>~b����&�V/]ֶn-���3���˧��ʴ�IL����F2���@����˹��͉�^��2I�"�FS8{�������(���z���Vag'�"'t���T��JJ�|6���)d���j�H�#e����?�2Ν���n�- QdGLE��Ǵ�4�[�k�������Qkj�gdd���Ş�qi���?'; �E�HR���]8N�D��-~���Ѹ�4`+�Fߩ�$W�AQZR� �՘N�4�5E�ѷ��e�.`�a���<��~W��G����螙����el�~�&wD�T�� R.m"]�ό���K(�|��
g���߽7�����E�%�=Zp���n��`�U�D:N�������~��qLO����BE�곚�&�!2.ej�����<*��,sI��od����2�YͿ*K������� �v���Y�����  33}�q�;�l�5�*�&��4N^TmR�FH�U�a����<oN�Vm��s�$�N����yz�f���s�|C���"�wj<m@=�O�{��c:�T�&t�q����*R@E�Ϲ]U�	 ����y�Ӟm�Z~�k����O����5\�O$�kd���<D~{�,�u���]<���.Di��..��+csq�S�/g
���n�x�12؁O���O����x��N�~�&z{��㯢\r��هǦI��bs� !��ťC$����뫋�����p�X��$fsmkkX���~&�ʹ�.��nu%C�ރWn\�gJ�\&�����l,/�����]s�0��X�Tb�O�*i��aA7�YP4>��Q���'�����h+]i�\�/���o���t�<v/�x"�T�!P��"'��˪9��U���,�HH�� cj�{%i��s7��2h�b5�(ܬ�g�*5ֻz�@W����D�������Rʈm��a�=E����|��9��4G6�Y���=�=�ujf�$*ɔ7�$�V�o���S�� ���ёN`j��^���'����������st$R���а�t�5U�l��O ��3.�k��=��\�A	�j� �'gi�s#eH�����7p�(�	�̱�u���X��c0��9�\ԜLB ��
����x�2E��j?�9o�/�o*��W�J��0o��7	�A+�I��4�P�V.�v��դ ��^֓fǯf{]��M�p�a=.~Ԯ��W�nol��|��fHe��ӷ�������۷?�o�~�������N����w>E�衐�#�����?���c�k��O>���6P�2�rXθ��������F��!�BO_
�|�	rdU�<uA������*[���F9C=�֜,���YTKUD�M%��+�azl���㧤,���G�$������&&�1=5������3s�W*y�H�{<a�害���a���Lf�4�{-b�k�^�G��юY��DM��f��&�Ar�4��$)���y�;p���[��)z8����d�3��RxE}�]ܮװ-kîJ  ��IDATU/ݭ\ez&��ߣ�_a�/K@W)��g뙩}��J ���7��(6�X��"ș���U�խ�(B7����ul��a~n��<z�=47�y�Yѭ�Lf��|�n@#�ɕW $���@������KW�ͯ^G.��7�6VH����|�ý]}������׮�����?|�޿���uz�5=��1��$����ڮ����ʑ�������q����.t��{�9��%I�Uay*�%~�����O�&C�-)�U�#T�T�x���(��6�)V�"5k�����
?r�-��r��<ޤ�S�|�j:~b\H���ʕ����~c�?��z?7F��n�?ik՞����U�>���$����וĢ0g��>��>f͢���`�`z�>�.���V����x�����M��,�-P��,�F��>�9*]׃��1y�������{ɚI#V�R��mb���5��=ܿ;����=X���|�����3{�Ǻ���TΟ�@���ɋf��F#F�9z��c4���|K��yK�X�A��?��5�o�����J��;W���͇��!=f�]�6�E�� ��,˸�uٜ.��|�Q5�9�Vy-[y )��un\��B�{�/�ww��T��M�H���u�l����s�{�O��"BBq{c��T9�J%�� �6�C���N��rG��	��]����E��ze�K�z�Fz���!�pin�{�k�=d�z,Kd�[����g����-����NM�ұ���/nc����i�/��+&Lf�B���t���#r�a����c�ӤW�3p0F��1���[a.�m�U'ϜE�T��^�BA�W$�]ў�*���J�v��/V���x(�R��Z��ѐI�1����_.�)�]/�"�ގ��g��p^ S���^H@�v+�?�L����~�_n���b���,��c�����m]ʺ:��896�Z��>�����x��5\�p?����NY��{��.^>��/buc�s��r��<<6���	)�;̕�z�Ew_���K�I���qw��7�L�.�v�ҸaI��I�'�E��� Ʒ���KV�=,�ϑ�_��Z"���;f{#��+{�[���z��'��(�Y����uV�\6�u����H�^a��d�Y��j�zA�V��di0o�7X����x>�5���p��\�����#_�`��4<3����܌e,�T�k�ZE<C�oÚG�&L������L���5\����<D��(�L�l��5p"��
���
У��� GO�7֥4Rz���k��N�I%b�[��0-��.ʌ�X��8�n�%t'�t�!|�+/ccm���A:݁ѱq�M�`iy5����F�1��MV}�o����*^��709:�p,�݃Q-Wt	��lpZ}�:��yc�b�Z||�;p+pn����c��P4����Ǉ��v�ȕ|�X�E#H�_�p�;�Ш䲺�_�9�����O�bD�]hfI%��>�Dn���|�tؤ�
͵�عe, ��§Oz��8������90�<�Zw�5s4����s�^L@o����ۖ'�J]�-[�2k��>�]J|l�r�'�V�,�������ٽC,�m���z��|�^�~��~��@�IOLM���29���X�����b�\>7����Ϭ��KWi�Q���caa�9lld���?0�K�O��&I#,\��g��# �`phD2[�������3$0G�\|���/��?�˴#ݏٙ��$%���/!��IJ�ϑ�a�MN!s�c�@��wb,�����p�y��/E��"�Zh���4�p]y4��-M�i�aɲEc��Cm�Y �ֆ�o*9��,���"��fb�j:Zc���D��FAP��Z�H�VA=&s��v+d��oL����ʻ�A�Gp���r�{�2D	��D��*�AB����\[�F�c��2��<&0_�)�<o�G������	4�8~|
��,���Y��l�)p�����i��T�p�����X��y�Jube}wfW�*Tq_.d�h��⳹��bn���._�w��m���۸p�*.�9����X��E\�=���	@�dZ ���mݜa����X� 0���i�)+�1.���Ċ8{4x~&H���%�?�j���6k!A������{����X�JV�b����A�@ϰ���sP��t��i�����.���%���Ih�@~_r,?�����E�ϯ�`�$ܯ� -���)+G2�Y�Y�G�nm�>�$�lŪ%qtW��j�xr���,!�cd�f����=���e����.z�.�BB5[�bf~;{����2�[�zCCH��|wf,`vn�S���,�P(�w֐����C��T����8�$���3W��63�[X��|�|�s���7?CwYؤ8�ju�ܲ��gK���*J՛������_�ם؍���^UuU���F��� �����HYgt�f���������	�����s,[ci4�F��(�� �X���������d��ވ�/2_�[j���������X��nq��m�sS�n���a�5��=A}^x�$\x�|~��6C��R��I���.EG���-mz]�K�!�RT@F��y��Z�\wG�6��h�}�E@����f׌�v���#���6�&�Wrĺ���_.�G��?���ȕ�Maq��c-ܼ�Hr�gn}��|+���o���ε���[�y%�Ç��=�
��vg���oa^汰O����:??皧�17�(��7[J[~�>|HQ��'�h��j���"ϝ8
g����3�[8'O�������'+���j�>l���:�ܼvn+Љz[pnm^Px�+�þ�X^|�ΟSB�}x��L[�R㳷���iӧfTM�\� G�g���6+O����3����=�aa�ϳO����U��4c9�2���V
����J5N����[�ZH�wN�^u�n���s��켓�|�Zz�>�Cyy[�Xax� ���^�J�c�m��"�6"����N��$5��f�h�Ś{x��$��Z�`�4�Sl�t�fv��Y4��?F�ĭ�tp��O����}8w�0?��N4�q��Ҫo����p��
�p���Wú�@��gtx���S8w��TZ��nߺ��a���[��)������� ^ڀ���G���A30���
��|�[���������¬b�����B�9S�a����-����gJ#["�&������@AA1��0���~���t���LZQNB�R��PM�
�ח�����|�F��Z�yL8��0��1+�v�����Q`��ß����4��y7"��c���5L�oQ�$�J��Y�?��
�����{����4g���+q����D&C��ʂ�??t��x�?:���M�X[���S���}s�	�Y��u�͓Y�ggN@K~<�4�%}���Ғ5�ŕ�s1UB���6�.=}��V���0�R�A%��y���S�3p��Yx�@{K	��4�{�G�?����w���[pY	�o�~���P���[�2��3��Oc���JI����z���:��������ڼ���ŕF��j����yPL]Y��f-%��ܗ�0G͢����^W!�)�5�t�ܽr���?���O����I|FX �["���H"u�2��9"�ysQD�߯O��<jıu��]�	�[���։P�7�)mLX+L{��"g�s:�@	�ӝ��$���O�����r:���S�T�Dp2���]�MfjP�iPH1mH�D�:״���*���Ҳ=))+[�oL�ƺ���"�^|�b��+M1z:I<���˷���U:����{1|v�f�x��*��Ōx�=UZ��$�e��f���gsw�փ��V���<U�K��y�.|:y��ͤk�0��3%,��۩�y����}�x��{?����k��f�둙45Q���ڦb:��0��zk42�3��If��%1�I�>-��Ƥ��z���m呔+�!��l�@B[�$Y"�;�	d�������8f�e8�G�pb������>�V�B��d�z����Jl�Տ�j��7orK�		mQ(���b���&"u�V�"�1ɋ~6�r��Lij�����:|��U���_U�~]o@	{�aG��g��o�@4g໿�-���I�������{qS�%�KG�Z��)8{�XYلO?�����3̯^��6� �����5W[JX�]اʮ�����*q��24[7���o�E3�2\z�%|<VMTmŃ��Z�e�&����(n��G_j�.ʎֆD�!�s���Б:¦�}(����6)ɀ6�[��w��"��:����R0�cb�H��:!5ɪ@�u@��G�:�Aj�8=_=gM�&�Y\\Tk$������]
�=r�8:p�@pnv����=
g�FtX��N�&r�����G71sL�8��\���v�P.G�I(�>2����Q��ov p^w�v�\��nڃ��$K�0h����ژ;�loc�]f�E�᝕�*5��=��^�txI�1�q��
N4��i�IYi��]�G�+R�p�~l��I��H�(�w::	
c�Β�H)��۴�A��P�����]�z����ĭg$��;�Ot�Ș"�;��v���9S�k��!�-����ܑ�&Y�%9t��r�?�v��9��)[��D��&ߣ#6�X������x0M������tk�W�:+���H G��hM���<s�@0B�1,�L�D���d�����i���n(0��A;�Q�Y���E�J�d[�&7����8�3����k��}�N�ɕ�����c��s��]4������{
��;�����|�޾I[�^8w��jmeV�6��W_�3g��}��ɣgp��g+��XО��hv��PlHcz�r�/����ɣ��ʯ<y�-]���V�~��ix��X|����Ok)�3�0�l�<x�Kkd�B!ǒ�Q:�5�y��B�/:~d�b��ߘ����]:c�G��h��*�[m:ۀ�@�T��E�͆Bv�h�8_{������;�����f��M԰�Z��N�c�L:h$aޥ]X؏����4'��h�{8p`����~��m��*��Ş��֍[�
����E�mCOH%q�!k�0�)b�;X7p��Pb�0�x�����O�����S#�:ۗ�@⾐��	�~��+$VD�Ij���iQF��C��d�Vjp��ٺ��\d�$���qt�����Y����lW��fkKi�m=�����>ZxH���>��ٜ�ٹy�}J�Ef�O�fB�4�MEi��llu�&��>#�W�z�)�����yX������C�c��ӑ��墋`uu���㶷�g�`a��l�{�{~P[;� ���� ��-LmŠ^8w
N�>)���*��|�$a�{�����h��R�ܧ�2�N��<l���In���5��ST�_܃ՕuP0g.iMdh�����Io�x!�}��RA}�^��̥;��h�4?7��S�M�w�p�턴�xzZ�Զc#|��]!֢�7)��Y�`.x>�r��洵cu�� �oa�:)����%(?��1ܺ�L��W_{���}q��߳jn�U���U�����7ށ�����+�9� ��;�x�*�PX�V�-�
TV�X��Zk0� �m�������xL{p~�*P�~�,/>%�I�v���GWa��XS�gͯn�)�"�H9;�1�~a��s��O���cy�7_gJ�_����y"��Ss��[5���������O��:��)JS�����б�c��4�T���k1�߷��/�gL����<X��1/9�o�X`��Vk��V)A��8�m�AO\�,Oh߹������ه�JH�"˄�Sz;-Z�?z@V:L���
y�)����L�U���c>�#_KQ����"�9{/�3����8 �\5>J���z]��
��YSݺ��UTޙs�Y�L*l���:i�F���4�S~k��@�L[1�%���R`{��ax����s��~��U���+
�4��`�����t._�
_~q�RlR����p��aZd����r�*ܻw����g�W.)�z�ݸ���g�x)�c�u��f�5��:|�߀o|�]��K�˰_��w~��p���*�����}���(ft��i�W�/a]	}�%����`�;���.�=~�)���*�����_�~�"�ݏ?����M��<K̬�;p����gp�~�E��o��?����)F��H������������9���o���w[k�ZPNg�^V��G���Lg��&1h�L6�3(K����h�^G12�TS5����C��/(@y��)�����Q�3���!����7�A�����#h��h�D����v����?�9	�`���+�c'���- ����ƶ�K����y��c��ן�~%�>x=Z"�x$�t�|.�|���V[������~���p��c�6�=��@���qn���m��>�z�[�j(V���;������$��R wo\����`m}]]�B��w�OTK�o��G@{����e4l�&�G�
}0J�Z�JM>{}��'C%�vT�]5�(v`"���}p���ƻ�RvēG���C��
@U=���觋�p��Qؿ?��E�?q��?y�ZWG���p����/�}芛��� >5�P�Z7�|�+o���Ν��ꫯ���2	�J�~�����7�x>���]�i��l�G����?I�":v9����:o����-��gJ��X��]%��/>?�L��3�s�3>zs�"�Sę�|�l]��ꃮ��a�s��jNE'f�'��3mCn��LW���Su،gc�}KqdRO�\ɘL�;�[����6�L7������|���������1���i�����{	�߸�O�=����[o����L �I�p��߆��v�g���
����
Џ+�u���~�+*|:ͪ���V+�����đ���)=t���Wa���;W)���Sp`_f�JCH������o|^>��|)e>��W����4����)8�����򗿂��֔���	ܹ݂���ûo� O��>U����4j�/�tF�}Μ:�4��p�����gO�lK�Q�uV	I�T�Ο>/�xf�f���������+o*�� m�YYi�����ٓ���o�iq��Yx�ҀϮ܁/o��&2[[R8rxA=���&;� _y]���k�m	�6��&���pHe L���}��B�;s�e��J��Z�y�2��PG������b
#�p�����9Z1�����S:I"��)�$4����T��J#=�+]:b��3c.���g�h�Ȍ�z�,�[p� �U8�4�EJR8���7^}��ڰ���ϟ�G��+a�*t֖�勯��s/�g�]'�jϷ�^��}30���˟�$@�����h��T���{�q�kO�£���5
HSm�@�ڴ:776)b}uU͇Cp��ax��O�b�����wU�G
�OS���O�)A艚c��Ru�A��z��yx����ߏ�p	�zW��(ƾ�<3�z����#����ϵ�Wi���Z3�����Cj�U�"떖���FS��^'�Iȥ��L���V���)���	)��q.��~�/R�r��9G�>��M��Ӱ|9��׬KK��ݥ�.UO�T	Jm���?tL�� �A����c�E#����l@U��hK����H��F��=�q�mE�ҡy''jH���O3��SޞJ_:���{��F/�KJ�>�$������ųG�w��U%��+�e��)��^�,�����kJs���]����߀��G��G����&�U�����0����'�~�їJ���v!L)���KJ�8vHib����=8����K����
<?�[�nþ��P:�f���;p������
Ig>�\<G��'�Tu��-�SJ���x��?��O֠��~J+[__S�t�~��y����F{�Au	��|TZw.\8�췾k+��~��g����M���ET��!]R�a��Y�I)a�ޅ�'����?�_}����~οx����7�TϞ���/�7��s���7Hh�~Wo�T�fJ�H�IB�ǏP��	��W�U?I8zx�:~ ���`y��4Ia������(`�u�X���80�'\�2���pr����"���3xK�<�KH�=��@��5݂Y��%�a�b�0 "��4�g
�����6l=Y���2�ir��#9.�f�ڴ�\:�.�S��X[^�#i���.ܹyn\�����}�O���u���~�%��7�]���8z�843J�N�ܺ����h�bnX������f\ �
H�+A��W�8�ӧO(�� 4���;Fp_���<T���S�ӧΨ�[���M%Ь)�� �3�K. ?~�|�͸I���槧Z�;`�5���U%�ޅ��z[=c�L�}���r�+�J�y������uf�E��VW�Q|�����)��%�"��c<�՚"�
����캉��GB�G����u�Mʗ��4'@����Hn&zztff�s.�VA��ΧQ��r�|hKtg?���tv���穪6=�K�������d*ԇ<�Q+Ч��c�����@�����.����:�7��O>z�����8~dΞ>���9��7�ֺH��g�^���߃�o�G�-����7�3g���r>��cU�&����O)-V&����E>���g���᭯��G�)bK1���j4���.\|���=]Z�-l[�)�-�[�\��+@<U�ꙺw���N-�Y��ߟ�%��ҫp�הprAiQk��<�b0����x���[�������ǟ��1�i�b"�<??��k��:�KhdFMNi Ep�x�_
�����q�>��
|�ɗ���chu+!CR֯>�z�u����wބ��յ���<K�k�����;�z������G(?�_��:�yԅ�o
�"юetSH%�W�}��1��?�S�؟J���U;�����U��@����az�Ӫ����D�Ȝ�F�Z� }^
+"��p �V:d�3�%%?(����7(i�V
Y3���X�.b�ǂ������XZ|B ��ڠ�0�cJi}��˰��]�p�������ڡ��966磛 *:�^i�
��7�[�|[	�_���>�'n����y�(l.=�}�.����p���%�?����au�1��w�՜��&�+!��=E�*��ڇ���Z^@g����Q��c�M�9�<�;�:q�:1���A�F�v���I	 ×���y�]z�J�o)�zvzn^����1�t�e% ߀��-%�*AUi�����<_y���کv�\��K��`S�K���ڼI�L�r$�O�9���X[�ߧO���'NS,����<��Q�MK��_�B�|�࿘r��,Y^Y��T(��1����e���Ȃ���r�n�]5s{Q~�">nݢ�4���Nkz%��ø��7���s}HJm��і��0�L�2ҟ�bb�2�Z��:s�����#Mxƨ���:�t���-�)�?wB1D�4��T�i�=|��|yUM�� I:&�ݣ�[SB��R�s��nM7�Сp��i�}���b&'�����J�p<�����������#GÈ{�$�߼?��?�k7��(m�5/)<�s���C� ��b�3Q���ƛ��4�{�nPV1d\�O���/����ý��J�P�H{D�����b��Sa4%ڲ��}����!h��s� qs�]4�ȑcp��>���e��җ������
����/W/=t���wo߂��W�p� �:qΝ\��an\��4��anv��GNM�3�]UBH�4H�AP�Q��a����}���'���y��@����t�l�A8�S/k�:q�YC!�����ݖ]�u�˕�[D�y�c���9�^�E��O(�a�8��l�������R���Lp
P=~��ށ׿�%��҅1�js�	J�z�f!���+���T㵶z�v8؄�/�R��M8t��z�2�:}��'��`iy����`��)�I/��c����ɜ�;mY�5h���i�~�0�oΜ���'O��hj�N�R�f$�p��E>�ޭsgi�-(a�%���1�m?m��UZ���g���T���L���f�j}�u�z�[Jx~E?���b8�ڀ����z�(�x@3;~�D�'�"��tcZ�ړ�aL��&{v�;LM� �h��=��2��#:�1�R����*/Q����D�a��>m���9\V��� 8;%3��B6Y����ֿ/oI���R�~l+^���Ι���P��]��y��oC�(���Oڂ��Z�G�OcJ@[#
♛=@ѫk
<�.>�3��(	EJSY�%�"���Ġ1��IcG�c#֑�3��Jc�*웛���U�Q�t1E���ۋ
x��~0:o��`=Z�^�g���6|q���<����������҂��%
�����33�����E�������20"���{����Ý�K����8"#ܐB�[�popjp���=N4B-���ل#G(F���ӊy탷��:���i�{�����u:R�W/������]<C������w�/>�
o�����K��ð��!�ꗟ��~	�^~^R?�_=�-�O~~D76�*Gp��q8|p.��W�|���-�7����/|x���nD�ut8Mj�ARި���(�Y.]���-��OWh��^�e���qE��G�]^9������O����CGQ�l)��ȱc�N���J�AU�̹���=�ץ Ğ9F=�1Eq�㣧+���Z�`im	f���܅W�#������C�qW�Q��O�7aqe֕py��c�{���ni��E�w�6�<��G[p���y�d�S}4���}�j.�����袋;B��S��i���S�@�;p�E���9lck�Lܛ��_<�;xBUQ��6�(VR��)8}aN���#�i%�. �%��s�����������g�z16Stuȏ��������S��c�E�zz=���L�['!��ڽ����2ɺ�W��[F(������Պ�͊�9)�:(�}W�K���bD�=ք/�e�)�jJD����a�s��+(2s��qAp���#�����\L1�]PJ�.��j3��ҍ&<s*Fh7c�>��\���p�+.��ǎ��|��p��G�?�)\��C���W�5�$��
�ĉ��z6n#YZ���,��Q�Қ�v�Q��k�p��8~�I���~F1��o�>sR�Elc�A{���	�)f5Kyܻ�~��ͯ��/?T����J���DB-�Y��j-����W��R��>8|(RZ�4:��4� 0��&��sp@I�=ф;����}�噖�?����t��l� ���ν�^���/���`��U8�4�#�N��shz_U�!��R�t��zG�zx��j�	"��R�s�z�m�Y�|�7�߅�� �?�4���+��Nŗ/_��g���w{�M��,�w��8t�<|��c��߿�NΝ;
���|M��qxU	���u%<����ޥaRd�x�S[��*���
znS��p��Ġpm}K�l�#K�^����':IQw���i���K�G����
S�=6Ke66zj�u	�������ǟ��.El'T�Z;3��W`�
�/�	q��3%P��?����|��~�)Y_��s��TF�방4q>x��h����?$�>�&M����E��#�=M4)-mL���L���Z{ ���;ܬ�Ч�o�$dc	7m��[P/�[�4p�a6:j�;�����0�ClJ
H�c`S����eR�#̥�n��t��\�3E�:���b:� *�f<��6�o+m<�ӫ�q��0g�A�.x첚����ۑ�:�xtP�{��0�wg4��@�xƖ$��%|��X"},����
���#Q�-Ŝ���j��$������z�UA'	�F�9z�G�=�ɏTd�G�u�~o�8SDlB�pD�������f%㗤,c���udR��:�2�y%����W����
䐙��.ߡEx��k������Y%�GJC����
ϖ�����8{�8������6�ʵgp�& E��i�G�\UZ�eJ��T@={� ,}Ii��&�W���\��'�)�V x��Ȯ����-x���
���`���µ���Ƶ�tZ��_ޅ~�,-������z�7$iCWo>P�>%d����pP�c�݃�kJ�;�����f�&���GK�	E&����8g;��1���>�I)o���<$��_\�
���Tm݄�w�~F��\�}Z��'�MS2M)�u��#%m���MM5()�����g�����s������1|��5X��$(��,��m��]���
\��*l)��~�bz<Z� &�Ҫ����|��@�3,�LZ���t�R�2�X;��թH 5W��Q~kNõ����\�w���O+A�uU�>1�ZD����')|~��>昩��=E 1Z2�$6���P��i�7h�>#���oTvm��6u6F����]}���j�q���c���$nA����@B�f>Y����O�0��z�L�O���$�Ӂ;5�]/:O	>؋�4]�*Zp�֚��̇�ʹ�W�I�l�%�A�۴�nv�	3�(�.Z����Љ�	|�M�?�=y��J~��u�Ѿ�������n���+�:מ��e��$A��5qo:�n^�A��a�̬�\Ugw�^�"�\f����#��8 �^&����}�!:�C��D��ߡ�r��#�H����r~ZAi�c�_:2��a��!�&�C�2L�)cz���a+�{��+O��/���_7�߃_*�\TR��^�^zn�Z! �:�O_���n�����U��q�����.Õ+x���_<�?����)�5�Oi�g�~gFT��{�6,�L�����J�<���Ӱ��Qx�t~��{�k_Q`|����O`~ׯ^�G����)�lue���G`y+���ו���=�P����,�'�[k�г'��_W��_[��M~ ��g���iª�ϯ݇ŕgp��)8u��.ܺun޼�S��=�������<\���\$�ϚǭBG��mC��<�f��p���G?y�?R��N!z��~��~���d�]��T���iy{�9Wn(�ل��eh+���o����	��l(m^1}�0�k阥޳���`�&�?ʾ/�&�AuQK�Z:}6���)�	��P�ԗ��*��>m��,O�`�@�8�%O�)`ё��IפmĞ�V۷��g�fr���OwF���vS$�%lE�쉘��-	d�A1��d��%��h��XN��4�����~���U��Ӫ}�G�*a��CJ�Acݱ���M��� S�x�[)9�����]�c�w���9�h��ѐRc�iORĽ�D'{�,��BH�����8���	Lȧ��n�F�
7�I~�M�Vs�9�eQ�]�� �`6��|���V��e&���0?��9��#������w	ʪd 5��ܡ�x�s@�K��-)��̥�Q��!R�4�]﯋�In2�[��~�&�4�H���&��n�#ŭ:�#-!5������7f�������=A�]|F���z
���|�����W��fu;)�a]���+�4����E�K��������	�]�lŰ~s������ 'Q�Y%��S�.�j?�|�����6|��g������_���!t^d�x�#����̅�m�5л>]��3ɬ����ω�Q�)cUDL��k��Mx��������;�m�)����(ٚ�z��O'���؅��w`��=��Ӂvs��{OSx���|~�+�5x��N��TǻO;�*��q�4nޣa�vz�.x���zH[�6{�eNi>SS�)�5�7� �&�,f�k�H���C��P � �nb2I:'^��&Q�1F32�03�i�T� ����� 瘜	��2�p���f�y���0�,ik�`¶���)�M�O2�;JFN+Ƶ�����	7G��h}�U��I'���w9�C,5&�Ȥ��:�`K ��3�q�=��ф��G�����p:X��&0��3��Hj;�@�T�e��[Ùu�P�o��X9�/�6-��g&�Y��-�(.�t�N��w(� �Ժ�]�VMy����SׇfC6�h"Ω����;�D%I��xr�`�\l�N�Ph��Z���y��k���y�b� 7���s�W?S��\�	^��F/��秭�%aΧ/��O*ӟȿH�����i�O�������o��i���θ 4M��bR�O�{k��aO���
iNF�C=�G����(M}� R��"�Z�z����Ӝ��\m��vG��	ˏV�iUL�惇2���)��4�v��E��ɲҊX^_�#�� ��L�ӕ�~W�F�a�jK}OVUje�m��z0%j#�w������܆ϯޅ��-�/�AO�|��24lD��5��nJfW=�ش��[�h�/	�y��5ub�L_E�}�?����nm0f1�� ��mv��Nn�0�_`�^s0F�71����o�w7Hw���G�z-��Z����w��ۙm�I�n5�)3fe��=��Lr�Y��?!]K%����y�,�}���DGڧ���K�	[Գk��s��"�9��۝��4fs2�u�ڈ���5t�w�~������n�i�B�N����t���]@r?
7���b��r�|PL�?�� ;h&P��I�7��^)'��Z�[����Jp���ҟ���e�/D!m���P<�9����9��u��Q0��r�=�7郀"s`��!��,�~Ӻa|L)���M8���-k ��T��e�CARŬAΘXS77�:a��r�Y��Sz���`� ���=��aR;�tzE� F2���C#C3Z���ܠ�J�J��bQ�?|/+m55��t&r��
���U؊ľj�|�����L�1��+Wn���!jL�֓:�Ǣ�Zv�6Y��?~�&复k���A�q���@�ڕ0L0rZ�0��#pʊ�Z��p,�ʤsAҁ��%/a�r�g�:H`mП�L�����V�P߁�Ǹ��P~���k=�����C=Մ�r~e���L��Q���Q��M�q_�V�!W���SF��� b�Ǥ�7O,X���c��O�@R����y����='�x`NI��-�?���K���=����O�k��͵N�##S� 6���k,ף���N���J���VoW%���H�xa+���\_ԣ*`n.��F��������v���8����!�s��j���g�K��e?�����.K>�W��_��f�KiS@
���<���4��v�fN�2L�
�dRc�Ʊ/B�_t�ms��VM��3 �����G��v�<��<���a��S�fט���9��d���P1�(�is�t̄L��P�}��G3a�������㎀�V���%��0eKH,#�H��z�X?4��c� Z��s�\f*��,��qfl����ب] >}G�I�y��Y}�T��:��c�4���#� 5���~rخ�:����"t�W��NS*��+'�x���	�,y�O�c�%���-;���B��Є�7�ƈR��9��<ᦍ>����5��wV����Ç)��uҬq2�s[v{�� �|����s��C�6��<^�Mg����V�T6�uZ[]*���h`kv��E$���͉x:�Pj�*%�d����6���ܻ�_қs�P����))P�l-��
c6��V`�J��f�355�܇^���t�C,����O����<�����بI�8�{m5a�А�BR���4�ў�liJe��:�e��&�5rpD�3:��Yf`#�هG]-�gzJ��J��Τ<e�%&H�cD�9�25e�q�����pܾK���	�`yJ�����8��l@P �z�{�����8G��Ї`Л��d�$M#2#!�3���?�}ԩ��7�kA@�"�-�:&}ߑ�rTӛH��1 `�8�B�[-<�)���/?
�ɵ���He�K+<f�gp����E���*s���h��i��>ܸ��d�\�s��"��SΘ蛍�.����f!̽`F/0ӱ���,�,ͳ����Nf��=��L5�L�ߙuQ�s;r副�;AB���%j�'�S�4`k���z�2�KN4$u���$=�6���:�i���Tc�	,��`c��؃9z��|��%���W�L#j�[��s@�K1i�En�jAm�2���c罌���u͒��I(0��5
�#��)`u�jf��m���Е�K�L�%���6�8B����Z]�LưZ(���p��L"�I�@�u����&�fR��
4�`P�1h4Y5��yǃQ0�&�Z�8M)e�(8�\)	���~��	}�J��-GS�O0:7`��0z� �lE"��d�o�8��=RoK�gzw�1�Z4�q��Yt-��K�Ǯ�"������D"f�"�cpS�j��5!8Ԃٛ��)��_�hȕ̭/�pp�i���<�}3��� �r�=�i�.#5�q�X�9�OSR�� L����9�r�v�, �KE���sݶ��n��7���|޾㈳�9$�s1m�6D�T#�>�D6�g;_����p����ݎ�,�O�K��YJ�r>����{:Ӏ�����FȔ&����|�9�n����<@�Wڦ+�;��W��xW׎�tNy��͌���ڂMu��o<�2}�H@6@��A#����>��Hϲ|��9���K�B(� e�c���i����̙4|�<�C���'V�O��=5�Cq�� I�����ln2Wc�FC:fI�i�#���G�.zb�7�ō�53�MO
�,b%��S龧�� I]�°^:�R=���&�W���������fb�sS�����
�	,�n%���V	��ݢm1�,k����9��M�m5R�~BO���3P�u]M����yR�8Wf�X��y `-�/N��ӻ�@)�� ޓH�0��2�l��tr��yු�p%qY����~������� �"2�X73�z��4U�&��"��{ᗵ�µl�yCn���3�K
f�+�6��X��m��ڼ{�����$N4Zқ&6A� <�7�r#"��(��|O��x�^�>X�����/a���<����[@[��:�
�SR؂h�Γ�� �h�����E��uG�	�f�
-X��E���{�A�n��Y`�@@��SQ_���v���#>#�ȕ���'U�t��y���$b��Fm-p+�5q�5����������dFMv�hMJ�>E{���0{����
�QCO#>�I�B�=�o�%�J�1�,8Rd�Ħ6Z4�Y��	ˑ�
�1��c�7}�
]mN^*������lopA}�t�hB�=i��$"i]�w�0��a�I��0J��ܑ=#` ��uTl�3w`��Ci���N���2�XG��ݼ5�j~349�?E�낦�I>�'[��	O,����ǀ�)Y��i!�e��9�ԕ�r�t�dC�0�0�[��G�s�>,�����,V��]�-�T?�a�}î	, ��7���x���O�s�E!����$5q ��0(M\p����7������ɝS��¬��w�Fx�r�<�-?A�<7��[�$���EF[F��M�g ��^j�  G�S�K�u�8�W�}�$@�:0*N�<e��zsc\z�����	�zJ�ȋ^���kSL󟌳���,����oR8�>��*��������x"��L˘li�6&�K+�[I�Qka�����ڤM��|G�(����xc�}�lV$a�@�ۖ���0�>V��vI����5 �S/�w�X�c�[.-��@���L��Gj	}3�~E�l��Թ���xt6��I��1��d���5���B��|"?��E�p�v��J�޿~5�?o�0�G�sF�#�/�5Kv��H׾|u6����(�T�l��{�ۖ|Ԅ���^��6�ٞ�m��$���8|��n�̌�t�ׇ�=f/����fMd��0��z��u!��1����MM|���&��P�u_�4�73����"1B ��'r>��[w��"�F�~�ꖹ�Y9\ۆ����+?5�т� �� @���E���"����Vd����Y�J�3,h}�$>p�v���om�f�3�g��>�֋��k��^�q� ���z�^�Ь�QW�/=}H�7�i?�W�L���,���������r:���dd����A5�'������u����%�����_�fX�� �%*�Q�=�-a�-G�1Fd����7M'P�!�F��t�U����(�eO�	е�E�h��Yg&ʪ�;F(��/�4Z�YS��d���(T������+=�p�5��m�Č��3{����*;��K�#�$h���ǹg��,��:��F�k��������F���Pk�:3y�>����h�^d������,���^�,5��Q٦ҌfIc��A� ��23�MW�
k���ECގg��6ʏoLM�ܟ���wۙ9 ��m�ֵI���r�D�&���On�� x�=!ƈ+�M���]��������������L���D��:�7?v�{K����{΂���u7m�0�C�� �y��<I�pF���b��{}�ɧ��^u�Zj��H�������Ȅ�bA{[��6Ū�P%d�gd�`Ѓ���[��;o�@?��i�y@gSfF{J�4ۨom�F��C���*!2�/�j���2�"�Y�MW�(�q��*�Pf&t0Ro���n������7Tkx)8=F��1r�rQ#��%!��^I���������X.�?�c����tt�9{�$�IajJ��(q_1P���`FS'����m������B�S�?�ef�m��.��DU�F$#��mg�<����(`��L;�_ھ�';��v�p)e�©��r'l�I�mV�{���;$?�;���AYli{Ud��]����r?	=�00�0S�;2ϱ*7ٽ�U*��7��Z�B[k�^n���������� s��Y���7��f�Ǎ��y�ƻHxٻ�Gh(7a����9=Rd�u#&Ji�v?YK�M�-ݣ�-�DU��1�0+��E�%�b�qܓ�ô� ��� ��d���^��0#A��΃8��x��@�$(���[|ᢗh��/�r$n,�6/#���0�ީ�p�V�a�`z��
Ơ��m��xر��#������0[��h�Z�Hs����hL�����Q�	\��!˲��Q��G�-Q�z�k�(��jR���N{s�+9 �FSphP��;!��*3n�k�m��m���Yܯ�����%�������y�L�%x�e����w�M��"�Se;e>W��"�k��n�KYd�w��v��� Á��'0g����&?��J&L���Q��M���p-�;@d��Fe,��t��άtJ �sȿ�k�7G��Td�5i�
<:z��ԷZ@�]t��m���`d/�?�{�O_�k�c'x[)�$�\���;�t'����V�n|�{v��B�׃�]7x�����9vQ�\�&����j�t�!;"�M^�8ɏk袦h���ބ��an-:����h��L�8i�~dd�x��L�(2�T3��4m�۾��"Ҝ3m���6�Ϛ�����7�5J�vb�j�y����V�F6�پ�@[�Z��M"f�&!�� s�vf�����5(F���j�3��I��� 2�I J�X�ܠt�B�O�K76���2/��옝+��x;g�c][`:3�~/�/l΍5����a�-�K~�Z=03@�,M4'}2�E��7/L��*-���a։�ǉjaB3N!}+���Ù>ȿ��<��?ɾ��f_C�e �����͞��素�kϋ�l_c�w��������[�0-��+H�ױn��|�|'�~�,#0���0���&�b��ذ�"�W2k�����.q���y��V���"�n|�-�0���,��gN�`��&����H�����k�h�h�f���o�f/Ǒ���/�0��Z�Tń��NJ�W3�#�)�����mA�#O�V	���������2&���3cno5�ϕ�Wa�}�mOc�g�YM�]pZB_�-г`��Mۮ�^/۵���}^Ƚ1E��,pa��ܸ
_�s��~��W��;�iO�G+�s�dBc[����E�����s7+V9a��������S�}�F��	w����>#�	F��� XBk�@Jw_��p/Xw�k�K�<Kdn��3|�;�M�
d:���Jã<y��-J9T-0w���~��ޡ�jQ��9�
H����"t�w�h?���j6{qc�����(r?�fwf�K0/�Lq�&�Cd婚cD�!�����@X�����;�v�{����M�~M��K�T^����q#�ܠmI����(}��d�D�O�>O@#)̩��	ύ*;+F�гF]�:s�^2?���F���G�Ϭ����~ɸ����*�y�C��X�qh
4�
���,`���r%BW�3���=ͷ��c�|P5�U	�(̏����־�ĉH��r���� }jj�7[���N����L���:Td�/�a���PB�{��ZE���!�` �s��������Ή���G��0�^�?��P����S���a�vu��ʹ�߁�U��4���
G�[0���2)����n3�9@o�Z�F���#�/)�Ѡ�WZ��$��yF��Ҹ��|�He�qӨÈ��_7bt' �K�TtO��2~߇��[�l��:�^��QiP�$�2�˴�q<s��;A�jc�y?)*�_��z�J�ɱ9?��l6�G�קf��J6n\Q.�\gK�g��x����Va�b�e�T1�V!��"��_� m���ޗ��w�
�C�'�a�~��r���4��v�~�0�w�q�3A��
��4��^v߰ϫӮ�Lu��.����(���
��vOP�C�7'�f�ヵ� ��h��(d��DR������U�6������<�u��<����>�Q�ې�<��43���V���L���gh|������:�h�uP�=&!3�UM�Ee|�Z��.MR�����q�/��´_�s��ߗi�*��1"f�����a��8�~8K]�(��2� ���y�O�I�"�g[Uj3�$�z��qi$!�_�u�t�̨�ײ1*z�Q�rT���<*�s��S�mU޷�%cT�N�0s�n������t[�}���2���4�9@ǃ~��_�>��)h�A�K_���'�U���]�t;)a$�\$_H
�q̤�}e�e�t��q�0L�h��YE[�$WP�lU�ȸ�TK�0l�¤�k\B�v��A�%���2� �q�Nc�%���H��z Rk6)s��\�A�c��ÿw��1��e�����f��?>,�n������;
�bbh�1/kK����I��'U�� C  �?+�:''a��4��R4��� ��r��<.��kϷ�է��/��q��V�LҶ\�m%��=G����Z��31�2�׹�ׅ��x�he�2�ݤ9�EM.�*��������Z�m��o	z�!W���sD��
����;O{�ч�WT� }d$�_�j�і��ipU��a��Ef|�s�w��4�4_3.�g��S�QVf����@s�ZX����SU��TVϸ ���՜�S�^����!~9�Q�j��B�z����̇��� c�'� �)ί�!Q����>�qx�3��ݵr�[�\�l�$-���0�2!!꾟޿?�}�6�4(�Z�=�fN��CʏY~<���Tl�̲U�:?B������E���*tE��sC������Hج+Ljg�κf�е�4�W�?E&�a]���*֬��%�l�ڿ�A����Vҹ� �42��v{+��=�Q���~�����
J����y��n�8�ƨUq!�5����ƥ�Wmk�����e��ҤL�E�4���e��.�i
	�e�9k�-b3�5пJx�����2C��NCg��i����G�lRG�1�ֶ�)?S��a��u�L{Ta���6���U����q�0&�B~�0?��AB	~S�	�fyЦy���z:�O���t+��=	�B�n�m5���	֗F� ���"�n�qP�7�F�ݴ�@��F^����Sc7,@2َ��\ uh��j��9�	�יv�&_6�_��n�Ї����LSх�=�q��P���An��n��H���$�?�:���y��5��f�S�s�>�u��:֑��f'��ؖ��j?��2a@��x��̎3�=�Hz��������1N�qL�:u�������n�q.�_G0�+T��A��!��(T��w[�Iޕ�ߍ
�øH�2U��l�:�뜷!���C�_�����/�g��8[[�;>�{БYC	u���o��]��� Be�[Ҿ�� �0Z�N�8�*�84_B�-�΢變[��Ӻ�BE�>�-�tC�������,��>tه6zܢ�Α� �7��M����$��>�1�a��q�O���hҚ��2��#u-�նq�y=�mȕ����h&A��w��ݶ���\_��֒C?�;o�}��%B��3�G�}�>��K[�z-�A@R�l^�Y������-�a-/�4�A��k�EEf�a�Tn'#ɋ���g�?\~��ݤ��vC�9^<T���3���׍����R��voa���(��$M���N��{U4�`;*J��ZE|��Q�{�zU6S^H6`ͯw?�w����LQ�u�q���;v��w�}�^To�����㠺�nݹZ���!������u��W�I�v����zm���������A��&�_w��B�8�Ȳ�Q��_�π�L�
�Ӧa�_E �BU4��3�q�M"�����f���q���:��v��&���R�)QE�V���kS�����"��|<��$�'�~g#���]����;̤�-Ҡ�լv;�z����!ԟ��8�Cv尾�: ʔ�P�״f�h`.������d���ܣy���!�{a.I`�{�t�ߦl]�s��=d��0���w�
��.�~X�����Ί�y�*�����r��}�_���;"R/&�N���۷�9�ץ�fQ�$����A�y�T��X&M;&.Wf��2�l,�M9���	iS,P��Ph�P�5O��$kO��(lO(�rW�$}���W'ƠP��Oi-f(�l�B)2�Cze����T鮪Zb��o
���(�'�j�_�2���Gd�ξK����2�5#̷��U�d]d����2�%n]K0�!�N®[�Htq3��Z����߮k�Q�PH� &����j�Ks�t/�����Xd1ʬ������7~�=��4�fҦ_�5HERi��9(]��{�d.���4�v���T� �c��a�~fJ�E�n�����-���Z����<���%չ��\]�7��`R�
�ƥ�5�K�eY}����>�|*i�(XI��u�zh�L��T�3Ӳ�jV2�LN!� �|�jg�8to����}��;���jK1U�����%�����9�Ϸ,��
�]�s��+���^�����7'�Ba���K�eí>a2��K�Ϳ�d�"�l�2�L}7�ch4��T�L�K�(eW��I{��{���k�u��Ts��=a�'�`����i��lw�N��'�����T�ꛅC�:���}�"0/���|�e}��q"�17�y�(}2��*vAxP7���ga�n�k�����.��q�=��:;M�|�s���h�֣0&J���HF�f�K���������0�"6��Z0���n5�<�3��_gX_�(�T�I2��f�e�&|�3����#lR�C�,����y����Iu|�LE.�*���v�E�����"�:.�� S�Ten8���̽!�s��N��(o�*(I��
�@��m�Y��fm����K,\o��s��bt�H�M^�c���"�Nh���8���@A_��+X&��!gr_�JE�_�X�;�[0�Au5�|��犞.p��8�+�Q-.��;��>�rX�ya+N�*�z��Z֦��_U�C�/A�:�+%�sə���	�T����
P�s����'2iPt�!��vfj���G��3�2����	V�1�Q��n�A�g��r>򰉏�j�:�}�>��_u^Ui[�`X��G�8��W�:��EV�qY�K��Cy��l��V��u�"~X���o������eB[���;�mֺB��>�"��û���9@��zQ�Kc��)ՒA ����ɭ��q�$��F�"�6���3����*Ϡ��}?�F�a��s�g]��5�*�7ȴ����r^�e��g�u����޲�W�J��m�"�|vϷQ�h�O}������s@��Ӥ��v�|A�_��O���$�E;��<�-8�U��ab����4h5Pd�yuP{��S�юڞ|�a�G]���~cՠ^~����*.��s��W�̰�]vO^8��g�0�$^֖a�2Kj�2�gq��~ Q����J�%E�~'�KG�S�� ��Mcա����5�?�2���n�~��X��8��S]�A]-h�}[�	�մ�����Q�o�i4�L�Z��3NK����S�z<YmPF��u0�޲����iR.:�[��4�:�[&d���(�����.ؚ��t��]�����)I�H�4e�D�q�A�}������yD��a��~�>�K�ۆI���B����4ȴ8�矿�:�Z��NS��W�sR�^�*���+0X��9�^Ud�
ġ6��WU#���e���Q��ٚ����Ҁ����D:yi��9@W���y��Ր�L	 �u��^�C=lB��d�]̫�����M��	\�g�E��е�Z��5]Eu�}��7�֨}��6�QY[�9����7����	�ܨ��h[�=U��u��J�5/yW]*�:��f�>��cݜqԬ�HD	�� ��0$��>����JY�p���p����lT���R���Ii{E>�"��f����E��O>ujY[��\U4�2fWfRnnLX�5���i�z}����>,��������ذ�x��\��5�:�ɁujCiۡ�B�B&��m,Gw-�O�����}Jk�D�c��d��$�s���ұ+���Y��`r�N�C���� �*����>(X��Q����QtXX)4)���,��jg�SB]a�(�Ơ�ŧX��"l�-2;�K�)��H� ��.�:���U�jQ23�̚+�*g�dL�Ṛ��ܫ*t��O�L��5��y�?emvUaD��zC�n�);;�5$0���3�(!��z�ש|�Q�1��3BRk�eJ�v��4��i���*�+ }���H0�k�S��s�q�1_�Ϭ��|�Z��y��3�Q�Y���L���T�j�SW�.Wk���R&tԢ�_k<cZ��e���:�1�O�ƹz�@��S��4��S�j��H��X���X �Kyy�Pq^�'�9@W��ĨBNl�K���Zǚ��C�sG��EU��hw�9�(����5ǲ��|���!͸T�Gնv�nw#�wyM�
����2�2�sb�	"ô����>kR��u\������hx�M�Qc�mP��P��b�~�s�Nz*%��d6��Qz<o>suNvټή�|;����#|1�U�i�����+�0m�W�P�Rʨ��_Tg�3F���z�8�� wI�&��^�:��"a4TnT�b5-s����xn��]�0����G�Sh6��՚���Ud�����ݡ��9@G�(������w��,�S�,��{��ښ83OF�8˾�B��I0`�l�[5�2�B^��M4��*� 	��nKѼ�6g���.k�A��;g��J��ʘ���r}d*��Q.{����� ��S֘���)�]�v���%v�\�-��d�'�.7Ȅ[F������:~?A��hq��P�EU���j3�g@K��"��������R#Ԇaߡ��AV�a]U�8��wP[�g�*܄�iPc$�J�F�5�UH��o�γ*�-�=�O]��r�fw4�'��d6�;BF��mw�ʞt�D�A��f���&;q�R�I;ٲAx?�{X�0�Ih$y�]�1�?�j�v�0:S6�egנ���s����:}7�\f�� h����s|p���<p	�9�U�=��;:u����Y���5�[� "��?9]�j6!��$�RG1ސ����2C��X�5 ^�\9p��
�i5?�N��ڠS�C��`>*�i�/��r�:��^�v�� Ԇ�@��yȊRIS�a�8nO��a���N��|�T$Dq��uA[�t�2ԾY����"��%I�"��pY�v�9@W�*�I��f���C8�|>k����$)/��'o�4��h'����q���/���~T���A�T��{�is/� ���z]��8����X�*>{m-��}�Lѽ��	��I=�)I��[��R�K"��e�K:oO����ϒR�v�Y�����x���O���!�l!)4�c���.cZ��V�eӿ�[h�q��b�VY����-�V�_�y�T�S.r��+���������_6__�uTԖ{�u�������c��*JZ3� 9�CB3;����6wO��]�X����K����_����h�D���`�i�l���g$�l�~�d�|�n�z��:�\��v�B~�<�M����;�؊����2[ge������]��b���,����5F���ې��A�v�]ːM��	�,��햔2�����]��� �g:a��'��2�!<� �@=OE�~��c��n��Ҝ�X���E 7�y@5}��&E����%�<i�����f���'^$\������!��Ny�2K��|����� \dNϗ�9!-�����U!�^�����"p��O�I^����'��8��e��nG��Ȼ�)l�)@�65��3���2z1��73�߂�@{��(�:Z�A�{��&}ƿ��F{ 1fyo~��^Y�0&�����^�8���1�A~T0�~�Sa��r�3����o�A���|�,%�U4ETط��l���2JR���+��1��;3D�/s-�=\?��#|ү��<�Y�c`ކ�^�ټs�Sf�oշB�������!���(�y� $��;@ʐ0Ȃ������+M� ����4�7�4�~Tjm��c���������������e!�����>�bn��컢F?#O�m�=�Mt)}V�o��e �j)un�&Z��{T3[�r��4�d��ba`�
4��TU�_+k3k�z6��7I53�NH�L����s�@���55��E�U�m��0�L�6�_��Jx}��Z�����+^/��?!7J�j��̖f�l�����~�����@�:I��5\v����t"D���L��u's����D���X�H �Lf{�2�'�8�����]�%h�h�~�b�3%��>�e��s}P�Af�zC���\^Vv7Q~��������/WV�OEV�0ױ�L��xYyV��w��ޚӧw:�'PG��GB6(�}w�\�s�>;���������d�p?��i��*f���Z�n�*�1�a�kX��0uW�"�b�����G����[��%�:4H��2uL�e��"S�_����ٿH��b	�Ae�S�>�6���Ipo�Ⱥ���Zyt��Z�Ԅ���@{Ч���.��c}�}Jy�g��}'iPȗ����qZ&Ie�Zյ1�6�i Y��!���.���̟u�1n�D��Ѫ�:m�EZ�ߖ�m��N3��_���=
�W��)�
�}<P�����韻����Z3=5 ��D�<P�	S�D^K�Xey�EQU��{=�{�+���ȼ<H�F��3檦�A@5,嵯���]�Y%�����]�۩M�[ֆ2-=O�����2z�g�e�G�Eu�S�:H/��]�4
4V×�:���v�9@�$�smK���(�I��r`��L�Q�-Қ&���$S��<S���ޝp#�բ�7C�}M	���*f�� �q��0��8˅��nH�6������0�V�y�+!��n7��̢�>Y��5�����������OEq"awh;{Н<D�-]2 ;X�� /�{Ʉ,� &m"ԋ��cU�����JUe�uM�em�}y��8�~��TG���yϝ�B4>!��Q���q�{�}U@�껄�Yǲ���_���о�M�����:�����B�8m�qoz����M@�sk���0p_f��z�h𰔬���L� �HzDU��U4�I�(�X���ms�Y���Uח�?3�0�����0Uyv�9Z�Ν2���e}Qw���2�ץ"wа<�o�8��]y�&T�~Ι�#s�g&�B��i�Q,�8n&��;���M@O�:�[�����?u|j����}�|���h��ݢŌBu�hR��Csh��=?����&º}R(�P]0�n�&��a��熯��܋�Z̫�o�"��_��E��p�<�N�*�(~`�u�ޠRɨ�����2CQ�ې��ODJ��1%��h4���&C��p��
f��Ap��.��M� Z.Tm7h�z�=e��kOEL;�$G�*��*m���y7q�n_��4���]h�_V�	EV._C��y����qP�y�k���o�	Ѷc�Ƴ��{�w�]���	�9@���p����)��`���|�f�����ɝ�����.�:�h72�ܓj\1^,s�<�0�"�λ� ��[��u����#@�Qf_Է~��=I*R���q�K���:�_����z�\�b
��(���!$d !.�	�A�.6����`�q5���O��݁{�U�!L'D�B���c��)��w	f\w�I�~�k�s{�ꂨro3}�y.c���%���T�,C	�>jTn�L~q����{y�+���Z��Cc��$T.db�3X_c*�>����Ec�nѻ���:@_U(�R��G!�
����.U�U�_������k���U5�AV�P�g���yz���
���ɟ��R��|��P�e� 2�qD��t{b�~.2��$�=^U}����8�w���!=�Q	6�-7��́,�{ewYMJ���UV��fUT�-"ը�pT(U�U�n������_.O㲆����+>�!V"�Рw�2�ARE}��'r¼��\+�^U���Uu�Ck��|.��гBBF���	���������w�@,���`�nA�=	�������Sf����0��J!�.DÂ�v�(��8������K3c0i�L>�b�eZOU��\~T������+mМP�S�^D��Yw��s݄�z�PtO~.��Ny�<Ԧ|?��ߍ3�;�0�\F�ϩ��:�RM�$MvCݓ�ɨ��B��4�1�K�0�Ikwys��]��^��a��(�L��R����qh��4�a��ElM����.���՚��W��Eu�A2�6i�������%!�yQ�E`>�-��;Zx��)����{ >���&��	�BTFf2�j*p=��c;Lr�Q�n��� 3f��W�?E��vS�9��a��a�q�g]��8i\�����l������}�"Ծq
�!0�+�QY!lrQ,��Ω���	~f�r�i�{�)\dl�:��'�~w�iEöq�Z�0T�؊���*�^DELm�P1�}E��˰	��p2���9׹7dN���<�k]���ahXM����iCQVq%��Qe�W�2��|!���n/5ep+�L�ۧS�\C����C�¤�+�`Xۍ4	FRX������m�����/b?�=_�N�/��|�U5��{V^*��W1���a x�T�Y������a��q[�����;��LU�J�g�L�EZ{�ސ&�տ?ߞ|���C����G�G/#�7G�(��M��'��3��Q(Ȳ���D�eT�b:Vj�l���`��ᄘ���?��i�!���jsU��0�]��I "R�v:	+ŤA=_f�m�瘟���y�p����3��3?�e��>�!�V�����T�y$�'�o[��A g�x�ֽ;a�>.p�I���a�Ѥ5���yѺ��M�ETĕ������Ft�fQ�e4nA��0\��W�&�.B�F�k�
QUP�j}��a��o��"<ˣ�m���>#���4��ߪ��Q����L���#��&/�NӞ���)J�ʟ�D�>	p&�2\O]`7���2��B�D�&Qg�&5�C��/v��7H@���u�V���L��8�l� �A�9h��	���ߦ�]V�2*3W�A�=�Z^ȃyC��" ���u ��oY9�[��_���~.x�P<CDd�U�$���蹆>	�:��!����M�l�8 �{�Bf*�<�m��2n�i��^�_�c~F��27�)����.��g��R�{'e./�:F����q�$�d�m���JL��Ȳ������:Tfj�\P���ɧ�e��N�t�b\��8ii�z���>O��붝�IF�E��n��IȮ�{�B�:�.������`܂G@�}F�C��	i�e��>��b��3�	��N�V� ��|@���s� ���0��gV��̛�Y-�ק��jWY;��7��:s���}� �q-{-;�8i�y���2�ޮ �=�H$��Ŝ�h��1�/�vצ�4Ml�\���ƁrB�Ad3������Ȓ�eVu��{o��%��D�(�̣ >0?�|�I.?�`�A��D��� -[�lB�E�2�����twU:#3�**:"3��g���bw^wWeF���_DdV���)<�X�S�vk&
|n��BZ�=ZW*�f��Uf�!��~J�P3VZ�O���B�}���~�W�M5
��O��}s��s��/������y�R�s�.����&�dԝ�3zT��F�u�����ڋ瞃���[ӶQ9�����\��p�I��P�i�8��j��w̟�x�����Lt�����_���(P�@�g�O����{ï���E:�C9��%��ڈ{#��
XR\%^��=i�����v��q��T�G5eK�K�k�s#Q�gɧ�p�W1�?~�Ҝ1��GkP^�bF��u���7gDI�N��Ds�j����!]j�m�H��F���^�k�����;�$8�5�=E��b��"ԣ�i�T���$�v�}�k�_=u�ReJ���~���y���/)ϼ�ΗY�h�F��4���Ws��Ƅ�G��-\>$�W6\�ĳ.�� x��8P#���`��H��j�k�]>�h��z�ېg����ƈ�i�5�Ŵ�<���!��&]s}Τ�I�S�ܪs?�!��#��n���CSP����:��%�O����kW5���a���r�9i���+kx�%-*P��ڱ�D=Kr{.匐��?>�50u��3_ɠ�zs�O���/�@�05}j�}5�JzR3�9_��iÈ��-��h$����3�ߙk���/^���5��i8e2(\Tlr�+ˎ^��Д�% �9�=�K�{��{�O����TB�<�%唗!U%E*�ɕ����9�Z�l��_/�S~O�����S �޵�LǽN�t�<N�o�Z�j����`:�,x���_B���\�^�"�����;��m�M,�!o��ѵ�8x�b����^��.I�^%o���y��$��҆�صu*E�FS����5͓ZR���r��c�#ߥz�!i<EO�M��cH�I�i�rBZ�T�P�;��t��ZM����3]n`e�#�د�t��ǆ�����\��qs�޶��h���n�gP���1&�Z�5]
aI�!��yD%�X+������
�~ǵ9�$/��QsT�%mj�p-��o_� *�*��EJ�k�s�9�S��Z��������2��S0� �0Ԏi���������v��:��=�Bu5�L|N�%0�%�M��7����m�I��ts��^4�N�l�A7XQ��0fr:\}�I����-�=��;��x�p���yk�7����>��-	pr�N�Ε��!���d�g.P�zԵ�\��V�s�d`����Y*/>�xz�ar�򈌄2�$�ԇ(���5�6'z�yP����Q��1�(A!��/�������\�.��\0��N9�Ǜ�RP\�ׅ�t)`�>�H��e�]�|j0��sϔ*9-�=�9���/.�ݫ�/)���x���o�����)���R8#B�!��8o�{�k��E�Z��f�r6��wjs�u.>&��8�x7�J�X�ɜ��CT,C�����ִױ��� �ի����z�:�Н'tI�O���T6,�yP�E��Hs��T���*���Ռ	�%`��R{K�_�&ގ^5�AM95m/E�2��˒ʛ��p�e E�� Vm:nx�N�P�Ƒ�m�m.���3�O�P���7���#zvl|�D��K��}��5�����9@G�'�:S!�t�|K��d���4�( v�[�8.1ٟCa,���Ҕ蚜.� -���8� g��W��uk��Fm�z�9޹~�����jǭ���a8����C!AO���pӁ����>=�ؚ�^�v�L̰�M�(<~:���v<җљ�������H�'Ϧ�AD�yq��.�z�p�sK(�!Ki%�D���%h��)��]�w�˦�#)�R�WuI���\*WK{��/�YqX�F+_�;s���c�y��!5yF�f���0FM�(�'����c[���=t��9�I�*���|��3=��G�Bz;>[����u��Bz�z�w]0����A��������+V��]�@ы��ӹ�Q��+�(�	��r��K^]m}j	��?pE+�F��]������k��A�/y4�N�P��&DIyi�y�s���i�y�!�=Ӿ������s�Bj��ʹT�q��B�d$gXict�Oj�4���;�~�7�Mǋ�����r�}IR�{��n؏E�`��-�+b��l� �����ڭ��9@�����X�w 8�����i�=�Ѻ4)�_N�\�4�"�c�p�(�\�.Y�sQ(� g.�tO��jy]����.cN;%��������7���H���������F�\D�Me�2��W*�G��S�}�q�W3*���S�E|l��81����{w&��+��Ǐ���~s�t�,]�A"����z�7~ ��A��<�	�/��d�xs�J �f�ϭK�����-)��Tޗ�%�v)��~_C������\�[J5s��-	��}���Z"��O�Y�g�k�<��!M�&�K�S��\���S�=W��q68Ɩ�uJb0Za����ze��n����7�==~�3lV01��lz��Z���IV��X�Zk��J�J�@%/?�jm)�[�t���|$p/Q-(��y)�ƨ��sxs �K�Q0W	j�59�
S��47<�T�8o���F5��y�y����6.5Q�漟�N�]Z�<m�����Iu���8��1�",)^����������4�ѝZ�@��Cj}x/:�z` ����?�����5˼F@��\�R٥IP
����"�t�BR���9u�c��xH�/	|OE��k��t���^�f``yH|]�f'^������59�c$jTk�O����'݌��02x�9��O#���siV?7�o�ֽ��V'ts�n�g�#���cc_F+2	��ۇ�{�p-m��4�B��˽�iY�>�k��|�K�K�D5^�%��y<%��֥��K��S����?��>����[�Ħ�i	�J�p���R���Q)Kk�'��6jYklA�1Z�,bT2�ji��L�v���i�qh�ֵ��
H�9@x�[w<>�jK	a�~���M��ސr)a>J5�v)�Jyj���6��yrП�]J���J�=gx����G󂴐�9�$L^��=���d)�47r!�!Q��M����-zR}KsWk��Fc�=��NLK�&�H�cL�����3xj��%q���)�s�W	�8�2�+y
�����޻����tX��O$<� ό��x���M��RvK �Vh�I
����x[�	�E%��P��p�e�K�A2R�w� �C�����[+W���K�vʋ��r]�Z0y-�pFx���<�k���%�p�s@ �����A��^�l��ƵW��n�?��Sg�.��&u0>B0	�8rjNc�������-G����sej�.�J��$)�\�FZ����)���tC�ZX*+����k��ғ�l��ij�R�t�RM8��چ��d�d�#��Ba��W���|�,��N�|k�xb���p�ݩ�~���i�֬˜G�O	����� ���bg�:�Ե���r�t�.��9��6��X4�0�N��ܤ�y�xMR��F;���>OI%9���)��xIO^S�K��9���5��=q-=Rig{���q?��j���9������9�ߤY�n��P>:�����9l֓��۷���<t��O��0��6=�1�s� ����C������u���*���J�=7$����O�_�j���<%*�sy�5c��;����g˽�%4כ�s��o��6l��C��O��ZJ����KZw�}	���Yp�k�M#4���1�.:o�M$��=�4�����	k�@vܜ0N<����ѐ��:�}2��\.A�`���d�"�yY�DZ��u�}Hu�$�g�/�CKC��ÉP�kxK�'�Wch��\O_t�ɣR�>�.x��5�5���NH���q�q�ȱ\�7�����i��!oL��0c1�N�񜴯C��̀�߶m������\�찆BB����M6zh�P�p�N����MpzMJ�m� ����&��+��@JT��wz��$k����\o{)���*,ɞ�'�Pv��J2/��ş�x�H��G*�m�1 1@R�i��C��G����R���Ѩ��V�{�����O�~V�O֌ag7 ��ﴏGߪ�x��,H������p����Щ����Kg��Q�\�iz��mm9A�)L�A������2���1+]T���yNQ=-qJO]�s�F�פ{*Ң*��������A��(��%���ӢQ%:'}�xʕA��D0��S3�j�ԉ88Ux��>�P�'��C�o4�d���O�1FC/��V�����U(�p��G���`��q�f�S��<C�����Q9-Qr9@����9��n���s��%��\�6l]J�M��n.ե���{��<�R�Y�@�D���m�@^���v-1 �QG�z� ���_҇��5Mo��o�mgs�$��|�w6��tC��.A��4%W��y�%�)����R{o�j�����Hk��,1�楷}�ꠥ�k��5|r�4�)�@3�)�i���ճ��Rt�9[��ڈax¿&2)E=��iRvhi��n�_�ze�nۂju�x�g����+]<���CbOFd~�h���!���^z��<�s&�owIyK=��T[�9�_
G�5S-,��.��ܳ��h��Ϲ^�k@���֝�����a�w�q�\��e��g���Euh=r����Ӳ�ޚ�csts����Is�ۑ�3�9���Q	F�j����Y�<]��r��熉����:WM�.a��:�Q�������R^2 �q��sǀ�l5�Z(3'kR�R�ι��G?y=����p�C�;j���$+�FUd��*9υ�y���1��ֵ��/�|m t�;7�d�Hvx�Ф=�ud��T�KM�s�Z#m�H�@U��F�Th�ٶ�z�u<��4s���Ds�f<�4��]�R�dh�r���ZoZ�++��#&�������lM}j#������yʯ&"����N�8�o�W�o����<��m�6z�聓g�7mn���#dI.��P,��k��R�Ry9�/�s��T�H�����ں��\1����� ��5/n���^7�k�l6�Ǩreֆ��p �-R%��e	̵���̉�p��a�.��4R,�ϣ�^;Y�%T�I�|ts�~<>��N�$��JO����7�t�.�s'o��SL�R�K�����_��PM����`EA�S�̅fk�0ר��Q��C�*K�0�V��@ �Vn�j���,���բ5u��5g��>y.P/�Rg�8�3J�ʢ�I�#����_3�@7�@�|C
��:C�tM�O&��z\J��L�Ð&qM��k^=�bnx��=�c��2�9�j�y�����ߩ,I��F�r�n�Sڹ2Y3�|�Hu��]j��^�sdl��7�.�"��W���P����~g~g��nЏ÷�J>�m�f�J���XV��1_�Ä҄ȅt�b[��s����x4��9!j-�S)�K�3.�w$k�^<��ja�9�d,r� �\?jz.w�G��y��:���^��ʏ�'?N���,H."���ě��d�Z�&l(�z�lY�܇�����}V�I@�Jc�&]��脉����g�0�z��)�-� �橗�q�
��O�S�R�$G�=׬�$�,g�Q%�o�^aNNJ����k�� D�Kis�6�@��h����%�F����9`��k<�9QN5:�ϳ���5������[�x;���@=�����N��]���wݡi�v�i7�ϙ�n�Ӻ���O2�߼��0V���&����!]|��F��*����O����am�[�	��ʗ�J��4x<ZvM��
ae��(ޟ�M j���ZE(�Cn,�{Z�5H:Ӟ��|%�'4�n�׈�����'�:keq��-�����"�W����G�ס��O��<v�>������6���9���t�7�[)/�[N�����^�o��0�]ļt�	��7�ry��.`9���m�W�#sts����ƣyۻ�"�t�~�dg�:�!���ƹ0Ɛc�����u�R��d���IS~K���$�))C���f�䌇%u��W�(��x5|�t��G2KyKުԎ%ޘ�[��{syS��gL�Ɉě�G^�WJSۦc��%�T�!/��s<������9ϫ��V&�!���!�/<dL�g�]�3#����h��6a��^�i������E��n-�m���J��D�	:z�44�u��(���r��x9��Q��_K+���C+Sj��F��m�<�Z��9c)�N�`a�;�sZ�1���s���#��y9 ��-���4����ʝ�?������+��y4x��tM\6���Ŝ~׌8Z�p漤��Z��s�T�%��M�r��`�@K��S3De�r%����#/ijB����]s4�;sts��u�����6�!=�n��9vGx�?v��B�.�w�'��8�d��^\LC��w�%����t�>�T��ESZ��T/:I�>X�	Onh9M<�`�s�v���-JZ�rF��ٗ(�g���z]��Mɘ��B�x��3W�����#{Z=h~>�9��,�z��f��\�1}�ĒP��+շ$�������p8��4� �y��;����j ��-(p��R��~�O�9@���{���-7���<��K��x����e�51�j�K�C8u�m��TR@��]�e�Mt>�j�Y��e�~�<�C��9 �=��һ��xR[j=�R�����kN=�R��+y�%~�2)Ѳ��2����~��̓�ɧ����P�K���h��Ơ(�0ר4��K�Յ���&>p�� �ml�3�����X0z��us��vwױ��� ��a]�tk���q�{��o���ϓ�$
JD7$Єl����R!����K�-mZ~��,�T�M���t�̹��e-P��_K^��H���iu��I=�\ٜ���k}Q��\���I�,�_C��O�7�Qcm��T��s7�s`[S�&󚬗�2��5�k� Q�к�~˕����I_Lۄ���9�Q@�����z1?|o�� ��{	��/߸�V@_B�������ϒ�)�K��݇�q�K������-�n5�𧓊Z|�䡔j�\��X����xY��ϟ���������yK���_</O'�+���5�O/}�eKF��})�֮ͩ37K<�>�S��^�0+�C0G��%`��/S\4�{y��L�h��K2(�d��9�\sJ�S2s�H�Ow���Iw��A&���v�Xt��ߦ]���h���i���Ë��/^�����7��r[�uqp;�����E�����p~�i�}�q/�
��sZ�KI^�j-�Z��sd�^�W�G��OTZ���TOD�oiܴ�RY9��ƨ�$�-m�nJ`0W!猝#H+��1vTص�o?�^2��99�5 ��%�M2|�oI�kd"gtj<r�7 %�sPs���-�wROc&K���pm�����!x�}���:^���&��������V@_Bm��}�κԇ�kb�%���%�3���$��M�
5�(Rͪ��D�$��h6��s�/�+�Zp�ڒ�a|p��IJ'w�\�k��P4�H���� �V��4��T�4/�������{m�s0�'j���$����_������C*_�})Ý�2�+��H�9|�qC��O�i����?��A�����O���>�$8	B�1"�5i�={�e=��j�%������������`vv�j��m��ܚ�Ik�@(i�=�5x��I�1����3WQ�WN���s'�Tw��4��O�`����{���-�o�~������9�Zӟ��D�6r>��r@]�R4����q�)���C���>%��ʍw�`�<J��9x/g�ִK���+��,�.��G����a��h�-�q}�8Ew�c�|�=vZ�;8��F8��>���?������~s������ַ���\��c�{? /`�"��>��.y��as��a m4 0d�������Q��(i�i����4/��D�xwzy6Lc�k�%��ݫQ���4^RZ-"@y�zp���H(]��G��"�x�Ȅv�{_5s�����#��C�ǘ4O��)�9 �i$}����R�0������Q�Zz��{���IF��-���#�Z8�c��b3\;�K��+s��;�h#x��!��w�m��7�ݻ7��m��o��������_������:P��۶�i����~1�a��'�5f�v-ƧќI�yQ��x��1�Z��1��F��8���y�H��Pa��̄�g��?�%-/
�j�O7m���RS>���A7gy�¦������v�T���>'x�PˡF��C��J��LyY��k��<�%��h�����~O�^��(o�7������ �5�ا�5Ɯ �s�|^wz=�K�1-��𕲆D°������Ѹ#�S]C�����h��ktO=�q���+m3�9�zL����=�|�~��X7�������%}�k��:�A
���7��1����ޫ�x�q�4��ڷ��~g����M����'?~��׿��?�7�`��nп����C������������#���I
�o�`�����o8`��� ��0�A�7��ӣ`r���=�x}��FA�s��>R��A4�a��	j}��r��P����s����( �����1��z��&MZgN��)Q���`���աl7f���[�'�[;Dy��i:e���ߚg��rY.$�ѩW�=��@��7� �Q����G��|x�P9�)��uCe?��Ʊ3(��+������]KN3�A���ӍN�:�y@?�mG�ƿ�Q�ϓ����/:w�#c��x�f��B�ɤ=K��1�45�"O�+��pbSq�qy��g�o:��_���<χ�C���vH��^����ｇ�?���Ǎp�o��O�Pyg޿g�/_���M���\�$�z׿>���y����q�������Qۍ� �����_�v-&��4����uQ� ͕�f�;w�+��*��:C��n�Ѹ8U��9IlI<Bǒ�-�����*�����o�A��o-�H�2�o�����g�,fk���4�N�X2��h��r�s'�m0:��!�Dh{8��M������(b�c>��1!{�pG~S�&�(ϧr�jF����������ѓ��?�?5�.]��z�Zt'��|ģ�����@�B�Q#?�?=Z�{��^ȇ׍{�X��h�z4�:1�G=`'�G^�����sݘhTzY��c{�; :��S���~v}@x�|q������}t���������I@��O~����O��_~������_x���w��j����ւ�4�K��� G8G���<8�Q6�̨�v�7�t�ԫ'k�� 9M-���:�����o:�������U�6��s�ӜHF�}��k������;�I�P^,���̋R8��.�F0�B!<T&k2>B}���~}h�6"H� �b�����&P�=Uі܄qĈA�B-������Rl���5�=�8~uC���O�q�z��rp&C3E�І�wv��~ƨdH�m2A���t� �c�QŇ�I�S���E0c�y
�M����{�=F�a��͗���m�wK�����d���I���M;
D�u�n,���ᐓ�=N��&?�R�It���k�ӆ�v�c2��1���tW��Rٸcwp��h������S�e܆��`8�>��O���'�ݦd����h�d�������q� ���䡐ǩ��n`���2C_���Z�݀w��w�ۼ�����w��w�Ͼ�ݿ����O�Z�&����n��������o�|���߹�ݽ���;ۦ��^��[�9��k�^	�j���@庄���l��-�Q�$��e�R]¿n�B �=�����!��Hƶ���	�G4f��>���Оxh��;��hK� N`gc����1M�����5Ӈ���3��nص�j��OM߶�?b�5p����
��c��5�q���m�%��W��9��<M�ARǊ�~@���Z�5����h��{ܵ�1d�[��k=׶�5�����ݭ�i�o�k�
�2�A��A�5�Px�򕵐�v�=*Pw�����:6X��(�U��@�<��7I��Ô��~���;6����l�p����+,x7p�I��᭄��eo}��ñ���n�=�������p�J��^Ǉ�v��A���2$x^t�q�Q��&~[D��q��I'2�n�Q���aB�0@�¼Io�_ܐ��h��*�ow<�)� }������x�C�����1����mۀ1�(~��X���ƅ��M r���m��ċ�O�� ������Ե��&�l6� �Ѱ�hl�hA`CiB�<}�/'�i���� ]_3�V >1|��~<�%z�u���O���?�.	�A�w�qᙶ�OFG���6�fR�tA+4ʰ.��&���qIv�񀾱�][�a`���W/�l����<��M �/^���1�6z�P�����_������w_����˿7WD7�?����������߽s���۷?�����
���>6aPM��`56����\���ܰC�Eiȴ
I.���G��Ȇ��Σ>�a���=f����md���y�C����!̗`&$�J�r�z�)	�Wa~v������ɫ�X�z1;׽:^a���Qǣ�s�c�4���Py�<���lP�[k�d1�.�}��a�tE�� `�����	Q�0P�G��i����m���ءݵ���v�U�<��k"�x���J���������z%	}�v�+P)�s���H�&���
��н��y���L��i�*����m ��}�Mw̭�lw�]�o���h�Ć�;�6���F�����`�$����	ӡk���`Au!��0l�Sz�� �.n�p\��}9?��4ۈ؆�9�Yշh$9���u���fg.��� :��'�'CܺA�a2���Dav�KcaC��@��G_�Ѝ ~M8k4�6W���$1A`�k��&���,�6v��i=������E,Fc�nmz'��ѝ��1 h���Ğ�����A�&�M0spNc�=ON��1Q1�G/���֋�6Lvx����n
����fD�h���A��m:hG3��A���Qko�x��Ϸ{c����y?٘BM�_Bt�c��ahN����%�؆5�� �w��>��I.N�0j��#��|��K�T;�^G_n���m7ǣ���_�	j�>������n�w��u�6?���~���o������M:���J+��ҕ?��Y۷�}�|�͛淿����O��xcj�nk�/��;|n�������}xx |��}��������� z��[��8��{�քw���{��E�C&D����k���, �m4.y+�[�@�}�u�;o�n�������{hވ��]�x<@�t��s���K�Z�t���>�݅�D�6p�[0"��&~����ML]�sm�>��TxӇ7�,����� *b�L�a��#����m�������v�v���m��7�jc��9���~��o��/��G����o���ٿ���B�y@_i��V�V��������_�����ޏ�+��=�����_�����	�?���	�F��_j������W����C�L[��N���x�|����7�� ��ׯ��o��O~g1��-y�y������5���.oڶy�->Ѳ�^���t�sn������GEot��/ �KQ��R��������}�Θ/� �/��wѝo� p�A�����B�"��y�������9���Χ���M���隸�lbn!�l�ݦi�/�;۸��no�{g�/���<�+��WZi�����Ž��s��uw�!� F|���q���5�
�+���J+����qC��nn�V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi��V@_i��VZi���?)��STq�    IEND�B`�PK
     uK\+B�<r <r /   images/9d915518-60ad-41a3-8ee2-5a1cc2d88e80.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx���dWu&�N�x���9�խ��	�Q��� ����ϼ��ě�a���g���`�,!		��Zju�s��n��Zk�]���s��v���~��Tu�>{�su����@ ~�!�.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B��@ ,��@� �.���@ K B���aZ�E�P�,+���>F���[�-�>����7���l7i��֭[��°뺅z�^(��a>����&���<;���|���m�u��8N�k�oO�_�|9��>47�/�\B�_x��D��{�:�}?�u�|ؾ݆�[�}������N:�$_��ϩ߅��=�����,��D�!�p_�{�9˖'��rD�8�&<���gy�c�=Ƅn۾���x�]��}�\��E�;�@	�6>>^5/8�O<�w�	S�Scy�`5�:U#�B���Sl߰����[�NC>_-��Z�rM�Xl��LV6j���a�� v�n4�<��f��X�4���� T�+>���8��3��AH���wͲ�y<���
��<����<���#G��{�)ܿ���;���X=2!tA�Ad=999��C�]ne<4���!�M>�ǭ1<g9~F��^rm�:�Y߹��*�W۱3<|� ���[��|�C��͡������CCC�AifV�+�m�^�s���8�4Ǒ;v�"����Y��0��P��j��
�b0P�~��<�p�7��"T$��Am5J��!���'�:06>>�s���������O�Gm��i������ �נ����ǊUpg�Z��ԑ�ם�LMMM#��y�f��'��v��Ϥ:::�pp����}�����8�D�Zhi�@K�J{_Ә3��2�Ih���0^�y��ݷ���]���gKϗ��'	k@Ϛ�>����?`9|���
^4��Z��0��?p�[x~�C]�u ��O�V;�uB=V�}=�9���%Pj,9
��H�lm�j�6��}�T.�;DL�������=�� nU�k��(�8����	�Ʒ>%R!��X ϲ��ON@�D�	��)���֚�_�9N��MV\��m�k\$����&s|�2X�b �r���y@1b"�bb���6�1jܨ��H��F#|��aٲe�ٙ�έT*|>�/ ���t�h����f~m�����A�P��;���*}���������l�u�&��j��6s9���{48S�繎� +$� ?V�]a���r��J ����9<����x�Q{ބZz�e�s%"G������<���i��Hh�{н��{ı�e~�>���6�~\L��,C]�Y����j����Ma��
_�k�S���& "��k|}-�&�h�	���@/rl+�m�����W*�A�̳��-+�v����,�M M�
��m��U� ;m]Yj�x��g�D�#sA�\�i��������3�S�iQ�&�1>�h?w�u��������s�ڵV�\	�Q�����g�Mm�@�?��s$�`��4�X=���x�>�me����A�%^�l��-M�-�<��չV�ڧgP*��$��Z��=o�|=V=N%셭���2
�ԛ�_���(>AF!�.�2F����_֗��� ����L��2��cǈ�j}k��s�5�f��z�ӧ�磀17������?�*�xM��� ~�F_��[�,39A���4�G�Sm���j�\ȷH?|6�6�D�����l�[H� �}�'x̃�"����k�&kD�:nR��"��C�\�ǯ��c1?��L���$l����4���U�Ze�u�$��|N�o���>��L�F`u�>7�O��宪T�����AF!�.�$HCn6�7��̜�D9�5)�'E��qS�KDq�}��7�HjOktMZ{֤j�E�W�����	���f��;��t��I�e-��ۡ�9NLL��JD�}�Z��Z�ٶ�M�H�>��纎/���8}H�65b����5i.HJ�{�k"�m��Ҳp�6LB���	j��ggg��cwI�� �BdS�3S�W�Q2��1s69���I&`��1_��K��?��^ڠL�f��a�N$\��
m���$J4�����6;ډ�نo�4Yk�:���m�me2/�	��k�;2:3��p��6��~���d�., �$���1�Q��d��v)��Gs`!�r�F��]���>}�l'9*1]�7�[�		6��� r�X�u��}QsLqp��E��AP�L!tA&!�.�$f��8��-�CC9��՘9X:1D��ɏ`�I�f;����$�v4��}�o�x���=l�������4p�jY�x�N0i��H���hw7h��[��k[�;,�7�?n�蘇@�Y��$8ݐ֮���
��c��D�!�� ��#��u�8p�$��� ��6�s��c���#B��M�T��/]���~π¤[&k>;[���^��C��##�l�4u���ȧ�p��f�HZ�|��!j�D&�t����4~&�@���6����x!�B�u �m�{�����������+˶�~���?^�:�汗/<�:��A��Y���8v��:�m��B��G���W�K��t+��p{X�� /P��''��B]�I��MQڬb+Q�� �4���f�S|������F��<I�#.$$	��U�]�����5c�S��%����@��:���:M��~�ڹi�h�4��>�x�f�m�m�s��&�:'@����v[��vt�m�rEwll�{'��#��لC�eۧdp����nE��hsOi��_���5�EF�zawjc�/�������n���D�F{���2�����j#so��m�Y�~�������dv�`�(?��_i�k&Yƣ����^����ײtN��3?GY B��߮#�D���%<-�� ��1�v���J�7J{���
Y�� ��)�*^���� �N߸I~m�z\C��԰酟��Fr�~��V�P�($��(r�۶;5\�'j�|��Ze�t2cl&��S[��S{����vK�5���ǵ��6����a)b&ÿ��g�͋
x�ǥ}��YuXP��H��<'z���h�d����y��^��@���ӹ9� �Bdvh5�0�\;ǹD\�;TiE�}��w��*O�UP�G>Q��mE��mFr�A�qX��m�֤����f���ճ�h3����J�a�-��¹՗}@����IJ5��$�=�e�ф��u�5*mO�Fh��Q$st��чƮ#S�O��Rns�)��<x�R����꣟��,&D�H�NT+��"@,(Yʗ��L[B��D �b��5y��Ǳ�����CID��3��-Pi��:˅���X|Q�Y�� ���M4#����A�c��ǡ�S=����e��B���}t!>�^�t�ަ�ʻ��M�]L[:H����m�0��R��`�*��՚��V�{4�'��c�+Hy�a�?4�����W(d��R�U�Y�2Ӝ K3��'��)j݂�(¼3Ū��=�����K���-p����z�izFA��a�`�#��9�9��m5������4V¾T�~糧n�9eB �(�����޴�&#3����N�v�x����]��X�=�����M�5�:�^ϩ�3]�},��k7҆��Hx֡e;�	����� ���Kf����	+D֛����4�T5׎��xC+��jE�x>0��k��8N��k;��̃jq���V�kT�]�	�`��,A��	5T¾�:� Bd�C׿c&wB?/�㩥'���}��ꌤ�'�^�v�)@�Ϗ���~q��X�V��]O��L���.�i����q�+O�Z�� �B�_�a�P�X@����.�f�o���=��OK��"�#��1A���Klj����|������+ui6��߼3�^��w�4�@E�k+	o��5�F�u���~@&�ж)4^|��B]�I8*�;4�reڎ�VA��;�y���<04�c�g������"�Ŷc
Z���Ε�N-3�
$������x4�A� �.�$
����~бz��kӧ�_��|N�2L������۶��o��V�H<.&����1��^���.-��s[�����K��3��G�V=����zz�X/�J�s[��uQ*2C�_��z�׸��l���׿���;����i�h7^�ki���,�E�-�xQѠf�###04<����)j���Ael��9��K���qݷ��
q����s�F�"�$׋��׍�!tA&:��/� �\�Az�B���%���w^ऽ~���2y�K��b���l�|�^��{��8���E�4�/�P�G�^��ʆ.[���Q�6¶ N�473; ^�N���˻׿�G����I�e���x�h����ЌJ���Q�Y$����(�?�<�(�Z���:W�������{���./�:==k֬�s�=NܴV�X���>�G��i[��h��'Dc�	s�%8�z� Q���� �pB���!�����U��>""vҮ=*1�0_��r���h���k���������������������>��O���;���n�[��V����v퀓N:	^�����٬��O��=���U���R����m��M+C�O;q��Ҹ�&�W	
������ډ�����˹/�������98����s΁�e�059�ڵ�>�<<��ðn�:��o���w�z�쫧���p��a(bۤ1���J�v�σ.��b#�ҷ��d25]�Y���0���L��EKZ&��K:S�z�����H)�/�v�@������L�?��O����6_|��p≛Y˦R�������|��_~6�t
j�yx�k^���'��	?���e/{��y�|
���7<<�[�2���َ�wۏ�8�b���{LQ҂0�z��E�H{.� �kГ}dz�-˗�������?�|�߄���8��]/�/섇{��&�Bx��U������^�����3�8�ix�{��x�;��+^�J�����:X�A%�C�n�A`���� �Bd�E��M�&L�t7�|R�����Ԫ**�����9�Z�^�&��I�^�~<���۷�9���i�ܹ~p�}L�+Vb��O<�$���p�QC��7��Xӓ��Y�1��KEx1`���Tup�I�|l��FVnǆ��QP��i>�:<Ώ���p��wþ}�`ժ5H��u7����۠00H��j��"�����I���{���ч��3�;��o�~;<����|�}˻��oz=��mZ��[ɫ�E]��sڂ��|u?f�~�C]�I4)���öf%~��4Y���^��3���%�o�T�� ly�9���;X�$-�������Z���0�N�y���Ӱw���:H(y$��~�Nx�ga5j�dM_�z<��,\}��p�%���3�h��En�ݏ�o��Ed���n:HN��Y=���nך�ȗ��H����TAo���੧��kO>�T�����9�p�ր5'.�؄<�K�2L�b\~��p���@5��Ń喏/���˿����ꪫ��h$�N��Θ8�Ft-���B�L"��60���AO���ť�˓�����l���0�=��p��g����o����o}�9g�y&��09=^��
dD��Fҡ���b�!��1

�9BU�U�W«^�*x�-l�'��ר���g�Z�Ǐ/�Q�fp\���=�l�\��:t�����?����(�
ES���ztt�8+Q[��V��Mp�:2׼�:x˛�w��.x�k_��s�>�:82����7l8�S�/:��\�!O���a0}.�#�� �.�&x�L;Z��� V�5�_����nq�4/+�8�L����w���u��w��]p饗�'��o8*��-OA��Dl�������7�	I�A8�y}�IX�b5�ر�O�É'���&�Ծ���޽{��֢�ND��T����㪩'�"3}��9���hdf�7Q���a��)�7�|3
2��o~�v��]w�\ �!����.���+X�'�<�*��L��������}^r�����p��Sp��a��/��28�����Nܼ�����'Z�L�\,�mkD���9��o�@�s�� ��q�P��;ҹ�]i-N���Z����Z$���,�`Skd�-���	�Οy�i��}v��	������΁O�oᓟ�����`�2��s�,�j�'�r�u�Y�w==;G�xv����/��]Ȥ��č�G�pj�������#��j��.R,}_T��p������Q�1���m��1�,�I�!���m6�s=^܏r�C0VK� ���&	I97͆G��(�}?��u���K��Kpι��o��;���L����_��+����a��+�
��Vj����!n�n�zؽ{7�سλ�R8I�"�à��֭��O��ɍ�|�`A#�
e�H��? �uk��Fk�;x,=�\ϭvWXM?l�BdB�L"�*q��\oO~	�fX;s:M͝>`��r��@��s��y����>7�t����I����Op����U+�0n�޳���s��lt����M��?�gp��87{��5�����/_�"	���)\x�Ũ�7�`[��]�&��`�k�GIlD�����$���y�N�`(A_�u�V�D���o�����o�k������:�ֻo��{��<ߏ���ѡaX�a=���]/�ƍ��SN��_�b�|��5x��y�!�#��026��z;\~�%<_SG���(��r�i�^}��2�~�5ObrdB�l"tY�L���&�n�dIDg���ÇO��4>*xB���v�G�w~��8����\p<��#��	ݧ1����	OB�{���]����������?�����_ع��
�u�K9B�H\W^�R��4�!���Lm�",���M��8s�z��
���R�Ô˃|-Y>��o>	[�<��?�� EZ9�����#j^H�q\ry���#���}Æpꩧ�SO<�L�������`���0?;�ׄK.� ���"��:��oBi�Ad���x]#�3 �۸m8��x�B���Ro�nZd���o��vh�� :7��๭�X�������4B������#��?�W0:>
�P�&-�H9g;p�9��Q"��+W�YyӦM�7=���?�������04XfSp��d၈���P��AkR�0�ޜ�$�I
��kB�fm�P�-vO���7�}zz��'���`zf�#�I���W�
�׮�[n�J�>�����Ffv�������{�z���LMmc��/����ڵ�~z��s���"^���*��ۂ���:Uq��֟X�����	B��l�AdB�l"��c`�F��l������k[����,|����X�����Б���!)�^�j�l߾�#�7�|3�oXw�j�n��u�8 ���q�i�.��ܿ�O�X+V��g~�����+�@l8���8��"޹Vy�A��H\�����N�:S�1�މ�&�ʥ���EAm��ao}�yص{/�����V�9��/��z���o��_qx� ���9��2���')B`���3p^صs�u��Y|>;��k���������(������P�G�fZf�����<,4����Z��̐�hn|;�<tA�!�.�(�V�{���
gI�h����J?�>�H�8���>���Z��ӨeVu&&ʍ~�G���+P�Ԙ0t-q��N�{ڦ���S�47-8��ÏB��!�-��<xv��}�X������L�EOb�f�����v���q��}=632�)��
�!r&��9�˿/��l>�p�	<'�q?��J��TX0���+�Z�p�܆u�y�ʱ��!�b�Y�~��Q�!���={������χ�O?�9����O����#�;�g��v�����t���*�� �P�c;)-N����7����y�&�z����x�g9��G�\��� G�7�>���������e��4챉1��a�~�%�""��������s]��<j�S��׏�C�s/އ4ˡ�҂൤��>.�ӮMRRB��!kB_�z��}4ir\�-2���ٷ�|o^����·�[���>���uԚI3�.x��敯����m۶�vM�t�f���l>�M�5(�ofr��a���a�[��7�Y	����[�p:z&��L��,p��=�ZW@��K�.�ۉC��t_�U ��C]�YX�7l��|s������n�)�驢$����|��g�9TDf�j�G�r�'�`��&�#���Bp����`-�ͩeBI+�\t"j�27�dt>GoS	S
���w�Yg�Ãe��jm���a��B��i�h6�q|nWE7���Z�a�"����FZ7���~�y�D��{Nn"k��i5�Grg�\L�N�u�/b�]���s�jY�f��sY��������B�w���u�?Os�-F��?WL5�ǅ���$*N�i�2�<�|˶�����\M�$!3��4f3?���\��@M�����,��&b%8����AP*��� ��ɁZH�D ;�m�y�8O>�d.Ns`�~ָi�0�$�
 V��x�!n�����_:NAy�mj笁�s��s����}/q�:(N��5o�y�[�y�o�;�F��!�)Y$N8q���>�1����pCes�򖷨�u\��ݻ�甴o:^mT��N�ӆ���G��6lbA������議|�Z�޵8'*NC�jzfV�b���u�M��k����3�$k� Jׁ�m�ҩ�LC]�I�9��z=ϋi���I�4�ۖþޟ<�`+oy��@��@�o5�g�/!y��/���LM3YyA���O[��In��k攚F� ����?{���r�v"3�ցp�h	Z I�8O2���n�iG���U�N�[�z5�����k�l�r�$H��s�w�������]�Q�d�&���a���4T��#����G}��ٳg����6��7���
���צ�{�>եv;ۉ�a��ڹ�>�1�4K-�A�!�.�*B 8f�(��	D����cO>�d��5r���K��]Ț�s�>���k�p��Aoi�@GZ7oT�\��=ػo��]��T@~���ƍ�0j�N�#C�܎6���]i�{�<��5���z�J镛N�j��Gn�Vlެ����N� �'��{��u6\z�EP�}��FAlԷm�o��gy]t���,"hx���6���(���eШU�/�wsLؔH����>r;�kdi G����޶�k��en'͹E�]�i�2��h\�M
�J�pI\�|��ܩ���]�R��7�� �]x�twl���id*&�qdd��E���{U$|���LdMDF���m���?���Hzy��s޵��(�H��� ����\,�����7)(��b҄s�*�K�F���
LL����>�}�G�M+��q����W��S�Ɨ-������G`ݺ5�W&s�����<��Z���o�`����Ͽ�\��>�@�V�g@���3�:[_H�h"ٷ�A�R��+ͨ�3j+�����}�<tA�!�.�("J�#8K���~��~t�96>Κa�o�f8�l�Ie�	��m�
����k��5l&3��?��~�i8�ʕV�g�����+V����[o��ۣ�@I�a��_��9�a><8��Eį�[���T�nc�Ͳ�<3ںV���~n�@�q��dRo4�lj���k�¦� K+V�⹣�n��ܾ�{aݚ�p�E�K���,����nA�����?��F��j$�}���}�, ���(<�z��p�M�w�u'[O6lX��4/K�!�.���Рa;T���):u-���f|����H �yB]�U�����������ؾ��._�E^��m�C�{�.�2��n~�Mp���s�WJ;#¥�*"�-�=�u���b4w�}7����5���?�?~v���>��P#(#�����$<� `�I�}�塗�t�b4�n0�mI�\��9��W.X#oxk�$̐`��3OC5g�����8��vs0w� t��=;�|r�BV*�K�
J\�z��U``���n#�LN�*w�V.g��@�k��7"�xP%�lg$�%i�I�����X|˲��.�,���08� �$4�B�C�a�zNg"�̵}���g�O��O�t�z�r=��I�&��{8���h�4����7�	�A��뮃7��F^K�VL�Z��Zl��������.��|�.(c�k����$��<N�i㏓�b��<��MU�!&�fŪ�p�%��|�#�Z���x.��؂1����WE{���'��'>��/�ê�k8Ӏ��(=�ș�����d�_�½?�6m�j}\y��z��`���U���v��7��&v����CoV���� �Pʪ��g�DLZ$�5_��N���Waj��>�����:��(j�����?{���r�Ȧr���W<X(�N$E>��N;�#�_�җ�c�=o;�,�U��دL���7������t�4����8��O���s�v,)m-���k������� �����~������և��k�D��r m���iܟ���a�S���o��7m�s����T(��M�L�K�:���o�n|=<���Q��azn�o{.{��l8x�0��u��w�"D�,�q���@��{�?�Bۑү�LC]�Iü��-�q�u����i�jM�6�S�^Cò���u��Q��乾�Q`���`��022�my���w��M�y��B��_X������uP��+�W��Z�A��?���ֳ���;�W]y%�s�=�m�V^:���+.�u�W�^k�m�������ڠ%Fi�s*�Jk����븣���Ͱ#
�I�Rep�Ulx?Uǣ�T��
�����=mҧ��G3]��^��K��u�����y<�����
)o��}{v�+b����w!�����5�y���/�;w~�s�����'��ul���N?�t��'�F�sρ��A.�s������~�x�x����������Gi�֪?��M��`�����v3��Ys.t;��=:�CdB肬��'?�2Z뤘�df6Mצo�	������Is|�[�
�z׻8��;��|��_���~�5O�S^:��)��4B"'�S�}���y����N�[���b0���_�5����{$�?�ݻ�@1���s<0+5�*�X<��`��%E�w�L����UD��!
$�h�C�,}����{衇8m���%K�m�݆Z�p�Yg�&�̿������v�j�����y��{Q ڼ�D��}�]\��4r�b*6s�)�Ae~I}�- :�>f]-����,�f�0�BU/6C�rdB�l_�[Dcd��WO�2_��mj溘�OD�$S��Ù/9���r&�����������+��I�/�VJ��g>�n묗��Z)	��qS4���q�q2ۿ��/��}��������,����atxRzU��6�kėO��ޚ#�9i�I�ϗa� p�9��FCU�+�
03;/��R���~���W������;�n
6$���?�q��Pⶶl�����;���C�}��p�	\T|f��5܏�N:��/r��6��Q�:�w��գ�5�������8G�\� !tAVA�S����I��~��R�f�<�^L~s�w�y��#��W���6	DFe�f`���f癴��H����T�4"�/~�L�D\�&���u ���0k��_~9��y!
(K"�|������n�{��M
�K�Smv�y�S�g�z.�]�Υ�޿��o�2���k_�Z�'���:�`�؁j������9Z�|9�3��kp�.��R���۶����|'�ի�<���_�W����蛴w-��1iX8�R-N�m��	�s�ڪ�m�W$w��i�����f�r���R8x`�!�m�wp �e�];w��B(���i�4�LD(d�'�#�~�'؇��~���?W]u\��`����SȻ\u�y׀��i��	i� ��'E�y�.>���9E�xh��"�c�	�z�����s��/}�������?��;��Uݮ���F��Pq*LS.�=��[���*�����}Aah�V�~�+_�J�� ����?T���V��YP��P�!��Ȝc.�ij}h�Q��O&�� �H�%���I���#�\���q���y�ԑ�h�"�o�n��+L�b����O?��;ab�J.K�����	��������KZ��C���p�E0��S��E]��t�\�a�!��g|݄����y2�w�b���aZ8Z�j��i"yR[D��~ ���/��/���9���A� C�uS�9i��3L��8唓`��\1�ڡ6h�ٹi.�C���|�s�c�gΦ����^�F��X��u&f������dB�l��,�|���Z~�(��2��}�j�p�V�e�IT���
�P�x�T�� ���)��|�S�Өu�����n��O��#���sЛ�5'�����M8��2�S�2j��/�W��z؏�����C�^��򫦀�W�#h���H:���E�6��OtX|o���s��ui��麏|5
Ad����y.�����t�`N�V�?���5�\���'��	7� k������O>3{�+�=�ȃ��F�鹝�i3�p�p��'�T�8�0�*���!:��Չ����W�[�n1浗��	JAA�!�.�&��Z���M����AqZ��ڙ����z�.�nB;*�������g�}|�k_�(m.e�r5�_�?�|��+oa2�6ׂW��Z �LOd��w�&�������K�I�`X��PO˹O�)H�l$i�$k����jMm��iZ�֫�5�[�,�2E�_r�%�O�����*y��	P�"�����Y��؄f���x(�}~��m��f�D�'m]ϝv	Ї�����~�:W�sU�o�sc��,�"�6����P�6硇�_۶v2yF��V�6�;�$wΙ�̯�q2�v�ףjEAh�����I��Λ��6عk�����l:���7��]z1�y��L�D�]r)��i��͛6q�����L���� -3uNk�of�C`�z�;^eN��~c�Kn��c�]Ж	mn�sG�Hۜ��G�5j�(-,Zo�.Dꍀ��4���{��ﺅ�"J�:�O?�Gů[���ꊨ�n�Zn��O�k�%��
W�#��~����D�z���yl��skBoS[�|��FB�2!tAF�oݠ����V��������OD�}�^�>V�4�(�jtd�#���*�|��p�-�p[*^�-'�;���)R�H��\��1A��ij�ȕ>Fĵ~���&Ң�M��2Dka�ƞ+8ma���hn�aj�:LN�Q���6o�"�=Ϳ^���"QJ�k��eZ���M�!��M+���G���39 N����� ��l;�E�ҡ�5B'9�+t�ض���V/찥��G7e4,�^#JKf��27��6qP�:U{#3�k_���{ciBT&�0"
M�Z��uڣ��n+�i��-7�������I����;,#��9���B2ë��9W�'`��o�0�:�+���S{H�q�I�����<R�A[
4�k�C[Z�Yi�I��p]�A�!�.�(FB�q� ��Z,��N:�`C�$��	�5��"/~ �TQ�$�z�	�g_�� Q� *B������M�q3{i��M��v�F.��G<R>�o[�s����-�OJQ3	^k˔��ZƔ������6���-?��gO�L�:����8 ��D�����5jG��=K�9V�xa��Z�LC]�Y�*ʝ��=ɴ���v�3efS;i��v�ENwX G�dG��E���oEXs9���9�Qz��dC��TT ��ES�e�qF�y���Ȩs.�S��y:e+��2���	@lM�0�S��M�bڋ��1M�D��B��(�T(p� i��!R�ω-�i	q7"�<������D���ѫx�ݞ$H���&dB肬"p\^�*�+O�G�Q<�X�A!�9��"*��&嗓?W��F�D6t�����-J�#F���l��D�H��oq3p\�6I�h���4���V����A�~��4i-�p��s-� �^�����ᖖM���t2�k�����on
G�A�0[�F�>����u	�dB肬"@���m=~Yw�b��]s�_�V�`M���Ky�d�eB�#����Z�T>謁vN�"soI��D�i��Q[��a+��9�K�I�h&������������ۡ���\J׼��\�E�4T����9��BK �oz�����;6�G~r3b�Sà�/7K��/���
��76Z���LC]�U��"���\q��횦w���$f��&#��j�P�)jmPk�0�&m�J���S�p�^ZTGٵMߪ�Zc�ef?���[�Aqiי�����~j[i��o4:#�yU�ȿ�;P�>e�P��do.�C���>0�sG��f���i	]Q�NK�χ����c�Pp�������� ���C┟"b&�s���Ya�d���O���U��N����i�?��E���d=?lEv��|��pך��AJگm��{iÉ�V`���{�*�YQ�r(t��u���β��{��s��]���"����[�g��4��c���D�o��}�lR�Թ��|GP[˺`EU���3���b<���I�t���Y�T�Р�F�
�B肌C]�U��5���&������I`Bv�>u�c7�Ls|��>d:'ZS��"3���'��'i�qk�y^���:��vA��q3����~$��QW4�����Z�m�?����n|�V$�.�4�����:�j��~_�I/�vp�ݪS�n�d�j�b3亮͔5��bM�i����k�E�ٽ�M8���ì2�糣�vI��C�ב�#�06�G�g�w��C?l�h肌C]�Y�K�Kť���i�F���&y$�����_p�������'�%�n�M�g�۬�ޭݣ9���혎hU�;�ؖ���|ƭ&�;�ҭ4�����4M����k��M(K�WA�!�.�*|��fd6�����"H=�nf�i�]��5���z���5�ϊu;~N�bǓ��i�/�B�%ͽ�<�%���ҳ���~m����Fn~�uA�ۭ_�E���G� :X@ �,��YE�/� N�%Ub&�$�w�	�}���g����sQ���'��� �i�նB}�	q�h���mŉ4�\�]/��>��Zh�I�l�Ǒ[�	�P��'���B 8�Bd6kE�H"�4$i��|�����n�	$d�"����ٶ>�#�i#���)};
�襍*B](\ġ�u��i���wB����B0����������)�3��5�M��{�/2!tAfZ!��CM<I�K���c�����v��&eH��&i�t<����B<& IsN՞�l����� 9�=�z ar�a����Ǫ�'�b�����5v�C]�Y��n���˷��M[O��<�`�$S�I�I�'�x�i}J���}��i�m^���Q�i�o+�/��$�y���,���x��$wJ���4+EҶ�*��'Ӌ��.�4��م�]�:.ZdF��ԗ��bG�}��|�I�/��Jԋ�HD$��r�nHH��(E.2��JP� �Bdv�>�ė�~��ӌ���'�Ny�/���-H�����.[����(�^�Fn��Ŵ6ĵ�^��.����h~���ۋ�	����>i_��?��g���Q�e5@]�i�2�0z�������jc���XI=n�N2��ċ�P ���?!���	��&�!H���r�:��n�HS����UZ�o��!tAVA��ay��t�K^+�|����P5ʩ-_g���(Z��.���'�yZ@<� -&!>�Z�ҞOl8�z�Ʉ����3H{Fi�M4a�
�]�i�����^�oٸ�n��y�m_�	���קEH/ƿk�w�}��$7ֽ��=���ѧ���5���Ƿ+�u�(��J�;�o[��\�y��
�pO]<�׋Y��f����E��Mˍkǋk�3�o��"�_S�9�{���4�w{VqA��K��[�tm��b`ZXL�㶶�@��!tAf��߹�U�%M��u<�ضLrҁp&�.FCW�F�����|��O񾥞�c��v�R�v��v�ZR�}��en��c"n�1�n�(�O�}+�� ��2!tAfQp-o6C��q�����,��Q@$���4�V���گ\��bW�m����}�!�h�vZ^�0��z�6��HB���jmǈ5�6z?�]L��V�ch��~:�Y�P��i4�R��K�ҽh�@]g���Z�m�Gぅ�ȩ^�ܷ�d�>ak���k������yq������5ѓ�L�5�A$4Һ�;8�3������� ����l�u}Sc���*b�̮I~��i>ޤ��j��>]�%-Z�����Y�4I�m�
g�W��Gu��]�9����z����� �sk~4̢/I��]4�J��crw�u1N�=���G��6�A�Z/z�x���u��%'���P.Ӎ��.�4��YE`Y�!|	7����z�Iē��5�}I�M�A�~�b/���z5�^Az��kӄ�&xh�FY��P(�Z�`bb�ϛ�����!��\����G��O�[ײ7��.���5Is۾ ,K���NsA��H�ћc7�A�Tm�'��ܜ50<ܹ
�@�A���0�8�H4S#'��$'!M�$�yY���x�o8�^�|�Z^��5���� &a��.HC���и��<��#C�,\��{ҹ�ڼ�Ή7�u HCS J������l��fj�R�d �,5�뿡b��ٖ^T�R�*�P�/������L�@�Q�2	|������J��6S"!��Z�x�<�D������wO+@�����������h��̾�"�0�ɝ�����?��ccc�MsFZ7�&h�f?�:i�F��x�jj��p�y~�X�6���$���2�q?|�ɝ,$x}�\���fg�ۻ��@ � ����8�����֙�eJ�	�$�$M݄�/QC��D��;�o�oS�H"�n�mI��M���l[�OT{�ɚ�pxxj�Z����ˁ���6�߽,���>s�;i�7}�f��:�ns���uN�8j�v��<on��aם΅���,kt��A]�Uff��)k�/���ï/���ڇ�6�7�$$�C70nF�#�z� =m�dtO�ԉl7o������.�-�|R�;k���=m��5ᦝ��nwR�:��eIB��F/��L�����5���`d9N���j���Z�*�u_�T}w� 3Bd��̚�����Bq�^���9�G�Zh<�J�$�xnw� ������'�O<�,-H+�?&!%�i�\���<�
�k��_L�t:��S� պ��9wi�9��ؒ���@?�\�.�^z���f��P+^�m �(:Ǚ��:B��ra�'x�s�� #Bd�ٹ����4�R�59XQ��~��"��(�^�g��q����r�{�篃��G7T�9��b#�F�5�����h�ڏn�JI4�7��nq�N@/HRb�-h���vM7�I���["zV���ZJ ��y�=�ޙ'�?���k7���u2!tA�/�ܾ��^�����R�r����7{�[�h��9������޴���n��5?��_����$�~1v/
�x�i�)���<�eR8����F�qn~���� ��W�Փ�[G19��ֶ:���B�q|�X?�5a��&ߏ�Ы���0�'LE�f�~����0���I#ޤ�'����#Tm�����'�|k�Z�X����+�e�j��؎�@��2���7W"�;�E�5t���7�Y#��zi�݂�L�5���z~?c�f���fj����yNڜ���b�ϳ��O�^�4��>u�u0�d������Fk�X�l���� ��,�����~�jͩ����䠪nZ���M��v,��Š�0�K�V��mc���K��5~,�wG[п���\�oI05rSHH�ԕ"~mdh���ߢ�,��� CBd��/SG���N�{�W`W/M�:�X��f_L=nM��O�[zYt{��A�����/i��s���ԽZ㏹ pXn��Um�g�2	�vZ�R�x1z�}����|����j��`1&y=�j�������h-'��w��;�^�9!���	���!/��	!tA6a�a@Edh}�Ҳ"=�Kz��=z�R���Zo� ׊�Lo
�,�r��������d�[�k�^a�yj�m-#���h���^Y�k��]�M�Hs��t
�&2���� �z�K 8Z�qE_�$^ih�fP\G�@���ɝ7@H]�)�2	?� �.tT$3�� 1��_��Ť}���S},(&��︊�}<�۪(�c��xHKs�ƭ�Z��]�g�w��\�^�3�Ӛ���Sv�g-��k���i�rG	$n���?;-�<'~�4�s�wߣ9�<~��
z�Zꬣ���S]`Vbk��H
���~�K�����4A򲳽����=��F�V���E��z�TS �E�Z�T!�r��lA]�9̂҈[�VF�d���4v����)��/�>єd����൦l��u3IY��i�Z��Z�"�;�R�`!��Pu"m[EB�J�;p6[���N���������H���Xl~ҵ�ڏ��h5�~�-��~��-p�x�0�:��ض��`�@�!�2	��#�$�����-�'b�Y�.6H���	�y�xQh��'Ҭ\|�Z�=AҦ��dIKS/i�g%,��x�)(
��F}��gf��iW��?mX�s"}.�Yp��&��O� ���%�M� ����"滙�����i�7�>ڠ�����Ð�w�4@[J�
�!tA&�D&t�$[i�T��4��j:n�]�)�f�����Dؤ[9��J�YP�!�|�ͤg�J�7�Ճ�e&�Ѿs�zg��p;:�!�. S|Y,*�"@��0TL,&Э�~M��w��ދH�i}�B��[��rx<��r��[�?��2�A�BdC�B�|[���o�b�ޥ|�*��964"h�m[L�Y[d��U]�&^����襌�u�W����'�2(b֤�$��5i��G%A�J����Q����)F��t�8}/h�����Y�K�﯄����OTw��qi��������ԏ&��h���������
�2!tA�0gYHζ~_Q�y*��#�u2w`�U/2�ڊt�
[�/-��9�R:��� ��*���p�:�ҁ|�6k�(?���;,_��$����`7M:Nm��x'����|
�c�,k���}<�]�_,����Z]�u�/m��ܿ�k��@�neDr�� ��h/��(�ˏ��5_"n_�)m׷-uUD�D�!���r�:��]�UZ3Rk�;��N{��O&�h���}���)�-��s|�?�{�9��u�����I��r ��������٬�o�9�	��M�G�7M�G�Kޯ){1Hnka �bH�[P�����V�c^��!tA�`��J��q�L�A���OߩEdO�ʿF&��)�Ȧ>ny�_��Ƥ[���
��`.$�*��N��FBB���i�nL�S�:if�ϑ��k�}+
���z�G$���pT;��qߔ��H�&���ʥ��>�"*��z�.�d��5��i�ǃD�����kގ���U�m^�OL�LA]�A�[�c�r�����=������}x
�B�I���H�y�������Xa5k�y�k�������rz~t j�*�*���(�(����R��~�r8O��T������P�oԡ�����:Xx_��T�P^13A¼�S'�<�P����K���Ck�	����N�4)����,����cǊ�v�ɋ�$!�dk�?��nB �7o�jZΗ�Owl�`PBd
B��a��~��M�AH�$l+�H�/��>������a��aY6S�T��B#�ò�Å7\k.� &��������>����S�E�كӮ��~�[ _.�deV���=�?�����e��jP>m���B�D��?�S��`�wT`iq(T�]��9P�Ф".�"4Q���x�/���p$�Gij>8���U5.���

KC\�=%y��VacL,<��	�!tA怄`�vT���~s�.!��F�8=V	�6PkϏ�7������*�s���&Tw>w��Sx���_w4��۴�8�lx�߄�G' ��ã��e���Ӡt�i0X��� ~�o߂�ݳp� j�H��k�����0�c�h�\a�[����ˁV����:n�p�6n��Ovm��������A��o��Gis*S��װ���^��:	�؂V�52+�wua�'t#K� :�q+�Q[(١(�.����Օ!�.�Ls�e��Z���.�����s�G>ts9��y���n���T�$�RŃ}�6X�yPq�<4׿�P{���l�/����������߇�U��x�9x����U�'@�v�����+a��!I7�u�|�c�t��.s�)p����m�����U�g�>/��\=��z�6�_��Qk���V�ݘ������Ʒ�~��w���b�;^H����Y�� kBdTd;����H�.�*��I�҇�*���r֞{6\�ΛQ����{�~�_a=��bt^8�?�,�^}9�?2	k��Ʒ����j�c!^��x�g��o�����!�0����X.|�L��`�
p�5�@����`a��C�� ز�����0�0~ޙ(@�$
%�P 9�Thx5��^l��P�o�
��>�^��m��~��w
��Γ��$��q��Z�	�"�Q ��@�-���Z�v�ꆖU*�� 4?�&�e�CBw���~o'�;TX��X������~ �=�`8�Gޅ��,+�!�zpdn�O�W��p���7,]	�V����!�����q6�F������=�����M둸Ce�y(�o~+�<��y�[o�y/|��O@�"S{�\��m��y=�S�sj����j����+�9�Uc_��'�R�ގG��qi?U���\�D���c���m�<�.`�����@]�9�K�r�Ц��:���Hr�v��`�`�l�rkP��p�5��sx^�'��6`hh�{f�5Z�������a07����W�3�<
��k�"�R���?x�Nl��3n�Ʈ���J@�jՇ��!�JP�:cCðǛ�y�#�k��Y0����As�UC~`��Q�4=N�s9U��;z7,��Ӎ�I�d�7�:i�����p��q��,�z�-��z
~�A�U{��2ˊ
���8�O����H�d���V���� j�Tnz�.���$Goj�r�#�A�+�^c���9l'�*��m�������Ai�	k�<L9�}Ge
W����.NS�lT���w�;܅C�y$��`�š�{M�5�P\6�������Pi�!�pa�D�>8�����Y(��f���x�'�G�����W�h��1�FU�#�F�(��UoC�j���Z���&2�k�2?�Q��P����yi�?G���A�z��H�͆Q%A-E�.dB���*YM�;w-( �U*(�B��P@�����b^�����= VށU�1~�n�<^w�;�+�y}�F��
~	|7��������������Їee�N¡p^s�{ �y�D! D��㡧O�哻PGB��\�������|���;y�oxPr�5�@�o��<_Oy�4��54��)C3t�k�s]{�gcoΥ���(Tp޻�|�k�(�@�����؟��b?r�D,	 ���C*�U�Y�R����\�Wϣ�:�7�~�a�Pt�UC�o���}�p��9����,a+|�K��b�����~~B7]y�ծ��7���6�p�����n��
�B�@-�CŁhl����/DB&A ����C_�M; �|��*�J%h )��U(�&�"AS�[,����_��� @�zr� �G�ī.�k����	x�HL��.r��-$b��&a��ka�λav�6(�ۻj{p��g@ἳa.h@�.��`"��RE�Ki�\d�Q�	i�sU&�n琌����x����f�d8a�Jf+j���fH-Gil�`��BǢ�L���v5��z�K�Rq&v:��k�*�J�uZz����DćĞ+8P��P(Y6<�U��^�A��+��� �[8���0�F�������*�?~^KN�o|��O}k�����7k��}�����y�*�9(�3�\�U��t�f���٢B��*���c7G���A]�I��re"$Ԍ�>�)�4(*���H֧�ݸ���W ����9�n�2��W�D'��t�/"�"�+k�� �rPm�ayq���q= �7Ch���o��J�Ņ�r0h�X���f��:�<i{�6i��^=6%/��[�D�t�G�ښ,�j� i�\*�q�T��~S���	����a�75����<k�d�,��ʵ��6��4LzUX�r������0߄l�RIWm6j<_�n���f=m����6����(3{�h�c�� `ot�Ѽt��8��A�?����s���[o�o�� 
�(�����8���u�~dv�M��Tl�R�j��?�BdB���k�p-�:��Pf���=[S>G����һ�����!D���/�F͇��!��.*��u��r�D6�}�����ldf*�Ǝā��*��ɶhоf��3A*R�v�҇ʸ6�$N<�HI��>nN�����(\�^�?������񺇭��6٤�Q:5l����N�峳YI�lO��������K�0U��s9��&�>��b �s۴><�oO��x�h�|�_���?C�uB��C�H�p�U���ل-g���F�&p2G�Z|��^o�2��Z�N����8f��iJ���5�t%�x�x�w}�<���ⳮUjP@����.ذ���^.8�l1N$��{��3Aes�W�2�jX~��UT˅9&���9(:H��B.���ėkyp�v�M�S�&ԭ
����/�X�+\�QE���G�Y�
=�By` ���;
��6eֆ���OQߴ���3�"�
P#!�E"Ķ�I:�-a�N��%�G"f)e~rV�G�R���D��$l��������1���@���Bs����9�&?���H j� ������W�Sfx�s��.���P+�v�S
c�4���]F��U���M�\Z����Z\ږ�녁<��<��O!����Dm� ��u"v��A�yBҠ�����o:�7��)@���ǯ�]���ՎW����Y�F)c*\�G�{rF���ܳ�tikᎭ���A]�9�I
B~S3ɡ�ɦf�Ŏ�M�94`lt9�ݽ���rj���p����U����/�r��<j�6���z&rB�ʴ��2إ2^3���X@��\��a5T~W�N�쳴���(Ԛ�r*x�A�h����n��uF�-RL o�/��QBa�a_�إ=������| ���<�#����\�����)�@�ꙿYN���ڷت`a�8�7��udŠ`;7�@�8�D����%�4Z^�t�Wr���,�X6�7��W&pN] ��U�,�YL�l���r�D�泬v��8����y{�u����o�5�q^�b��"�(R�S&sn+|A	��[�:*
�2!tA��y��k��fGo�j��-W+06���$�"A�;��HM�7�(����5a��L��]�9�F�c��<�p[�^�#�욟���
�!!�"��*8HrȞ̆ags������qd��G��xնC�= yS�[c��ʔ�����A�\י�����WwU;4����� �0$R �H��#�	Ehb~�݉X�c�����vcG� eIс	Z�{o�mU�}�|f��ν'_�W�UW�P9�����ܼ���s��/���[i�Ӌ�*���f�ǂ#2��d ����K�x�P����y���y�&�s�X��V<^������B�,�[g��_�F�-n�ӿF^��L�i�ȴ��Rd1�yn�k�����=/�u{�{�׳�4��_�6�yX��1��Gν�ㅞ����Pk��gPX����&��u�I��\��Y����Y��t�
-Ǡ��H.����տ�I����mZk���su@xc/2��;{�mx�>�Q�^R��#\ꛇr�ѢZ�N^�:sf��Ӻ�`�m� r��m�C&}���S�:教-t�o}�&x�[�B߱MBК_��]������8��W���D�r�FS%�dE^���76u�>��QV�<^8�w�R�=��e��OP�ǌܽ��z%�SDb��K������/��]H���-����`CvWJ�b.����W��X;:��{IAO�_<Ɛ�<)I��}���g��p=(#</��s���'�v;��u��d���ߑZt\��/P�����]�)�*�?�O6�a����5�;˔9@w�=kyR@X1-a4���T`�=�C��$��8o�=��vS�ދlURt3�܊�x� �b�D��ɢ1�_*�|�J�g�L{�?��7���g��u�<��d���w�誖�+���t��7I_v1��U)!C� �o��e��s���A� � m�9jA��DAK�ͭUe1��s�!H��x��'݌Z2�+"W+]ܐ�tu"s��Ԇ���Ol�q5��N�h⒳�(
�@��F��)y�dB��Cz�O���Il�!�3�l�ey��U�����T����+y�vC�'/�(�� t�<��Ah���i��oDR<Bl����h�V&7��Yv����ڧJ�2����r5~_g@,��w��D�2;�>�ö<��AQV`a{ k1�#�>Y�HX{uq�J#ey��S�Qb��+�cT��)B9Oa�D�+�421I++��et�<���T`���&'�m!�Z<*8��Yk���'^n�ݑZt	��x�/uZ��8F�<ʋ��,2�n7ے��E��\�He��U�z+�#�_��ݡ�A5��@�zx�z�zսa��F(r�����8�v�����D�r-)�RR`��!���C�	�=�z>���8䳴��s������\�#pc"�?g�Ջ��O��N�~�+���Y&���Lڧ",*-F;mM^�G�1s=�Z�E�|���i���y0#W-ĭNL��2��u-W(����w��4v���F	��h�o��h�o++"356J�����hll��QY��z����#�m����vpŘ�æ�}x�[='"�@> ��E!���x��V�I�P��N]~Cc����z)���u%_�lwdS~�{>g��-�OC�'�2�s�e�4S~f��6t�?�*�����w^�������x�C�1���C��"���p:|�#�{a~�-c��L/49wO�t�[g��y���ZK�� ڎm>Oֳ�F�-%Y�r(g[pˋ��<] fζ'E<��f�r����j
1j�RaO:���_YX���q��������y�����1�OL����- 
��(��� 	�/H8�����|!�)��M�@�c+S8F���A�Ls�k	X�E��c�y{�J�
HFqޖ��%�����]�1:��:*ԍh�o���_���w���G`Dg�rۀ�ؾz��}��]�u�S�AzZ��\O����,=����舔�/`Y���Լ� s�RG����$�c�9K�tg�2x拋G�x�\�UA(�g>��+a��ϳw`�@���*����Ԅ���v����0�������I�j�*L�)�'*Vh5jIn�X��6Eh��Ԅw\�P2�|��1�j�>::"���-32���E��P67
�9�A���CYp �e��P��P-��7��4�)��^����(�y�����Z��GF��j�p8Y���5τ��C�m���&�P�yAb��%�F����"���8�Ǒn��x�ｦ��%Υ~�����zj���o	�/6��zl���)�s�g�����.l$�!��v�.<�9ˌ9@w�)C�����~�>r��E%�mX��_yMj�Q�&�= �##�����ej�j˫�櫯Kyڙg��@���ʞ���Z\�7�|��=�L����F^�+PP(KS���Q�i�?vX��J�/-����j��y�Yھ}��*#�[m�x�	ɷ�r%�s/,/�$������}��Y�6:�q eDPO�V������t��<����3t�i�I���-[��k��Fo���m���s�9���aPʷ���%��&G���g�_cˠS|�@��x҂��Zj���-��P���2�#�y���z�'�����e�u_c�:���zƞ���75�Q�Ꙗp��^�]l�^7�o.q�Yη,�lͽ�P�;˔9@w�9���6�'�z�-�� ��l����OK+˔+�i�/ ����ݻw�u�\C���M����|�a�����R]�|���}���ᔫν�@�~�)m[]l�J�[g��+.�}��PmmU���=��c��C��?�)񐛨�f���; �Ѷ����������ޡÇ��7�D���Ð�
Б�:w1D<����*/B��&�{�^|�ej3�r�)� ���O��?N�R��:=�����:�,*tBA%���=�&׈6$j�;O{�����h6Y.`eۄ�c�#/�<,�&<���B$�o!Й���W[�0���z����j���� Nȋ�~d��X��2�ؖ�I9�6��	�"�����[.��,c� �Y�!���C��Ld��mʳ犰3# �%W\*9�*���=��S�8�홿y:}����o�E�?���}����~�w�=|�~��iI�4��)�N��f���Qoы/=+���w�xN��OV��{����w��i!��hjѿ�կ
腭6���ѳ/</�~�g���c�� r?�%/�Ȟ��O<I�w>�p����H_������넗��_������>��FH�W��=���s�y$ۥ��zLڨ$�2��4|�"UjC��x�9��yQ"�#�[��0�=�y.�f��}�O�=��^���S��w��H�ރu�&\n�w���7����۪�`�q��8��aa�%o�M�l�\:_�ː�~M�ӄQ�9@w�5s��,s�u� �.��(B������f�=r�^���ܾ���z獷hnn����<2BW_w}�;ߦ{o��g�g����z�.d����N�v�!�k}�A���t���wu��˴�<GO<�5�-!�MM������ig�N��^\ HZ����'x������#���/�Їh|j��"�R@FHi�������o���;�&�|�)�喏��jw:t�UWѾ}���<>8�������n����*��@�zu��f�H�Ʀ)�	�Z�6(���F�9%�c�ߵ,�j�Ц�̇1����0{��Ƣa#�nO4ES��M�𱠉�u�[L[\߄�=��C��DI�IS��B jH�x��ƲНe��;ˠ>�Ч�`$��?��x�|_f�v�֭Ңt�=t� �x/VW����ŗ\BϽ�=��>��ܹ�>���ΞuJ`�Ю1����� ���y:u�^�R�Z�Fb`޾}��P��p��qn��gggi�Ze���Y_z饲8 �GM�:��R��?>.�y|��+��[o�%рs�=�.��bY@��	_�>�,��,--I�a�H�]�R#�5#h�P�J�L��L& �G�ɞ �%���S�.s#]�b��W��(�!M	g�1߳���o:H�}�6�鋀{�e���D��ϛ:t)[Ӧ0^���3g��� �Y���Hqx��C^/��� �;��4l����2ͳw~{�e���.��Rz��;>0_s��411IG���I:��4���?����A@+3��s��R��s����(O[�� �����a$�K(�����/��@jSb�����;L��Ev`�>�v�c���Rw�E�z�X�<��s�c�^�3�u��*��P}�R�(
� �_�e�-���}-X�m�[=mꊱ!_�z�`��I�~/`��{O�D66^�$��]0��bG�;˔9@w�5�B�/��g�`�j� @x� J 9~߱c]}�u�ٞ'2liuE����.���[^O?�t�;:'9lx�`�>z�.��"�꤫�a�i�������K/�I{�P�R6����b,-~l�\y���x�m�&^�#�<B{��+��"���i��|�;�7h�s����e����ù�����X*�`Q �����i��Yڳgv!Q*�c[�o���l�:N�n̄�����LM;u5̣�o�eՓi���mZ�=1�:���M�ԉm���~��9�8g�3��2g�ԑ�i�v#�Hc'�|2}�S�2�Ȋe���V��Mw/���d�٭3��Z�-S[E���$U��d��5�2=C�^r���'F����������mJ��XT`L*� F�������;<kx�+  dQ��`���'�|,�E	�}�8��#�}^|�E:餓$B��`a��SO	g��SO�q�����f.��{$sa�V^գ�h=�����M����������}���>{��<��G��?Q뗔=���=׵q�z�Μe��;˞�a�H�mEL
��h��.����)+�$��ۊ�*{ҍ��H����N%//$���/��Y�}�5#�+��y�k���t[P}�?�������?M;v�y�p�~����o��6#�7Ұ��g���O����%��&,�9Ǳ�cǢ�����>��/Pmu��y��	^��m_�.�,#=�3B.
�=��6��9?� 4Iw3�$"��N���<�.x��?hK�+����~��=� g�2gНeͼ�$��G& oX�� z����1��45>!�f�n���ML�n��E��n�b��|�q:��;��9^������g�����-CrUϏE<�Q�_�u����O>�$��g?��i���.�Ƙ�8��#o���O~�:p��x���|��rnl��\<��ۿ��=B��董�\��⣲��@./�v�m��ּ�K�9ɱw�ʊ3G�O�!����i�{W/>�|~/pޯ����cU�x]��6yw��3g�2��2hݧ��Nǲ���v�Y���+�ibrBr� y0�A�FF+���z���2{�&D����"?z�=��3�8��[>N�gf���<gD��2[�T��;w��P'R���5�����,���+�M��0������?����q~�9��ǎ��W^y��@��k���k�1k�'MX����9,̌vA̳]ٴ�a�o�-�˽P*��pL��5�I�lTִ:Z��.��������,�^ϓ�L$�c������u��9;As��,s� (j&��6��F����:itQk6�5;-Q�`-��P�W��<0�D�9����f_���RuuUd\��� y�"/��B^ �������2A./8�����^��1������D,�?����Z�>��/I;����#��d�r��P_�Mt�G��cb����2�cς���L8������
�ݷ-G	ѣ��lIc�������#ɌKy�DAx���D��\A^�
�9\�-�0��7y��y��d�U.����f�Է�z
�ݹ��Ѡ֫͠�q�q1)!9s�!s��,�WӚ>���3u��a���@��Q:t�0�8���Df�Ȝ��>�Mh�=�\� V��K���#e��;@lϞ�42>&,dapn	������rJ�S.��Ǳ4e��}� � ����a���:l�%mX�w <���B�Q����~�1C�3�%��'�xE����
�:�R0�A��S�4"�Q��)[g�*c����&�/����hb&)DK`2W��� �z�o���0�%m:s�%s��,k�8���k��s#�I��n�)���[o�)g�F'�j�m�;�ٻ�:�I����f40���_ �� š���-�߁�P�NL'�9Yu6�ܠ\��6�.=ɩK���*���S�ց�����K���AÛŶ��9[����	ُ��q��3�?��X?��d4�Kj���z�)�D0�A���g��K�U�k���P�7
t��gfw�j���+I� �,8��l�ըt�Ü֫uz�9�5���h��"�?G��Ʈ{�Μe��;˚1&D�C~L@	�,��,㲫>Lw��G��|�^~�5����C�LR�(ߊ�n��0������	ڽ�$ڽs]y�et�����HSr�`�o�o���˶�5KȊ�r�w����C�1��#g_o�7t`���(�[��k<�� ~���Bjw�]�=�g��J�C۰�Q;�P�3�&�dv�v���Ͼ�}��w��O<�s���ұy�,�cvMm�B�>�h��|����G+�4;�����j���|��f˲@A� �Z��l�~������(W�a������2�9ˈ9@w�9�"/q�V:�V���VC�����;��׿�-������5ɫ��mW�Ҟ���8������\����?@͕5*20~��[���_�w��2)��c4:�^j���x��A����������g�:�G}T�� v0�gff��>�6t ��u�]���g�!�X�  X��?�r5��#�ܽ�Ά�_:_�0�S���̷�Ԓ���{���w���?���@�__�簘��}\�y��D/�~�D!�����
Ԭ��Pu��8����R�������{���/��[Ϣ*o�A����f��3���F�βeНe���eAJrB~�2=A��?��?��d��f��ZԠȏ��(��R>�֗������s��*�^�A�=���)����
p�����b��- ;66!�aԑ�w]hh~_�7�Qb���?O��O�$�uԡ�3�7D�����&������W_0s�q�^����\B�P�CI����|EHyP�CiJ����K��wozb��i��B�v���7�(�1h��Ez�������[�:i��^�0�7b߈򅲄ݥ��A��/I�`:���r��W�E� ��͗^�?����������O=<u?�7B�ƙ"y�b �@�y�\��Y�����yj
��<�'����OP�������z��"՚1�{�b'�%�}}�^�>�m f�?t��B;&�iˎY��wы/�$������M��-��c�-h��N�����2�}��'�O|�Ic���r�-���_T� �_��0;�������#�ZB�h�
�4��9�gnL�^�uzΒ�KH��.`�|�x죓t��'���#4}�NZi��IT�)�)�x1��>6
�`���
��:�Gh1Oe޶�\��cK�����履��s��㟠7^yմ-��6[Z���٬RܰqE��rw�=s��,����4k��!˄�s�������4P	=����*%�r�y%�.I�\4Ul��$�C���R(Pci���@�hz�,��i~i��9�\�?:g��G�a�<����;<\m#׍P9���/�8բ�g���/~�T�;�X��ǎ�!�<;z�Ð�Ƕ8'��ct�y�\�b(^
�ksH�ƶ�w�z�h����T�EZ��y }��AGT��|`�!�%
�r�xaSy�,�٪֨�\%/��(_w+�
ߧ��e���ʈa�N}�
�}Ρ�WK�ը��`���3g��;˜�>�,oC=R��B% ɨ�{���:3A�fK�Gi�����O���Y�q7a8�#9~��^v�����r������R8���&ƥ��HP��ؠ�Xh�c�5*��	��`�⛒�������,W��@�`A���ⵣ�*t�u�@�WHłD�w���l5�_��Dݩ����� H�i�O�	R�)��i�� �F��ŲD0P�Nh[�$��,^�
0�a�x�趆F�r�B�L��*UFG�_kKu�e�\��s�ruP��%`&�'����I��H��[g�yO_���K�~��J�"�C�Cw�5s��,k�G*����އ���}�؛�13K��1Z<|�ƶOQ��B��&
�`�h$��G�U$������1C��4���8 XȾ"�ݬ���xdY�A��ũ�i�R��/ ��/K��8����:~Cx���/�;Y�#�]��h���� �ժ�0 ߞ_s�:k����RiVX�6i�L��Z�����?z}�����Brõ6�VOŋ#Y\T�%^�<'�8�~�9�D-�xS)V�z�֪˭����BI�t��H�'������r'܇����Ay��Cw�Es��,k��e�ҽ���Ko��a~����w��[��|�/��k����$�������@<`����\����w� T�5h"W��s4]����wRk�ڨ&����!�ŉw��Q/ �a_�Bݾ뤤�֥k��Nj m�r��8����=р�`2�thԂ0~��L΅K�G'��~/8)����B>'����V���;�w��[�����v�����w��B>`�����z$Q� �慖�_�;���hP��������l����c�1��;] a�K"76��`���Нe��;˜EQ�
װ�x썐֎�Зo��<����As˒���T�T*X遭gO2D�׋%�\b`Yd`�����t�ŗ���o�-]p�Y4w�S!/H�^g��i'�r^@�<M����X �"ﺲB���~� u�7����ַ��r�Ç��{��sGKV, dXL�����2���\���
�ݦ*��vX��0R��E��t�Fxt��!���������5z���h˶-dtۉ�~��GW�����EYa�� ���h�ʹ�i�N��#������g�.�?� ����8u�Q*����U�'��ü�_�Y�;G�s�)s��,s�y�:����_�z���2�]�/~�v�����Cs�i���H�c, �3�h�a/�J�޾S�PZ��<��{B��S�tl�K1����a��n�g�y�������w�QK���oK��ݻw�g��jx�`�?0��9��ak?�@�&"+�������ې�;F���X�S�ޢ"��6�Ѣ��st�%��/���-�j�*�D�B�cD���U��D宔g@GS�"��y�rln��k416�ǩ`��K�{���������9˔9@w�=�"��\'U�g ���Z�hI�U�֐2�]�[�]{��*r綵hD�=L�z�bާ��Hӑ�C�R��^A�@7�YFvZ�솀ՃT�V���=��#yq�~��j��`�#���k�� 9�e�3G�9�?�я�?��!�1��vکt����9���N�0OV��M�l'�E�!_�5Uc�Ja�CͨC�o���Bwh�ĸ�ec��ۈ�ow">F�ڢ:o��E����|�ɱ	��������^�S��OWpO�]��{-�s�,�� �Y�̋���~L��al���'�-��֨5��sT.���l��@�i�b���nIwph��ث،�F��ˬ�>���x��a�����<�rGm��}���q���� 	�2��ؑ߾}���߾}�$���M7�$ �c�z�P�MMMl�d�����=p�/�W*���.�XB
v|j�-F{��@���~��|@�^Mw:�yl�S��(�)�b351!���[f$Z���wx�����M��9��	c�oi@�h��;Pw��gs��,s��qB�TΔ|&���HY��
�ݖ*�ZC;�Qi�:�3 G�a ����P�V�n4�=_r�%�]-M��\��|�69M��??��� gͩ�{�v��O�ԱZ��q,0�N��eT-��[�g��tsn������kC�J��B	㜙�yX)����x�O�L�@D�8ՊI3��;���ZsM�TC+��bf��-Lע�ǭ���yY�3�
",�6�j���s�Y�e��;˚yrOٛ����Bɋ#��kS�T��X,��8������Qzz�@��BEB��*�l0>�&�N �PڊJh��y�T�5�u�&���J̵�\z���W�Dj���ⷖ�.�|-ڴ����'� ��!z`gL��8Գ���D4�:�r�kGIw
��s�4'�9�1i��+��^rd���Hz��'�<��Ӵ���N�-JyP����w��8�ع��;e���:O>��(�AuO�J����F��侭��{C��^��<ۃ>�#r�,k� �Ym�b�x�@�6�6�J
�/�8�d1Ru2�lsU��x)o��@I=�h&��+!�rEB�0 @u� tU�S����x_��Q������;H�r����u�7ki�|�;M�>�^�o���}���Ԥ��yL}��*���������s�5�~�C�=����	� v%�a>x��~ɇ>D��}��@����@��M�gß�|�	�8s�us��,{��~���CY ��E�~����!S��B*qj�֤��lk�w�� �����{���Pζ�pL���tW58Ճ�׺g�9��E �� 9�"���\�^���=HN]Z�xf���\A:m�������aj1��Ez�OLOѡ#���e0�I�b����*zꩧ�{���r��N�B5� ��	�v�<��kW9\Kd����G��O����d����>���@�Y����̙�J��w�a���hn9��
������p��F��K���]@`c������l����+���06���$`ᅞr�)vM#Ԯ ���n�t���Y����^���ը�u�o�Z�H�"-��)��I� ����D�v��g�����|hts��C%}�nǜ���f|���=�6�ѝ������ޙ��~����?ν�%L��^ڼK���Q��S��F�����?x`N�Ȼ�k�o��G�1+�MX���>(`t��W�t�m3 �� �đg���/�w�!^*�A�^�Vr~�����<��3�Y�߷0H����5�P�FRW��h�"|�F�@b��G��fffe��rE s���"�\��v��C�mf�����PͽS�{?�u]ș��tgٳh=�}�	aI���9�K4{��՛��$��4�L&��~�dC���p�-�~o�1"8vxېo����mCl���ܜ���C+�h�D������~뭷ұcǨT.&%j+`���8�ʌ��.O�����s�*�I�����m���h��7�25�`c��+Z���1(��c髞��� Pđ�m���b�βgНe���U���g=��h��b=�
���v܏|C�ħ�9���{=y�!g���ƒaJt{������җ�$`�����K/=��|�Ft :>�3�g :f ���v�����W���-�F-aҿoާgcJ\wH_Q��'�'cHnA"�Ӗ����5�����^��{�f�l`~����G{����7��ۗ_~Y��k����??ɕ�7���A��9JC4���49�8g4�βg�gG� �R*�4�]ּ�o� �:�ܮ���
� ��|1��_������O?���饗^��;_<t����D��_|Q�_1>x� �j����A���6c�˧�U��K>�������R2Cq�n�Dh&0!t�_�,/,&�6p�����h�A����8�Y� ��:�!'���vi⛪߽!��I�ɷ��5g�2�βf^E��O;!{x���Д$��9�s<��I���m�N��� <�cK���Ep%\y~��@��?P?�,i��r����� �ԉ�&��m�9qM{���b�y�1:c�496) ������
��/~Ir����c�ѿ�׿/�����7�p���ri=s�l���+�}Ƕ�Mx�`�{�sh`'9�H���.��y��s��/N7U��&�\��u�DJ���1���q�:��%G��k����g�{� �G�Ǩ��o�O������hA_xhܯ,-�������{��� r�����p�F�qfJx��w�0�==v�yo���6v�,#� �Y�,�b-'Pּ�
��3�C�����b��I 0xs��'&���-m2�2C���8 yk�x�5"���*ߊ�7Lz}�S�eQOG\��o�Yƀ��3���+��'}X�������΢����?���
��2���� �=����N[�7*L�!�������H�o�c�u@�vp �;�<?�y��_�n��I��Ԏ�D( ��Dw��w��d|�;0�L�A9w�4r�8g�2�βf(|�%�����{Ł��&
h����!�]�޹��!ԫ!Y-kR�qӑ�g�����y�U�k��T4���@v�����RL8c@Q�ux��ÎWx�-' ��h���s������ְc���P�B�� �O7�a�������@���e�7�F\��\���m�����k����:΁�u8��p��?�� ~.������Q��>���Bϙ���tg��Xj��g�GW� �-W0V�� � U���І׮�=  ���
�$�:~��]�U��)ʖN��O����0����.(T8���Ɓm)�4�?��O4�����A��	��'���r��0����	��8t萴����� �S�R��yp 7j�a���7�:�[&�仯}��e�����je_?HK7�I���B��2eНeͼ8���n��&��%�or� Z�EX������5B�x�m��Z��x�	s�J��x�)j��@_�e-�	�<p���F�=<B(��a
���n�)y�8x��Ǆ����!7FXy�g��Q������~&�q o��|�����k����L���e��T��u�'�6����q]W��Q��2E���ɼ���_�!�Կ�կ�O�Sz�g貋/�������������i줨�~����}s���Y�����Y�efi_�NǨ~XQ���WۀE�6��D��+�H��.�^H�b{�9HV(�¾�`�~��O�ϨwƹP3���L(L����+2^5�� h0��	�=�����>�Lr�����N9~�w�;��;��������!��潠�^ӽߛ��v-�+����sa!�mP1f�5#�7�i���sϓ����W_%���s��p�7�O�c|�,��s�L����Y�,]ڜ���t��V�� �ݻw��P.´ I '��\s��`G_q�<a��A��[��sǎ]t�E���Ͽ���<N�7�|[ itt�=�J�2�H�h_��ŃCϫ��|�S� 7�p=}��ߦ���o������w�+9��/���k���O�D�Է�r�D#������ҋ�����N&���?Qt��E�0���V��� ;�)�o@[�`a���z����������#2���k�	ٷ;!}�6�A��ŽM�9ˀ9@w�9�ZʴmhR��&=��R�0C�L���� ���6��GoWs�
�"j��xh#�o��bj�6����)�j8<l����o�]B�_��E��g�8�����b ��/Y�W������C)���Ajh:w�ޟ�#�m�����׆{�9��q/0�k�F�^Q0��Xü�Tw�r�!��{v�i���bw���;N����tg����nX���n{]�P�l5貳/@�G$�R0 J��{�0"�y\ "@#�����3��? -� X ���.W�,9�c�o�)�C���I�Q����V��c���(���O|"!������>������G�UL�EQ*쮞p��DK�6u/�'���1���}@N}��IqL�}��.6D�9;p�m���yY[Y�{��]�J��/��{ӛZ*��1,�((H�nn<o���3g��� �Y�+�iB�-�[���!��:<��y#��4:�ၮ�8���_��!����\ �x��%��}��,�����B7fv�M��E��	x��=����a�i-q3=��B���;Ht >\;����a��Ø��B�x�y�5\�FF�p�!�T�5�{�Z����u�z��B��n�{l^jյ����/l63�a�M���q�1s��,�&�t�I����/5��0���?"�c�6:�ܳ%0F�zϞݢH�%c ��}�3�����s��^)2��kk�S��Kl��1����E�.p�����:Ή���A4	۾��o�_ȫ#��c`��у�+~GD%��ց�p����#=?��d3���L\7"#;�ip���u�|ڐ��P(&u���`�{s�w
yq�i��<��%�OP�֡kj�i�<�R��9��S��մ�9��;˚9@w�5cw+� 檅n�聼�+�ÿ�h&�x�c[  >Ã�þc�Z�mT�Ek�� (��P@�<Lu��8Ή X��#�\7ƦHv���jh�?�Խ�?F�@;��r���qz��&�/�0��Ȼ�1�H�*�a{�ٱp@� ���,X>��7��<�\�� q��s�P��j�����ۻ��ȋ9��m�9R��L�tg�%<H�~����=���:{��bcɑ����ku l������o�� Y@����YRx�c�f{zj������"K���;o�.i�f]t�G��e ���"���>Ʀ �d>	O�5���F�����w+J�^�`nq_>�������߉Zޮۅ�E��k��F����k׈˧>}��:*�����v�k�]=u%T����Ͻ�~��;s�~�tg�3๾W��e�S!�*�Z���|�KHV�r�s�0�ޕԦ �R��ѫG+D+� Ӡٯ��/Ueg�t�i{��rn���Ņ�������0�� rc�	�~����]���z��t�p��j����@n��=4.�������0G��"^�aA����c"0�?�(@:�~���'�m��{.��,s� �Y��PVE6<��Pm�FB5���W�o�?_�}~
�x�c;�DW�x���D������Q��N ��ϟ�R��H9)���@GY��8�	J�4������䚰 �z� 	���͠EFB���$��m�oC�@�?����rσH�Z!e4���o�guy)��žX��~�	�o=�}39��M^�9��������R��x� �B�D� �o��* �Q"�}��~Z���oeE�;�Np����\ >��L�y#��rV2��X���`��3��qk�T =�����w��R�(cO�$����uIq�Y���t�������j����U^��^:�r�_�^���3��K�<���?���� o}���=�uy��Νe��;˘M@���+6�Y���F�x�b�@��`�<��?ԟ{�y(��7�6h�	�4@p��d�[o\<����ރ<E��te��B�v�J��qڙ�$�.� �5m�װ��`J�>?C,!���~R��cU�VAY�������nё���}d�`s��.�!wa���E�@���{�kP@�<W���~��_
cA�܀�o��Z�!�E�M��~���&�W_72��-[�E����cV[����rv��^�F5z98��Cw�5s��,k懱����J���i������"Tr�%����ߐj�4!�
mw��P&2~�Z$D�;9r�0����x���9�k��7�wKS�%l𾡌��j�8]��g�;#�6�z��(�{U�m71�a^�f8�O^�:��>[X��΃>(�8��&0��5\"�q5r�l���F^�mn35��a�EΜe��;˘U�COғ�d��5T�裏J9@0b�:�^������4}��w�M7�,��F �|��8�LQf��~@u��������������k�;��T��q#�,`�{���G���q}P�;�����Բ9�*[����ǐ&��e��{�Я7Ȏ��?�%)�xQ�9"�?"�^��$U�~Z>c�ṃ? ���J�����a ���U�_=������A�>o��Qg�2cНe΢TQ�A ��C�o Cx� �B�$@��9��J%è.�M���I��7�n4������-�!���h�w%SHO�6�Z*��ZX� ��b�Z���EELu\*3,�-�1t%#o�B`���n=]\��ϵ@־�Ǖ�(�1�/�V9��q���ת�r�sWҡD.�H�KsލmB-Ι�̘tgٳ��*�` 1
�7�����+�y��S鬳Ρ�v�,�9<'=�WW֨X�Su�&9�Ņe�<ő'࿴�"��JŲh�cq��;@�5�ǳ�����u���qhVa ���38!/@�2�z�i-yτ܇ע��a'"��~ƪ*p�:�B	�~�K��+;ax,�00�Ȥ	��]�h�޽{eۀ4��ՅL�|/�w��k��ّ�Нe��;˚yq'�����p��:�p����o
��A���e���ڐ(�������){�����h� W��r\4?�CK�Y���[�A�!�l5��Y䃾W@�>9��h���`��Ǉ)�MC��O�?w@�ʵ�L�xl���Y�*��ty3�(�5���^W|�b��Λo�)�AE��7i%j��g�={�Z�>h����3g2��2g t&}��Ј~�g���W^u�����>>1J�_q��qw��FK�t��o��K������#����J��Z]���6ab0�G��k��5��a�A�ђ5�^���4r!����>&�����fIq�������*����\"��7H���9P�g�=R�v���7���^{��G�]����Z*��I.^9�?8�k;��s�4r�,C� �Y��C�y���J�*�
�� �0@tO���ࣣ|H�V�5?(���=�A�B���=�L��r�J5��)����Ѣ ��bE��>��~����Gq4\�����$:��xw#��S/�o�4��׈�1� i���g?KO?�� ;�ª��9r� �[�~�`�����~�5�$u�:��~��:�_{�;vJq�2gНe�<��AZ|E[k�0I��<���H�L�+KT[]��I���₈��������G�E�����"ML�X㍣['!�aQ�j!?�'��K�x�H���ܵ����),���z�J���wewk8Y�^�{�������dA.�&������/6*Y�/�Kk��XLZFץr� b4��+B�JpS%8=o�J��;D1��-���j�]ǧ�����r�T�a�`�za!���[(8s�A�tgٲZ�ף޲��>�[��%��	[�ru�Ⱦ�n���y�C2�uraS$�@ �K'6-�R��blR��0����2��d鴖|�*��i�.b0~  ��t��W,z��~K����)ŝAl#b��j�Cs�0�����~���	�A4�-�@�s���o�@J� ʩ$�.,�_��[��t���ϟݠ'��q>OΜe��;˜�q� j�\|���>�G%��CJ�k@��G=F� S��k_۔�3Ҥ�T
ǚ���m5��ƫ� ��Dn\Ρ]��;Us�. J:.#[L�W[;�a� W���&4ͺ��.�
���o*l����z���|�&̋F0�����2*ZjB��"LC��*���� �^H�*������7j�溣��N����"�;˜9@w�-�CG<�<��{UO@	�5d���|��NI��+�J[U��
�h�T��h�6��~�2)�kq ��U�E��ņU�q l�;�F���f#��|b|R����c<0�ɮ�:0ѯ�����I�����/�(��{�y¼i�D��B�@@&=��x���I#!�8�p:[YQ�@:��i���;�ߕ:���.��,[� �Y֌��q��`S��b<� ��۶��x��;���
�sGM�/�)�R��N^�= ˥
���;�ƛ#z����]�4���O=#�$΁P����p���,�c�B �Cn�S������=divF�p�	[�9�#ߡ��'�z <�ľP{���~��5�a��\c�p͚�{�>mU��Q����[Cp�
���"��i��'�?-uS�����0�F�5(t��Y���������5��� _5���U���h�M7�$���}O�x�C���K/��,���|��e�"O�4@R�(����k陧��5��6����b�ȑ#R3~���x��~�e�ё��е�'�S�2����s���1�ǎ��4'���ya���C)������/���3�k}�$z��0
ri�}>���h��Y��������>��G�=T��Kǽo �� ��b�P�u�C�s���
���HH�bFy�7�7�ae�i3�v�\��~�*�9� ���l��ɳV?*#~ AuiE��np{����Š��o�����}��x�	�.��DI�m;�k���ꦣ��7-��)i����>ˠ>����F�ڟ�/^���c���dL e�S*��w�R�s�;�~�����U��1,�ԅ} �?��O����XƊ�do��p?���A��9����o��s�Z_z�e�j�u<��Sr?�j�����oX4�����T��n�p�~��r��F���{N�_vI���'����J�6��6G�}��|9s�A�tg4a+�;����xb�^y��b��^�}{O�� < �i��˾�= y���D "Sƅ�: D�x�~�^"��m 08��\t����k�H�K.�Q����C<F�o��������sΦg�z�J#�q�.Z��Q'�h�����$�G�h��k��B��UE�4m�u�
����m�������6���+����cQ��Ƕ����������E]$ ���x�PT�w�Ek�d`14:6BG����8H�����$�b�'\�!��~��f�Z�r'ל�Y����lY�A�3b<����VeK#4wl�r�"���z��g���}�ctֹgѭ��*@p�]wѾ3�B�#�#�ӏ��> ܓ��.rPC�:�>��mߵ�λ��V�eZ� }�g?KO<�� ���(��B�K�����t�YgS�ǘc�y��'�_�O~��459-a�N;�xDP�>��sdqrٕWP��Q��}�i�聇�[n���@?��Oi�I;y�c�Cˈ��!��[�vo�n�vDǞ<�X�8�[��I�x'
�ch��Se|!_g�ա='�,�����I��3Ζ��[�����yQrd~.ɕy~~�Q	�_���1Z\Y�4�_}ݵ�[��f�9�����Z%�V�."��6��łɾ��u n=Q�[��%չ$���tgY3�>���Δ�~�ɻ�ͷߒ0-�4�]��'�m���<a����CV�����!`.D9��n��=��C��^8@��\ ����~����'���<r����4=9%�xx�XL��G'5����	�ر#a�+���-�_��ʆG����O#e�|��;e��������]��޳�a�q$9��bJ:S�?�YU�p�Pg��9�ø�q��`��x�O�,1�{�^=�O%]�Y:�;Ҝ%����z�8�O�X_��ѹ��y��="���Y�����k�� H�<��A�uvVr௽�������Gr�BX"T���4k�9�������m��g`9��y'g$_@ �s���vmeU�ğ|�I\orr�=�1�x��ˋt��=46R���3�8X^\�r�(��@-�Fxa�^,����"���[���Syt����{�9t�i��x&&�%�,`f{�A�J�:Q{��� f{����#�شp���$��)�����PX�1 ?��C<�;e����j���4[����5�����~�>3+cFU��H���9���΅!�N�%�5&;0w�9s��,k��sIs���F�&�p�򊄥�&G޵٨����1����c�2���i�T����@_35�h�^& �����c)Q��4��6�F=G��=ƌ�@���!��q.�.�vv� ߵ��Q�$<�mTTE�j�x� ))�ʏ���ވԶ��ӯ��)��p�w�!��P)Z��GdB�~�h��Tf�V����I�|3׸QyZ?�oqə��tg�6x�Fڕ=���z#��V[��E*���@Y�̵|@�~㘪�N��6Z5*�Mw.�B��@������F��;!�۵D�u�=���1j��v����/XaÈ����QZ]Z�|�(�^�B,�L�]ZδiA��Zaƿ���b#��,{�a�𤟸�=Tu:x�X�D��XC(�S�!�iyy1i,`JŮV?�� B�#��>6:b�=
)��v�-^���-ds�����]ﻜ���ű�;˚9@w�1�� ��?��o�ht�t&r�͖ -�w����!܎�@ZX$�e):��EKkR���WC\sݪ�:�&z m�|�1�{���*��*t�O�ِc� ��c�-���i����w�z-i;���*���9)�?A�<ٍ�������;����?��@;�5Xt{����:U�+�ڧ�Ss�m�:ȥ^}��]ZtG����y�;˜9@w�IӇ'Z����,ȥ9�!L����-�[6^��-S�ƃ�^��[��M�w@hZ}wi�rV*T��>�ײ�]��!|�{�>�����&��+P�I��s|�	�Ӗ��Y��ԭWUa��x=����C�|����NkSs�}U�w۠��R�B׽������P����p:J�p�+��T����֫ܫV8�ek�6*��Ez�T�G���r1����sWw��s��,{�u]���1��%��-y����x5��Ji�OS]��z�f�G�p��'	�Q �}��
����3~��f�'ji)�6��+!,�J�u��{Ӳ�a�����ԓ�(���Iq'�S��>iiXo73�u"������ȨDU��Ke���Ru�������9��{�r�e�;�6�=��h���9s�%s��,kf�XS.x�Zo=�!��6:�y�Ũ>|��4�k�QR�$]�x���a�x{%�SCp�U�2����8W�x|��{�i 5��������M, yd��.v;� d\�U�`�ʶ谓�����ߓP~�Ք��e�8;�r3�r<탮i]�D�^�yq�Q�j�ӎz�q"�C�\���S�CwEj�|�����os+c[��{��)|@|;���c����x�yé�M�o}ު�լ0�V'L4�������BDP�,.4�m�{��md���(OӅ�.0L_wl�w��,S� �Y�8��(� L��y�:am��r��e���GMh�a�K�{lȃ=��ρ��lM�9��;d��r���c@ġ=��ݺe���x ���"�$}U��m���.>l�d�X7Nk�ۨ�F�����zˋ(���\n$!�I>(��f��S-�+_��n��K�/�	��@vS��'�x�ń-g�G�cj��Br������UU�-�������J膺X��<Y��0")��U���Bl��c�/���t�uל6��#ˣ��Qī����9�u�tgٲ:Q!��፛���
��:����3 �6�g��̔0m$�v��M54l
�l�!@�X^<�6ګ�\YDl (Ǖ�C��<�z���  D��� *@�D��;쑓��)�=/����B���ī�t��6���
�� x� .D��;r�⨔��ls�@������J��|�Kܳs�54^)�ƾ�h#/n��yiF����b0Pݖ���U�i�UyE�^>�?� ������	�.�B���>d(!N���U�&>�~q,wg�2�βe1�nq��n�X�2��B6y�^*,�%}eC����,���s �[��,gu�����\���A��F9B��|�Nw!�&�:J� �6ߝ��91�㞑�PS �v�J��\;t�s&�!a�S')�3d�v:O�t�Ї0ÒMM{�x�xo�=�!�)��l�Y��h��\_L+:��U���"&hjj$L*$���޻���T����F��G�&a��.Eme5�!� d� O����]�U������������{���9}���,�� �Y��Ra�<C 1`��ԦA`�Y�!����-Lû��C� �g�	�P��P��Q_K�����Y�sM�s6��ώN@M-0�x8�	��~�c�5�/��3�������P�X��1j�%\���30�)�ɡ~Ξ�K"X���l�ÇK��Хr �N}`)`o�L��v	�k5�S�]�*#S�E*B�K@؎O�lXj��L��Rw���@�EI�=fr��.*,�ba"������Qɇ��� ����{�)����7������ޕc`a9{=z�0����(�8s��tg���ju���U�_\<&�0��  �����g��T��xvE�� �����<�"��h�\aO��4k������w(�	0[B���v�ir� �,��%�y����i���0��u�͆Y�����O��HG���R�J^|	�wх����P�+'ҩ��%`���2뽮�:��_ g���|�]Y���)��U,��bh�6�P�l���P�B�K��A���u�m`
|��Ցk�H	oS�
p&*�i��ck���s{��{�P�:mI�Ș��b'6U:kuj�uC�Ҳȟ/WW%Ͱ��H�����jJ�^_����ͫ%��U5��[�;s��fНe��Vayyijk ��٭"�	P�b��VȄ?G�'��ǻ���O�Łx��a#?�fi>n��=������$�;5- ���7陆.��<�rU�P��Zd^sAR�&��oI)�ޭ>{�=i0���ء#�ů,-
��"&��
HfE<���B�]/Ҽ���kt���"Y���vʛ�1��t�m��e��a[�ړb! e> ��b�.��9e����%��\,��A�OB��fҌE�p�ب��"?*�����^v�S��;���29e���@r輀(��4^^t�ZZ"I��.��K�g��ޭj��Нe��;˔�J�ptt��t���sV:��:�0�@o��}�2� ���6�/RQ\0�:��7M��\�8�1����D��~�>ш�c�������t饗R������� �o�p�h|bTR  Ǒ�1.x��OLOɘ��L0����� �P7��wQ��A�=�q���ϐ��J��x<{�yѐ)�X�^�#�
�t�s�Q%���d.t z��L���$�td�R�d���Z���//�t��:@sG���*�/װ����,�{�7�6����=U�^q�?�nܯW_}U�n���4=9!�����X�IiƸ�����7xn&�\Q�\��۱c_OE����6x��ꫯ��^��O�Pz�u5/i��]��&)�5��H8�,�zk��nIŅr���J�8s�s��,k�+#mSo�I����
傂���4��x��+	Q�mj�����!�G�(�Vimm��*��!�JB�k���0��!�`dK�"�TW��W�}�U�3�5Q`��؂ ��k�YX=�b_|�����5ّ��Ls��)�mF>����qTFGȟ������>��`�gZVX�2��J��$.f&r�F���({�kU�U���_a =&��cP5e�hXB�:�����@Go#�]�ѩ1z�����˯�W�Q�
_�O";�j�ŞDB��W> Z��$Yox:��s7��|�~_8 Ddǅ��z����j8V�����A��[៎�o�H+(1�<jߧ&�ڏ�5-�jȢJ瀒P���<H���/�X:��G��-�"�;˖9@w�1���!���Y������Fs�5�z���4>V��/�Dw~�����Q%U>o����Qt0cOy���6����lX>HylRwM�5��'�˲VA!My�e��<@3���F����!X��;z�#���P���t`q�����1���c!�a<9ɝ�Uz˯4ԍ�,r�h��NJ�E�_���`�뀂�3e�FT���-3tΖ�T`ﶄ��{��G0�d��BP�Y`��+��xx�W�򱘈Q��4��gD@�9|/"/<ǝ����-�]�j�}B^��F�'��s���|�>�o~�ր��g/��'����+�2UY\�Y������W�r��t>��pM5��d/���T��c4�`��������B<�S���xƃ?��~d���#�-S<�{�����G,�F\�iE��n#a��Gj�n�p@���'��7k$=tzc(����`/x��d��-�Ջ�OZ�]u�M�[��?Hq��U� WJ ��`��_�`��8Q]>Z(�D���S���?/�(�X����x����o�[��M4�p�M��l��{�}%S�G�����oG澘?��	 =�/�_��s�\���e�Ieަ�������]-�(���2ܝ��,S� �Y�M�"�aq������KRf�B_r���3��p���d���x@#qGj�!&V 0�c�0(�����S[�D�����f���yj'x���m=x?�ś�ơQ��;O�[<�,�,��qѣf�A�F]�2R*�8��;�\������ACiM�4��ш!��������/*�R�t{dB�^�C�$k�B�Ћ�/:"e����c)�$,��Y$��/����%�li���Q���-���LD&�Y'P�_$�������|���n[f��3 4��"&�P�֨�s2�+P-n���j'�?�7ǽ�8hQ��YV���LY���ϰ�ӍZ`�`�@j-u'l�?����nU�T�of.� ��=�^-c`��D�:��X�Q�H�&�M�=S�[��x�N^n����|��v����,��&*u�޶�@�c[��tmڃ��~ Bηٴ޹��62:N�/�L�BܺW�Ô��o� ����yL�+�J�ն�pr�f?߲��Y,:�6t ��V��� s �k�7�s	��U���q����ܿ��-���P:�UFǄ4WC�}u�(�r�D�<������yM�Y��Z���Нe��;˚��� ��A^Q���� ��|.��*�Ŷ��?�!��i4�0
��_d�������|�6 Q�O��6�c����)�w��	��'�k����g+L�"��(�I���3^)�l����cl&O��G�U�+_r�A��N/�u����j�k�kؾ��H���'����-|b��͛<zlJ�����Em�PB&Z��@"$c0�>��&�@*��g ��o#��i(ҺZ��[�۷�j?Vn��&��-�͉;�1Q{#�k� ��Ƌ�[/��H�@��*�GG����Fz�]�KŤ��Y��;ˠ9@w�9�S�)Ӟ��R��F��햰���.xa �����W�L~\��Ȕ��IJ� aw����]�P[�9z�?�I�ۂHl�~�~R���;��
���B2�N:t�h晅�����v��D:62�wTD�A�&s�Pv,��"s�a�iw2�#̞Σ�mi4� �%Z`4��pMd��QvF\)���#G%~��4�a�5���E��໺�Z'N4Ye?�^�/}�{Z�i��ld�p�=��q���Ev�<6N��Y�<t���oclf-4þpz�땧Iq��	�9ˎ9@w�9��ܤaaP}�h�(�0�E*��Jc����:�[|ū�S�n���t:3aT�T Ȓ�L��ԝS�~�%�y�<�D|����P��0u�ѢB�$�g{� 䄱���>�҄�Mr+�v"�?�����vl�U]�� F����L�B��;]���*0�kHK�J��eo���c��HF�Q¢Q��H]^���&$��3c���|6����%�)�ܷ~��<l���3�t��9�^�����B�NK+�4���NT-�3�.�;�Wg�3��2evss�\�*c0e�{֫�)hIx*a�P���ad4�� o��@�ė���;x0�M��v(K��� S�y�و�-Y.�����R6�8q�@&��^���Q(��y
r�~$���HS��0m�&?�@���#M��f��n��cɟ�P��+�tx�F��z��!�a
�a�v ��oEm�0H�������GM�'}�}� '6Z I�;�,b|Y<ج�g ��c�]{e[����RUk�};{�s�t�ۦm�I�X�(��Ȳ�DQA�E(AB ����|�o��$\>��p%D����v��n�s����e�UU���3ƘsV�}����W�UU������g<#�V��m�x�'Vk�nY���[���SO��rnP��=$���� �ɍ�<l�v�*�I˝j�c�p�j�]����ڥY&�����nE�33N��uK�;�_c�cU��}9�F�N斋��:oe���d.�m��V�e�5��Q1�o���Lȥ�oDYW�7&��۫�F����ԹQ'Ɖha���� �~�N6�pk�G��y^t��6>�T�W#k]�i�-��;�	\��k�2�MP�=���gc89'��O�"n#9�8�����1��\C�������)S�Ž�L>C��PV�T�'<{�|GZff~;2��?�:�cM��vq��j�f�~^n��y� }�	��zR�2�4�n啾 #dD�{G;���MjsZ[��.d'e��u�&�1�����`c3>�T���	|N�o��N�'G3�� �Q{��k�6���I�"�X4��\':%vlj� ��z �`Js��������
���rv���!/f��sB����2[��z	'���>ǒDu
�GN!��:���'d�k	��me��5���ʾO=��׏J�g�y�e��N���\m�K��W�4c����>#"����6)�M�t����fM R�Fq�����
.���Jϖ<�c$�����QىpӉ�/�;{�w�j���v�*��|؉_����V�z�����:�sW���?Yh�������x�g�#m���}���c�(�Y�R��E/�xn�H�'�i���}�D�a���E�`5T���&|��i�We���}
��U?L�����;O�/�Fk�����
�]��#���v�'Mt��Ҁ�cT��p�g�[ 9ZWvtҖ�o���ϞFgu�lD0�P���?�����}ދ蒕�`)x�uPQ�:ku9.�ʾB����d�L�mk<��ۡ�.6=M�Е�H��&�R�C�ueJՊ:;Asp�C���W>fM}ס�Kx������:X/��;+�ݜ����Soy�s�	z�yS�`J�O|��h���ZZQ�w
�2;�l�N����	v����:NE���l����{Xk�]����ڥY(����jïE��C������mWH+S;O1��-��Z����(1�޸L�1��D�q�s/r����9v隭�+���F����c�4]�>y(�!��0�]�<��Y���D�xeV� 3D潉׸�-���p\6����w U�C�]Ep"�P¨]�S�9�7��۵ �ѧ �Sõ��˜N���|�B��<�@�I�,����;�(>4���O?.�~/�1N���>���������څ�
�]��aԤ��L�j�˛��֒h_6�3��D��7[�v�m8���n���jd�g������=S)1u���&�2����Mq"vΕ�	4eE�Z�څ�^�����+�'���d	~h>4�ۧ4���|\�&Ϲ��.+-��D�Y�wP���M�F� 8��=#�Qv���фe�L<ճ'�.�)kA����
��8w@����w���H�Ep�|��ءQU8�y��r��K���	\����b^�AXm���W�0�, ��HIh9Cڣ�r�GTX��4�V�Pnѽ(K<k�;g_G��֌ؓ2�(pb=ݮq�D8NT��c�t���tx-މoK��}Ј��2Zղn��c���A����d���༕���5f����@-��3���N�Ċ	�,I|����$Af>��a������5K�¨ml�X$��NO�q���`=�COY���� �Dla�eB��-�dM�A����s��G�>�CT'�������T��N[٪jf��y5b%ŭvi��jfmj�:��p�,�$�z3�J�of���b�f����4W[�{	���a��?���F��O�;��hmj�(u�vmD*�����O��]��Jԇ�~��+����;��5oo��P�G9 lKH�#�IP�CmQgד��Q��8µ��S�F�	��cʱG�ԍ�)��w�ٮ�9�{�3�,�V�@:S�[�sM��j��d�V���z�Wr��N���9D'�i���vhR<N����ޒ�I�jW��-�*�b �'����׉��U��r@�?6���rv��K�i�ۭ���L�\=3�?sQ����`�7�\1=h-��va��j��mJo`�p��A$cOz����~/(�Z1e|[5�&g��$tR��IEv���+���K����Az���L�`�?#D?|�f8��#j��  "G(��L`���ct	�֩���h��Ѯ^�D^���<��G��%j�E郥���H�o,KR�P2g<�S��ڵ#���X��5�O��v�flm�"�0ջe������|����5sKˋ��S�||&U��/I�X�Z32��7�gv����i'Ŝj?+q�����W�([}��Ն^m 4#�JS� 1�ooۍ���D�<(7�-R�%r����Dg�t�=�����Έ/Qk�R����x52�t����]��}��l����De8��1��f��7я^�ה|m$3��r][�^���-�0���\�Ol�����:��]
��w��Yu, �����Zv3t�	�2��f��W��zj�1S����Gm�K���-�pv�Z��SVX�pGFTeoȪ�߉"#K\c��e�J	t�[��f�'~��:�jl+��vif=��n�E�T���i�>������C���ݡ�C%�;�͇����K�mQ����)jS���Od)l����`���##S�F�v�����֩�\���J��!q8�M��cNw3h�#:�x�J��~.�3�m]8��hЋo9�ۯe��$˛-:�\2��c� �ҠĀ�J�SG�f��e�0^�L�*���jt�y��Ś1�f`]��g!��#��؝_U�չ�����vMp��r\2 !��g�y>N�q礸��j��n��W�4C��;���(f�WB2h�2�����.?�<~"��?���#���\�����"Z�dLS
�Ҫܿ�7�c�f	O�ȧ�����\�����
8�(K���p����\�^�C����[QPF,c���f�%���xZ;8�)�<��/�Ԃa�g4�zY/D��u����~�� ��;��c[����9��w�A����T�m9v��	{ۡ���Ą�V��r��v��㓥�e��T�.���-�o������V@_��m���4�P]e���1M�:!���,/ �G��Pk�swybǣ݊#@]��X�!-R���T/�I��֋�,��E��3��Z{�U���A䏬B�Ҭ=#I���t������vO�t��8�S��?��z�+0�Z�"B�ƙ�S�K6>�kX��*��;Q�F�����t6��L�|�2���T0�-ρ�F�%威׋���r\�?�l��uq�{s&DGކl����8Z�����v�>;$���j�c+��vi���&���z��QSǜ�w�}O�������P��G��a/7햓ؚ�kjy+�MML��)��s�-]���+��-�Wo�o;���� J���0D�Cy�X�?L6C�^��|$�kH:M��_���y0�`�e�V�:l��q�� ��H_?| 3�Q����VGwfT'NuhF��D# �c���#oo,���G�:�y:�7F�i�Zd��#5�ԗ�11��>�r���q,�_�u��D�G�U5���f�K'��d��.�V@_��o2-�Z1Sڣ��"a0��y�]����;��!e?�/�wr}��utց��u�q�v���}EBWu���F�>唕F<О��4�6TA�uk��Ɗ-]�-` ; �X��<ȫrl��a��P��P�r�ʿ��ai �ș�Z�����FM۟��Ed�ﾦ�x& ��d�ؕ�+Q񰿗-VIo�\�:Ǵ �@�z�*�v^�u �t����XKg�k�9��1���������Tۍ����5���u�c�]m������`�l�r_���6���w��8s��Y��W�0[}���`q0XĉP�2�v��<yZ��8��a�W�Z~�7~]�������͍��ܿz)�J۟��*{���̬��������}eѷR��k=X�gK7�����,*^b�3�X�0��q��}�w�16ʹ�L�`�y�m��t"Ҵ�wW|�ߣ>N�{Z �E�� r��YC7�Ěz����YM��v��CΓ����A��O_<�o�淤}�H��;�8D��S�|�29��Ѫ5�Qa�&����<:+}�	ʎ�{�p}7��	mU�N1���D��{���~_u�(���x�cS�~p������ξ����ͅ�T�&�7g:V[�i+��va֎!�a9e췋�XH��fk�������a�g{�Y��Agd�0`J�:[ߺ�$-*����#6he��lG��T6Z]A�+�Nڊ%
L�5��*��Z�b��Ⱥ|� �[������~����W�: �O8�Tp\D�K����"(1�9mo/�sC�Y�S
���8gNwkJ�ƶ�T���)Mr�C\B�a/e]u|��?g����ٷg���ٹS`���2�O�+U��à��2��F��S� {[��x���M#_x�]y��3�=��X�s=��k��Ӛ������
�]��{e�s���{i$�E����3e\�����������'�  �-IZx_S�QeU��2�i�8�d�{�(�S�Qw&!��u�l�Q���z��VZ��c:+Q#�1�P#�U�����~��2��zh ��	�ѢEW�;Y�%LdJ������s�����|�>:��Օ����r��:�C?)��!`�|��m"�|�F��~��Ȏ�V��Z�_����Y��E��K/B����A׼*����HE�������$�)�`>�����/&3k�|�K��W�(�k����z������5�1�ڦTdP�
i �:ݗ�<qi���k0 ��lL�6�4+�x��ڣ8k�bRٙ�ӽ^� ��M]OH�<~�|��jbl������{F�#�ce���������4�m���sp�'>�3`�/�����E�r�t�IЎS��y�ݵ���+�Y�>���M5+�����_3��&�c��ʢ~ң��è厈,D�Y�U��N��o�zqގ������Y{���7��D�<��(}����W�,;���.�v����~dXyS4�O�����ܼ��4ñD�YU��#n�[���)Jg��T���%�)�s��hQg\�f*��8�ʀ����ޣ^�$�>d��%�-�=i�"�}q:6�m�,F0�[�p�>_��L���%��_D��V����ն���	:����/���+y���:���Ίg0�7�1f�����{9#�> �ZSw���M����Fg�+���E�J�4����)�l���l���Db�p,?���W�N�ge��UR弍�&�U�}���W�(�-�>3�_yn�}S�>�_�b���?��S�������0JA45����Sn5ͭk2ش5h~���X
�P�%i�����(�sL���}K�|���MF�~O��c�G�LбY/�A| ���m�9���x<J��0%/H�#�f��4���@=����ߔrg�2'ΓG�6� �A1WUCq��MT�<�>����	�U�r��ps.j��U(&�*�2���kf��قv�NP%����$��QE��%��-����/'s�ֽ��}d����Vz��S��2�u��)+�X3;��j�j+��vQ���,��N��>�F�7YSVSє���v �}�˲��ql���QrU�֫.l�ڀ�@�c\*	�gJ���+�{ٶ�6�96V�:�8Y;����ZnA���F>HoƂ'�����D�xZ��m+�^�+`~(�7��cW0��x���炑G�^.x��Z�2)�-�{�$nb������G���F���^g�#"����G�QG�n*eҷM�Hާ�9@c=����L@4 ��À���؈����}mH�����Ю���1]�\"�
|�}y�-�1��;ذ�s���:x��?�)��R �~��.�V@_�l��T� �L�y�f�S0���6h��SP�G~������������<�5�6R�H�A�2�/�&j�W"I���{1�MPu4��j�Z��cN�{
~�&��Έ���6������-޶[�O��ֻAE�u��|Q6�%]�E�`����(w���c�Z�M>�<����m�$#��L�J������r���F6���h�y�9	��4O��6���CD�}4�W�_���(Y��!aЦ�a�ΐ�q���NL
�N��l�ܨ�)#+��^�� �1d��k���n����N�:�]�y1��G�J�HK�\� ־��.�V@_����*��Q�GJΌ�Hj(Ǯ�M����;�B�zB]A����������
��P����N#;�UiK��*?�LG<-�`��Y���Ĺ��$���~�]6��������|]�
�r,`t���tP"�}پ/�G��xW�	3��� ���z��Ϥ�X1;�-W���2^icq����N��;U[:r�I��k1�[����P���]�p{/mPu��@QSc+���	��xmɶ6�fX��L||�����ꠓ��92)H��ZȃN�#i���^���Q^�:�}�ܑ��c�^TJ��s��Yb�wWr[�Cw����Aq���߬E��.�V@_���:�$�~��V�nK�ݕ��D�Á$�C���Ͽ&O�<���bZ�"_�z��5�]q �c?	�l˾���t+Y�2���I��?/�������-�>YZ>��:3��nH��:��c�H���n��́I�8���N��D-��-L�Y���+VF�m�8������
cm�#8�&+��ܺ�"ʮ���\��B���ՙ��:x-9U�9�}�V.�ɈΫ_�����Iri�:\��dƹ�=�~0�[�\l�*�s�7q�\��#�[�Nͱ멫���̂TQ�ӻ���W�,[}���#��z�W Lot��x$�y*�?vx�J�����|�7��rS���Օ������m�)�DıWP����p�I�S��7�R�B�Iv|�����6J�����fT��:�t����|�J���+�L3yJ�}ĳ�i}�g�mwQ�vtj4ͬ��+sZuu#$�e}9��tᏨ��)��� �7ގ��3��det��̄j��3x}���%�=�i��Y�w]���LI��YvU���	���0���`�X�\�&Y�c�g�oͶ2�k��ymˁ��r�Ǖ!��E�
�]����Rk���%L�H�z��/�O�������_��P��x���gmG�� u��	���VcOe�xeҧ2����S��c�d>I���Q��;:c_N���������2���cq.H�ӲAT���dn��e��h)�;;Gs�h����FU�>2�!w
�8��@h����K>���ͫ�5���Ѯ:h�c0ȴ��+��J9���l�^�A�Am��ɮ=��Ѯay"��tguzj �0j6e�p%�eu�*��[T�$��렵�.�V@_�=该2O���k tD�藞��I>y��|����ɳ��}�C���K�)�o
(� ���	�S��2�z�L�+%����ҰS� �w"�OKY����*��PM�����-��A���G<�4r����Hr�^h_����*ھ(;G�d�e8��U���Mо:K"�ף�Wt�C{��5D��ޮM��Gi���X���ϞYў�l��ܥE��烫gu{M�i�� �ȶC�~�Cєxms�u�h���E�|��.�k-y�:2}6e9�F04��Ϡ�B��=�Z��1XS�]��������9:��,:�q���V=Z�K�v}s#���w����GM�)XL4[���z�g%��/"@�Y�7�iN��,~���y�6/���`B/01Ǒ�f�i�DuƳF���Kqk�d��m����+��-����B�O�J{���L����I��b)!i�����Q�H�1�X�}����9�%Z+�̵�A��o�b�LZ���^-�=���`�t$-�46L���f. �c��v�j���O��s&zX����y �@�/6�r4�����q��~���j�f� �	������4u֭el<H;�R�A��w~S��������M%�WEfd`d�H�G{��{��H�i4<�À���4c�4�\;��2������X����8�=��^L'7n$Y�6:aj�B=}�)oL����������AH���.^$&�b	��A'��9��U�6��U�El�0�4HE35�9m��:���t9o>sk�#�âZ�
�6A���C���f���A�:/���ߙ�Ck��/���QY�R�/�PPb_�irV�'Y��*.$
�֞�F�]�����EY`�t0Lɯ�,��Q3�k�l1t
f}w�ts�q��W�[��*8-r >ޏv2��C��Dr�A��g�*Gf�˿zZ��)���p����j�ԗ�sy�461�'�z�VD[�TUNt�+r�]R��@@eTPCVbtÔ�?=���g��:X� �A���ؓ�c�T�M��5��t���-�cO6~��䤙X��a�3�dX�Ae���,�-7o��V¡~1�,b��Y���R�-oJ*�7M%MLZ'��lu�c��y�y�,,Q�z��|��'�[8���vy��jf�5t��@/�`�7�1F��*�=���-�!�]+o���O�:��C�M�� ��_J��ia�T1�p}���63Xγ�w��M�{.LLm�֣��,�W����:p(�~4@T���3$��#-����r8ԑQ��
��U�Qx[������jُNM[������qz���4�l83�2�!҂Q�P��:���rӶ|@E��\G��o=3�|�m/i��8���8Pc�������$e��}kZ�����l��`n���)���C�.!g��<+̀d��mO��@�Hv����T2��V�([}����v�s���wek'�T��Xۺ� �/}�۲�����^ɠ�i�=�Gé�gt�����)k� Jp��G�ڙ���;��F�"a��4`� ��9��v7�s��r_��m�io��%7`_������ܳ|��.�y(�iK�z<(��6�!�dS�:��O&�������vr<�8ȱ?�a<�zۇNt��<l�r���Ecl��Bi-������/�|}οa���:���UN��>��0��X<��W;�(���C�m��qS�����d:a�D9 �@^q}��D�1t+��va��j�+l"uY[��gjy�W{�'HUT!+���/���|�B�핤��Oߢ�m`��ȵ�'R��Eԕ���ؖ�k�J�	�Vwz��(/�@�2�	�r�	&)��i�@*5�����p*�xlvd��o�/��Ṇ)d�8G��!*OyS��� �`��U��2� ��W��Ԡ';��ϒz��}��;UѫKd^��i9�MY��-Ȯ�嚎FMiW
� �����l��̳��7�;Yj��g�_:�	�e)�Z�t;�pԞ��y^]��no�6�妪����n�%��y'
�^o�-k���=�Y�1���t7]���W�([}����j��~Ѕַ�I������1�ݕ�z�@>x��/�&KS�CBZ��P$a�����,�ю�y��]�F�r ��l��4}`i����9`R<C���C���p��؂]P �0P��~�I�J��c��nJ�y{O6��"�jT�0���^���84z�A0����/n	vm��s8`U�:��@�G�"�?�|.�/>!��)���^��̈`0wY��8���z�X�O:f.�9rgm�J�����m�b1�ev,=҄8gy2��+N�k������o~�C���P֥��/�N��]q�0�m���0��+��g�s��8Qn��.�V@_��,��͞�}Tb��/�����F��}��[��Y�]��M�;C�<k5ۭmo���Үq��&='m��گ$m���o�7G�a"��4E{����z�W�s�x��
Ju ��(|��Sy��l{\s��P�ǃ��^�6��jM2���?�L��<��r�/��ȇ��5���Y�]�
�y��}Hr �Z�8)�9���p,�8t�A�kJD[�Ry�����a��"_xE���!��A
� ��x��x��A3 �;��]�e�8��c�k���h+�_���'��SǮ\ۓj+_�>���+i�yGrY_��5��l7[:t�r��<��f�2:[��A{ʡ[m������eY�2�)�O�ꔬ�i��r��NCʸ?�L�b��%
�{�R�`�s���}�`?����6zT�yL���Tx��hX�e�}�V�3����~��@�'�?NP(��JL^y�^���oˣ'���������2��>����W��#J�3o� 6{9�}򛫝�~�[����<��<�>␑o�տ!��o���8^;Ȇ`͗}F��d:Pw��7e�>�����nȜ��7� `#���df]{^���y�f��iu��GQ�F�ќ�S��ʾ��I�ǈ���F0~����W�~�G�����[���w�+?��d��3y�{(�%2q��o�Rh7�8Xg���s'o2�~-������W�0�
�aYC�Z6�]�,�2�]���.7�z������'=�{��뇶��Ƀ�d=7�pjn��G#Q��`N��4�-�ZU� ��~h7 �9��D�%��U�?foz����Ih`�W%��.��i%��|�w~EB7�M#\��g2�1�ZH��62B�tm#_bz�*Q�Fڗ}y��ݷ?(N��e����m�6#༢��h�g��H|=U���F\��5Y��D��@)�Ѵ�4�%*��*�S~�)�P���s �1�oJ�;i����} �A�q�Y�5��������,��w�c3���-���_�a������G�������՝ܗ��<�!!q� 5�]�+�NW�еk���e�
�]�!>��o�I�icj+�#:�cL�B���������e<8a� ~��g�!���r��  Z�(\bd66�T�3 òX�R��*+�����_c|�)� �p�9��kzCgBqHB��[%�~��q������K$�Gu2Hd��z�Bqj��w��4���Ԉ4˚\��ꝨN<��G7�2�r����~Ǚu]���V�'@����T�r�H���3����p��s}ȼGV�=q�(������u��纈��/~'Sl�k��f�>�5�@ikѩvu�2M����8I7�����Gr������/���o����W�������|����;��O?�T�2�Ҷ�7�����3�KYm���W�(+AO8���y� oM0 �帿���g�v(�9�부�]'�g/��ߋ�|!�{�վ���+�=j��b�'�����
jݱ��Eꬽ�:���@��g���F��b㧪=JO���4�-A���^��/��pgjmB�LL?'MGC��沶�����My�H�zj�#E�1�6�B<H�g�1/ʯ���^v\�)�>��f�L�dg�%���B��vU�Y/O�8���hg���e�|���t^��jS���@-{��v��XG��t̕�7�r����/NN�y�����V�)}�R~�/�������������/�+�-߷(:q�FF�8L-���YjXm�K��W�,Ӓi���2��X�� w�^���F�z�ы}_"�{i>{.��@��M��߃E��"��k��{� Y}Y�]F��"�q_{����^��|?�N�,�MK��RL�}T�N>��̪���%���!�r�!�Ca��G�)~��G�tr�,��� ��m�'NKc�t2N����Q�i]���N,�5�d��$���c����zg�^��s@ߦݰ���z�����(LԶ�br\�
���5<�z(������-��;�˟�/������7�K��'�����l �q��W�4[}���^��:���x�"1�^�,��B�j��7����������2�Gy�Ħ#eBt�q���cֱ��j�Kp~P/�F˖ۛz��=o[����52XX��Ν��k�iSâ��;�}Q��{�<�r!s��$����b�_�kN�� :n)���w�T�N����ea��
�&�;c"~�d�K;���:͊!�M?�ӧOYba&'g�< f|
ȷ�f@����wr��F�������u�@�z��쏃�[���6����]�����EY����nFY��rF�u���� ����N��A��?c�K��F�V��Zj���4V��ܠ? \s}��e����<2�)`.��X��9 C�捚�fK�ز�����%~R����|��S�</S4[d����!.�+��t�3;?��E�;k���isA�><E3e���5����y{--��J��q�<ǚ�8��c׷�xPX�ר�0�s�済��C����J^|�R�>~R<����W���|��w�o��"���3���(u��f��]Iq�]�����eYM�*z�S���� ���%R� jRn��ǂJ����%���ٺ��ZT�|�J��Ekֵiw8Q��40�Z�Ц �!&a��e�� b���df���S���e�k�Z2�K�����m�juӾ`m*#���ie��>�i4������~^�F��<�yF-�3}���Yg�7b��m4����ܥ����rVGK���pxB�8����G����'f=����\�oH���.�I�?�ێ�����7Dszٿ��|��;����������~?����mK��ɪ��e�
�]�!-�����<�ە���ۺ'PU �� ��<��7���Z��٣,�C>,9�3��ֈחѷ$�V�&���'P^2ח栃�X��/#]��"���2�����~e�G��S*�����0*�ɲw�;?���tӗ��<_3#pS�[�����q�׳
>�}��vH��yvc��˶�ײY&^���v0��h������oJ�}`J@?�A?| �rM}��q����?�����ʧl�2� ���J��je+��vQֶMuu�oʍ@q��2rvp��h���-R/�K|�JZ��]]����� ���U�l�����к��h�)�6��u;I}8Ta�w���يv������1O�hlb�)a�y��@y
��)��@ЅY�05�	��T/_F���۱Ҥ;����58� �6N\>���N��m9L�M��l�G	��])����S�,g��|~�m �� Y�Mh��W_����ky��|��OA"|�h��#��m�\m�˱�W�,�B������%يLnD��F�hX�xL�t���@��-M;3����[NA�E\P�o�y~�[�u��h����$n��C�(,�-��8c���	<hٳM}Ԩ�=���4]ֻ�k���n��g�׫%�S�����5����C���kR�{��Y/,��i@��\X�����9�EC�N~#JG�D�N������w�P�k�Wt����j���:jI  q�IDAT�?��vH\]oK����ɍ������MDUHV[�l��.�P�����~/�?捗z����eD�lQ*7p�*�\u���u�;}Ӵ�j_���T�m�i�ڢ�ƈg�0N�ü��K��'�k����IH����+]����Mj{=��z(�ϴ�������v��1pl?����s��+�_��)�Ua&��i�R�J���2����u�n���u���k�5p�q�M}O�tJ���n*�����2�ܽ�mo�y�9$^��l�[*ٶ��p�ڭl+��x�M���e;._A�n/ҁ
ȘWo=(���]+��vY��jem�tϞ=����'�b�2ɀ"&�cG�{	�e,�����RF������^�7�ȹ�oJW/�����m����������/_'��՜�O^�7�@XWs� �T��E�st�4B?���4�i��t\q�0����syS�w���=םjy����~Ys��9z۞�|N9 ��E=�9�׺�)#t�n�69���2�c(m�g�� G��s9tX\m�������Y��n���Q���d@�9�0�\C�rC��6�,m@G}�3Y�� �Ƚ�`���MӵNs��T�������=�K@_���w8U?�s0�s�@vB[��U���Y2�ŕ�D��3�<�����kQ� ��癳}�y�~-���דҜ���s��z������|A�]х�%q<[�eB�D��x�סM���pbߨ]ɘ|#�c�3�	���ݿ|!y���kdW����2�� �����
�]�Kt8t�i*��|x�@�@�N�<|�X�_���g���y%H���j��g,��X"u��'������ނ��s���j')��sK�9�1+��F��Q:�<��P�	H���^Kί�v5�5�%��l.��&[�2��y$_ɼVΚ??��O��k�������}�c����3�wq8~�/�C������br9)i�$��7Fض�<|x#��d�l�}���^�u��jh+��vq�1m�P�Б�����ߖ�����r��r���?�	�,�[4���"��Ӵ�"�׼ߴ�F�3k{�X毟��7,��4w1�����E���̰7;>TƥR==��Y�gܑ����L��+AN���)`>�b���� ���Q�'1���h�ɺ��QƓ�y�`n�Sr$�4(�pbR�m�������(��GA�a���\�|�;�%O�z$M�h��rHU�~W[�l��.�6�m��*�q����g��'���+��uus-�$�|�b1%2�F� `�� d�~��ǀ��2��u���nfot�s�_F���Jr���7����x˨]7����;'%�<������Ҳ���ֵ近��y��1�i�J���%{�{0n{��y�Z^�W���~��`}OR�^cϳ~[ Ӽ�(#�4�rؔ�VgD��3����š��������={*Ǉd��ֳ����r_�l��.�H_K��P%=�Q�yeΚM+��+y�����HU��y��ܮ8Z�5 ^ޜ��$0�X�7��cXD�¿�)Q����l�ˈ})��<�[��k �[q�l�R��x�y�� �0������r�x^nX:�3XOv�~t8C]�9a:'#�����m��k�c=5�'�;�j��y�2�bW�������i�\	�q��A��-,���k��^��h=��
�SP���oل�P�>������3y���^�(?T���A]h��.�V@_�"́x��w��p��R_]ˣ'��q��>�����<E�)L���Ka(���M�"�?�Ѥ��v=�w�Q#�Mx�5M{赱��dH��S�{�_�F#�`%�G��Փ���`��Hy	��� 	h
&k����ɥ�=���9���#O�6A-|�s�k�G%�	�&�ؙ��U�]���8�q&�`��2��/`�ex�}!��F\C%a�O%f'a~=�aS����H
�xH���2Ο�eY���ݫ�r}}-��k�_����E���(�����W�0Ӊݜ5�>�j\�u͡;�l�]�a���<|�m��r�~kw�T- ��(��Kr͛=�dИS{�M�1���1�}`x�t�Z��CFF0�pq�K���J֖��h�F5�U��,�RW[�?��������Qwn����AX4�����2NCE*��q�����6�)�Z ���L��`_ְ�q��y��d耞LK��י�$q�W=��򕾞� ��v���E,B�:'�>/�ls���Q��<G�oUM$:��)�8V,�@�Y��C�BC�5��v'��^Z����lCf���G�.�c��܍��1���f���g����V@_�¬�Ƴ�{�`Fk�ZO�z�&���i��Q���m	:L�ƙp��$�g���[gG;dC�?W1;�_k]V�SҨ)�1�*N���8��U�&��T�ƶy�t|������WZY� :�T��Zb��q���ܵ�]).U�J7N;g��l3�+S�k/�["w�¨��eY�>&�G{=�Z�u%"�z'���'��%��9���M�Y'pfĝT�'-����h�=����zjs��ߕ�M��^HI[�(�[�@vm�CA�Jr����[�x˟1S�}��.�V@_���¬s����52;0z4V[4��tl(��J� �	k���O�>�i�w:Z�c0j��������_�ɂ��hҬ��e�vX�Ͳ���O�u��n�% #��L��k��!/�|�r���<���S��)�UNP��9\?�e�hO��������� YtO��h�J�j��7�i��PV�Y�iY��>�5��b@��W\W-'ߏ��ߦƾ�O���kX�ml�����8=�L�~Dͱ�wfb�σn�G���j�]����ڥ�	���uSpU F�x�l)4K���u'8�.b5Ra�0�[�����f�EF���������R����,-bkD8��/Z��"u�Z{\Un%*@�����,�����0 Z琋uGkZX��Dr�Q����_���ڮ��@�����o;��l��<9�z�+#������taU <.H�2;G#R�彘w^/�s�T;Η�b8�����
��+�!	����a?E����L '���Ή��Q@i���Ƴ.�1}�
�]����ڥY����~*R2Gp�sn}��5&H+�3b��e�qφF8��}��轴V�E�7�QS��2��t�	,zL��xʨ�����G^H$	mB֋�2�v0�1N�*T,5�Y�1L�*Z4O`�6���M�sG#Z!#)9-�9U�)n��B��2iZ���<��>�GS�� �ffs�ŲZjH��I��ϩ~;S��@���F�8c-z��v�p=��|���69�B' ����B�aqj��{#@z���1˝�jw%�qyC�Bp.�j�]����څY�`�4���Z�? �e��"}��'S�ؠ�ɿk�U�c��Xk��R��&�\�z�F�3iN��q����a?c<n����t9_��`e��Gi��i�5>B�eWQs�I��~�>���B	��	�1LهZdr,��}HÔVf�a����2d�c�x�5����:]H0䶢mtѲ���[�h)�A��Aң#��5��L��7G��(�����@���W=(ǡ)���v2ԕ���k�V7���	� ۫������*���.ϵ��W]��.�V@_�ҌH����T>�|�;9������	ajczi�Ѵ�ep�02�u�ϰ�~�ک�e�k�i�{��4���p2Ii#�'Kh'F���<]ֆ5�����n`ҟTv�ȳNy�Z��Z���E����Y�&z�'�9��A��sT硞�c�RE�ط��lr��׭�3�W�� �
�-@(Uʞ���>�MlG��4+	h�	����qя�N�JU��W��vW<:vNĺ�T�(�j�yO���E ��8��W[�Rl��.�r*7�1�M�i�[k��R�Ul=1�,��.�n��6�v��p�8R'Mq�������U8X���Y݋�(������v �?X����;�}�4�(�^��r�x6���G����ґ�ld��)u��;�X�#��*O=��X�a���p�s�dn-s�������7����CjXə�R�����e��5f�|	�蔤�I��m������$��W|�C����?�!��ۆe�[LX���$cӤJg�蝐k�}����W�8��s�ܾ�ne�+� �(R����M[n�*V��mL�Q�DLF%��#������#�`���6����Ϯ �ٲ7 %\axR�>k�詭,)�n
� %:V�-��K)Zg��Tٍ���(�m��nD�p8���R[ym[%�x�CR>���=w{�J�@A��w�3��Em��g��S9΀�7�U��꘺�Zߜ���=�ei���g��:�vGG��=df4Т�|w2�H�����,M�5,;��U��Q�QQ�×�?�)���ȉk�N�}�_���p�'򸋟�W�8[}�K�C��.gXQg�}@��{( �=� %�S��F*-ڕ��`�l���!X�6�"b5^��I�}�'�{��5tı�E�Sԟ�lg�΢9�Һ:��Il��bJ�i~�da��q�>=��_E
�$#����^x���af�O��]���yA������;�5����N�����'��2g ؙ�q���8> ��c:� ��TaN&R"�D>�X�<g%�d��, �����s�%_,D�p�z�Bh�@����jP�z�w��2�A
���ƾ��V�([}�K�r�J�γl��5�Lm`�%�u���Z����0�n
H�� K
�4�u���Ո�b��G�zF���������1J�B�ZQ���:"u��*�γ��;�e�Ǒ�1���RAy%����E�$QOAS�n��סy\Y:B��������m���8��9��:D��h��D��j��ͨ��^�	�Xo��ُ�8;h�"���)q1q�6]dT|,��f�������)Q2���`�$h#���@�}��;<�:�}w$�S=Д�T�G����NU����V��P����><y�dm[[�l��.�Bt��Y4��sk�ҍ4bm��\�������} y4$@��P@7o���LD�mH�N��yb�/&�Z��8��S6������@�5aM�,�vV��5f�c�
)�`��G�Hyk�~�6�2��A�j��'l�2O\S��z���Nىu<�k_h�35M}[�h�e,��[�����Nf��ԶcV�ⵊɪRa�8]9��Y eUo([m���m��(��H�M5y8n�O6����d<8u�4����rܮ|7�a4���f?+�y�"P>�*�����(?�����۽fa���%�����
�]���fړ�,c'�+��ԕ���F���`�m-ՋHw^�|��8_�-Vh{�l�-{���u6B��Q�'�`{{��Q�8���aV�����'�e��_�<u\�������ɑ�@$ZQ�,yN5sT��b�~����s��JyNٮ�����@�6-z3�� c���J�!3V��.|]�f���tm� Y�o�h��F9t��}:Oϲ܅},K�����iӶ���є}�VG��8���.�s�!��a�k�׾���	?t����I�����e�
�]�q�U�5҉�U�=.��x�_��C�d��vn�@�͹S C�?�Ef��-QV�e��tާ�ޔz�rҖ��������qx
Ĵ��j�Z������F0F��j�*{�p=�[�2��q&�Q������_��{��9�+�㞧�@��ҴV�d�	���fW����d���dJqd��9�xX�n�'�-�����\]]���I�QF�5�~�,�K���e-!$�ciUvCr���Y��bd9��a`%#���FL� ��}FZZ8��S��Ϙ�nb\w��Ճ�W�,[}�˲C�rm���^Y�
��ޞ����[O�����)‛?�=�EMA�:u��^Z��ez���w:�0E��:2��,Ԃ�H���� ��A��Q��`�[d�~���HG�`?�N���J.`�1�� ���V�HQc��`"6�a��N.�e6gd�[}n��.��g���Ȏ��|���˵��Gr\�ڥtAb�o���Qa���"�����QO �R0���WT�!�s�(׉g����E�.�l�@?��ɋ�����=#��J`	�T����,�`ꨀ)�3?�3ַ�3�p{?{��C_�l��.�B�H�'*�;�"2Y��PٔJ�P�m���G�`h�(�ϡū�@8�'RU��X�0"����Ȕ��h��գ����Y�xWn���-�Q��Y9��+y��e�;���D8���*�r#��V{^D����L+
4��+��/~I�^]s�;�m��L��۹,ws|����CB5�	��T��������B �Ǳ�ï~𭲦�x�=�I������N^�44Q������߳���G�Ǜ����'b/��0����l:]�vD�;����Hn��~��ŋVv�LM��)�H����-�|��@9x���vQ��j�e���q�U����Qz�l�X�%2od+5���r��Cٝ�c.yԱ� ��D�c��Ht�KV�Y�S;�P��ĶlѰf�)\BQ�s�� �;"�lwr��)�N =UBCD���>>�1�3��*����g~,��C?�"����7�8���UyNS���O��٬�
o.�B�;��}�J��lHWG��W�{ 0�!���ɢ�]?1���O�����X$���y��{uK�� ��l�����'����z�%��}M�Iv�P/��ȹ|��x�����!K>p:Dw���iv,k���rw��V� [}�˲�H>�2iVy����)�&�R �Jk̈��#<�1!+ȡ�|A�ͦ)bŰ��,�Qg}7rΞ�>/���R�>r��e�E�Όt�c���Z�B]k
�HV�+�*5ZKe�g4���ܲ��Ⱥ@���r�m-6��j�F�[��O�裫؉qd��Uum�1Ng&h�>�X�dD0J���;I�pB�N��l���eQ?G�҃9.S���\+�=jݻ�Nz�d8k���O}.���A�!뱫����8��)���'�|g@�C�!d���֦g��$���@�i�ݪ ��ư"{�P�\�_W�([}�˲��JD���F�����'��,���
�4�p�ܻ�^��^v�ʇ�?�6��g�'�$T�66u�CW8��R�u�,j�M���)Y}ݙ��6�~n}�����BN�rњme,��j�^
 aKĶ��cը��"�\B�j���hK^qJb���2�3�猃=?m���X�#A596�[�>F�޽�@#զ �Ҫ>b���;�����7e�v���u��|%u�T�u�}6�[��5ݮ�.�#F�T��;N����� �wL�C{f?t�g�-�)�l�F�IZ����{��r�:K���Zm���W�,c=7�rZ�G�j�Zvf:t��Z�m�>�L�6�L�������PG���ͺ�G���ƃF�l��~kgc%o[��e�y���%&�P�b�72U.�����Y�Ǯ>�ii����:��
'��V��S-�=rO����\!�k�K;���':���t;_�t�����q̬֦�aC.Be���������!2��`�:D�k+ [�hk�)k�I��`mu9Y[��xc�B?]-�+��L��d��te͚�*?[��Q�h��{U�kLH���!��4�S.r����O������Q����GO����j�]����څY�<�Dn�����k-Bj��뤺z$ͣ� �A���޽�ݦ��jE  �|#*' B�>2��	ed֣���9��}�Q�a�Y�	l�2�f�Ϟ�HV=������x���9f�>� �����\$UK4��A���H&wA䜙o������pڏ�,��45o����9x�������ѿA˙e)�)�Ѣv��8�#C1�UN3���W �� ���U~����d=�oH3��r��m�g'��C��+�A�gy�z顣_�������f��Ue��e%�A������'O��#�{�H�[�M��~��.�V@_�J��8�O���� /^�޴��E���oʏ\?*QW�>�f�D�冽}��8�q���k�����`��6�4*S��i�{�T�UL�5�>"ܦ`�7kLt������ݍ��"L3W����s�D*(r%r���jj�Lyazԡ,�{6�=��Ѧџ2?N��ϏFl�y�yjc��B����+��W�ё����5��s�^��˶W����4�J��}cu{����W+8瀏K�_�G��]�OgCfe�}��7��w������(��|.�kyq�'j�C�_���Ʋo��K������g���a�Ƀ�Ym�K��W�(�u��T�Y��J�ך|50�U�;�#�O���������oɓ�y��S�77�ñ���(W��^����+L�#���
�r���K�� ���B\����b�7U^���;��)v�m+���Q2g�U7�v*֛�7|�QV��Ñ:�CK����2���TϜ V\R���M(����u^��L�=Yk���a�)����ֲ�|T�!Z�E'�ٹO�����@7@	hp��6��N�2��������X�"1�Y�N����١zRՍqn���ȧ�A>ٖ����ǮٽEU�P ��#�3,�(���?�G勿�k�Q�J�:�a~,���f���5B_�l��.�rN�����Oz�yG����<~��;��"����n�Rc�i�9#2ZwFd�����| �}��tw�jo���w�5��#� X�َ��/@�ly>AX���ez;��)#��#8���EkÌޭ���mT�S���ؙ�-"O`ʸhC����J�>�v���-&!�`6_��r�W�	�,O8�A���lo�9"���6'����\����ep�M��D0�!5����i��"�����0�z���- "T�-�����s�Y�y�D~�����������C���.��=&���ل�����}���O$?���8�h�ܔmЦ}{3�j�]�����E�f#�9�j�;�f�m��7�0��V#M:4;�`#�����X���ϴ�0ӻ6*�9������o�_�s���:d�%�U�a/3g��h1ڸL'���q���6�O
DH\�7W��/JƩg?*�:� !�a00����`���v�c>f��:�34n拗}4�j��_�Iex�v:[\Veo۲�)��]p����E#��M�CT�'� W����\=���w޵^~�~L'��z�Nқ	�L����e���}O��/�#ySO�
�>���:F��ں ��H������X�?͓������;�G��K����*����������(��Ǝ�9�;����B�j�C��e���꽬���
�]�=x�����_��o|�O<z����&����{H�&C_���Qk_n��+�A��8vG�:�N³�������?���_�Y
���wGp�Ȉ�I �I�;Ou���!{�(d�ށ(V�����ړM�Wh��s�A'=��uN(C�U9�]�����3M=DH��u{�i�u8r�(�u'�7;9z���J]����V��(� ��"'�µ<�l2�*+�Ϙ�0�{.�\G	�;^�^B�g�N���l�s��D��{�_��7����Ϫ!M��o���g��02�~sP�;ϗ�N�tH�i�d�w��}�R��S?)?�'��4�#���y*��kѫtZ[�Xv�q�l[>��� o��T�ݱ�=�����d��.�V@_�܈�V��o~�[���x��7M����:�'�f�;�2��xsfZ�\ �����ػ�Ȳ ̫�^�r�~���O�G������/�w�����%j��q�J�m#}�Y���l�5Vl�! &7��W��+S��w��-��z�I�f�?ǹ-��꤯J#���X3�\����Ӷl_�@u�^;��_���o�5-G3k�WF$�w{��TW7r�������S�'h�]/�8߶�(����G�l�K:��D��(�C����Z���jk�Hd-P,�[��Pk�q�XU�O\��nQ�~?,R�NƆd>m[SQ�������͖�?��?-�gO���[9@ÿ�<2�IPǉ�AtB�7�nK�����+[}��6�P���j�]������Y�W|�[��_����(�_+7�v��v*���5���y�=�%�ie_�aߦE
˴�����������t%�z��E	��U��Q��L,��}Wh�*7z
����t:��չ�y\�صM_`αw*��כZ��N&��H� #��e�SAZzT}�r��ȓ�O�[�����ȯ��7���k?�H=��Z6.$�OT�������f8vt ��5�����#e_���"֫m�,%(��x�:7����ￕ���Ei�v��PB�T�����	�|_>��c��f�Q�a��y4�0��gȎ��{���������~���=z��rM���je+��v���;_����������,7��V�Q:��D��)QY贫��Fĸ1c�i8���F�m[Q;� w�9�s��z���\��&H1r��3�NA�l���SY >mW�2ע�,��D���b�+�k{���&��5eF��[�cd=d�<��ݫJ���O�ѷ~]����R��|����}��+��v�N���-�U�y8y����r�yr`��fM'��r�J��Ш3`�� ƾ�놳�A�Hv�C��M��O�F�[J�&�cZړ��ؾ��էt��t_�Gr���F����|�z�Q������<�=�s幗��jf+��v�Vn�C����7��Ϳ[~�P��$.��*��a)��2�=Ⱥ�~Ȳ۩�L_"ʮ?Pt ���\�\��}�����fW��{�߾���0P�U�t1j5] )���q��،"��G����)���2#��C�,P�y�s�݁��o�Z��2
�o0�. �����҅A�}���	ԄxsE��p�^x��/��S[]������3�u�p$Ƴ�Ü�_:?'�gA�a���[��h��HI��*؁7�V��n�x��(Q1��<mjI%*�m�cP'��>����,{�� �����͍���}��g���{_�����~UV[�m��.�?�?���Y�V���Sآ���2�r�'�e��TA���7%2Cd����ϳ��MJb�����z��w�z����0�0��ӡD����~��
d���8Xg@�M�y�:6TJ�]S����n|��F%<Y����/}��_���%�.�~��������+���oO���9a�N���|�����$.�*�����[ �xꙷTFỏ;y�����;���!͎l�q�#�y�{�+Az�|����7r�n9f9���+$��L'��E_?�c���o���=y��+���(�X���v���jk/^��@�R�!W��q�'�T:Ϛ�)��6vT'~�ϾDh�S�8���|���t��;�V)Hd��LfC���Q�(2W1�����֗��2�����߶�z�z�^�Z��?��dJm���U�lb��~4�8J
:kf�mu��A�Ƥ2��|R~�տm7���O�@@��z��uG�d���ljyK0_f����É�C���h=[(�A@} -�}q���4$�0h�2��DY��:��B���s��80sA:�jT�7�=�v�aL�v+�wwh��L��"#���^�<z�k��/|��6Ym���W�X{Tכ�|������; ��� �Q1�?�t�3��
z��%ʉ�T9sa���`m��휬����!W���7�����qׁ�z��q;��m
(�Y���Ѣ�M�b3�&�'in0��uº����l���8A�<�X|-��
il�lw0�$�@�+`������0J������9ID��l�g����Q�Ӥ[��|� �QZf�8fY���_�e������*���><��K�kψwٔ��1P�c_q�<v��wL݇�%�O�����>���ܯ`��E�
�]��c%�F�g���ק4��o�H���6CSa3�+O�@U˽��
����m��AXd�T�%oi�S�2-��,��s;ѩ�~G#������t�z}ԣ'��c����Gu���O�����1����A�V�_�����-�2��3J_����$�f�7�q��҄zq}���#�{j�tߧ���ZO[���Rޒ�w�~w'L�q��w��E�
�]���!����&0?�}>�����,X�Y�	�,��^�E��2:�:�yK�o�<�s�^>�~n;_Q1˩U���K��uX֓�y�}�����|;n�&�����kZ���Hk��}���63�g�
�َ�������I��yǖ��Mv���õMm����W�dSq��{�"���N��Ξ���}�$U��W�ݓgvfg�˲��MDD��   ��~$^��ǀ��z��E�"ȕ_Iꕠ�p�Q`�ɛ�����������ߩS}��zf}�n�~�w����+�sz��˟�ve_����E����K�6�a�7��u�"(������|L8�:����8�b�>m��C�q! ���]�=�_\P���Ǐ1�S�Db�[b,���_{�{W����#���!�.(c�Q���I�a���EW���������ʍ������f�9�ν"��(Jha�Y�;�5����L�N��J�,9J>�"�y��1���~{���� .�X����
�:��5��z�Y���z��pܽ!��߅Y�q���?��e�pL~���/v���>ֱL�q��97,�b]&���D��s����^���k��/u-��m�3�ʍ[�y��$���4�����i��k�� {��b�U|�:<�K���b4K��^�8�~��&����eg���R���M6���;l��Q�ei��+�l�!z�m��!כ��ne�1�Z�ٟ��Eĵw�Wз]����̾�q�����͘��빖�L�FX*^C7qMC�/P�y7�h�u��|XRּ�'H��sM�f��mr�Zb�s� >{�~�{��3a�A�B]P�qri�F��F���6Iǅ��8Y7�kz���k\�j�I�X�U���U�&о��&uS��k��K�[��q-6�����e�f5��=h���`&�4���Ml¦7�Awq0q{!����Ԉ�.(o���a���w�}�i'�ř�qL���j�2��fw�%��3H�]WW�����h�aH	�{�ۚ;k�i�������;Ĺ��4y�EB��p�����5�l6�5X�3P�}�s�W��Ua{X{ݢ$���YW�4_1�l��-�hK�`�'���j\k?�+�q1 �m�a}�q?�=���9)�ڇ�B�����:N�.I�w
Y�����~���a�d��@PB�-��5�s��HJ�
��K���0n;~\��@0 :p�������m/�����)��I�I����W7�a\����s��{닶���-�ڿ.�����o�n�[@�z�Ċ2��_��e~)�Ĭ���m�(L�ƃ����v�v��)�.(o���A�Rh:3{/c��L��~��{�n���c�{G��6s3���!c�60��s���n����D�{]=�xT�Z��O�ʖ&�y�5)yIf�R.�RV��ݶpDH�?�᱆h9�??��Skj�B��ĭ��,��!n��{��������ȵU�u�u2_��
~�#d.(��P�PT�U豴�$�i���ɦ��@lҷM� 
��!v����k�S��5�m4w�0�o�Y]�	��(GI=��m�J� 0&�/߾n<z�>7ɲ7��q�z�kQߺY�p=]?�7�;5]Ѻ�:�@D�����j�0��Xc��	��K�%j���ў��У��Gh��!�.([8�<���8�������L�q����U��#�fk����n��A,x�$l�L��6�<��~�AU�kP�c���֋�
�$Y%l�5B�9'�{_��&��>s��nH�h�Fȱ��2�u'�^����sY]�ao�&N�HS�L���~���TDދ 5��o���>����-qǏ��ײ0�kWU�CM;I�Kc���8J�B�5��e���U9x��c4������I�Vj��I����Ē�م`�h�r�h� �I\���V�w �v��~6��Z �Bn{�>���ϞC�%#R/ YЖ��w�����n=�{�|���9>i>6��������qb-�O����}׮]�ט�A���ܣk�����}c�X=b����$RR^ (K����9K���O��J����u��l��1����qҳI��#��n�	$�!m_Gs#�N��Ƞ����T��	F/p������_�F��׬���ެaܴn������7Do�i�ֱ��}޾_�B���{���&n	�����yoo/���?�&=>��B�4�o��)�AyB]P�p<ǫ&]Lq=|7��u�,[s-��s�qѼ퐘��Î��Z�z��a:F�5h�Aj���|j����b�);��x��ꢾ�>�����AE>�*�2f���h��d�7Nަ@��$�5�R>t�9T�t��x�������)�Lwn���Øs�@���f��7^��"������M�5�L�X[��΍��W⧂Nt��^�$E����J
m�Zb5��B育�� t��a����]�~Y-��I#���)�	"�&Z�4����ӡ�x:�������S�kl�}���<&ōϸW&�KÎ(��k�cS0�3<��ں~mݺYGj+��u��p�3Dm����n���������0�����Q@�J(�{ِ���_�-�����?�F���2U��^?V����s�q�z�SuU��W��کyC������Z��֭[y�յ5j�4�g������������j�0�{l���W��}�ه��Z�߰��쑇����3�߽=㹼,K\Yd�M]���wrR�Zڇ_�X0�q)W�w�$�]P�B�1<�}2��
j2�9
�uM�v��e���B)��Z���y��ܪ��ޮ�ё� ���q��k7��uk����I~�"�|v���#a��iӦq �I�y�. ��?+ҟ6c?ڹm+��8��sU@�qߵ���Y���٭a��
t�u�d����q���� ��
��qC��B
��u�5V��"ZD�����vZ�v��f--<h�ܹ�6o�L�{.�\�����ymkp����g����wO?bM�u|�Ʀ>�X�S�Ӷm�X�ºC8�����(�-Xu�Y����M,1�S�������!�.([8���bdSL�؋����oL�������"OE�����S�"��O��T�3�R���#3Y�X����piܸqԾ��fL���i˖-�l�2E>���c����]�d�2�9��6�[#
�����2JXhU$��B@��.�s���ߡ6Mj�ES�lb�M�c��K��>p;N���Wk�ֹ����y����p�yZ}��c�^����.����_x��v(-^�����s���ǚ9�����ٳgS�"꧟��Z�=t�{�KM�h�����g�myQ�QQkk���q>z��mq�j']�=^	�^��vp��O�5���
�����r`�S��r�l��jbcS>k�����&輧��违Ni��_�;�n�B��vu�w҆�����6�f[G'w����q-�x��#��{ｏ{�1Z��H:餓��h�F���u��fE�5����8���qL�����5^?Z�%�f4}������q; �6l�i��`چ렮����Қ5k��f�8Э�~DͯO	F��/��"����48<@{v���+_�w��j�o�{��4����5������Y���}�"��a���K��Z�`v��̏uĶ����ߋ�5u����YzԪ�έ��5AyC]P�p}���GC���G��?���Ѥn�`�<���ݹlNi�M�������������$1i�jV�9s�6E�^�A�۲u�Y���ް��t5e����|���Aڽ���>�h�?.�J�����o3�_��6���ÃA�x�5vH1�;�Jvd��a����/��9�qsU�X�6�f*��}���Smm=���^��|��-���k�j����*E©L��IS�|�Ѷ���h�����4{΁��OR�$������U�_�O|�cю5jmm����������|a���^^��,��c����0��ߌ��.�7���/�g��f�����mR���h��.���9�e6�� ����Fi��RV؎��4N�����Î���LW���$�'��{hO� -Yz}�+_Q�imq͚�t�e����+i�ʗ�.��閖&GC�U���Li�Tʣ��G��gf��>�ӱ=;��>�p�h>��nq{�c�ݤ��.a��z <oƌ��o���N���J�����+mٱ�v)g��)�U���ٳ�����ϘI���9�3��-�4{�<z���8^�m���&}��ߡ�����ӭ��N�{����	�z��E�c}�vnK̚�>u�4�3E�u�	Kt}�o)��~��#�%���
_i�����z)_p�����E�M0W����rY�'>bR�������p�N{��z�z��X��M��wC�y��4o�ڭ�ͅ-�%������_���x�m�9c?��_p�Et���ӳ�?K���:��w���.����wSs��ʕ�K�n�~��0k��<�^����x��"���E������5K!���jSAw�T	>gR:��Ii�E�Ҹ�m�A7�p�t�M�܊��;���p�I�~�f�6m�J�����/��4]��+���m��;0H�W��s>�a�j\y��2~�����i�&���[o�E���V������tvv�~L�تZ�+���I�-��"�^�X��B�rl��t�%��69�u��c��c� MT<�8a2�|�-�ګo������G���F&�M����o�M�~8������VRG�.ڳ����_@�����t��n��Τ�l�������3��>�%��O�o}�
�;g-]����z�甆��_W_����	fl�4_r� ������Q>�v�<K�kf�d�:`��&g�0� N�<�n����o~C/^��˗�f}�eߠ�s��������&�؁��f#���9��6m�L���g�C�K<x?}��O��=ʾ�:Z�q3tw�6�Ϟs �w������azG�"���Ȏ�́z��~�S����YI���u���A�C]P�H�gl�zк��mF��f�i���=��|Ǻ�Y:Hm�EN@�#���U��-���h��I������Ѷm���2�N{����}�N=�t:��#8�����2U5�=L��]s��3J�<H�8���B˗/�����������E�꼆��UD�ޣ4Q\�u�M���W7�y&G�k��8�5��'�J-`|��*`眇�u�f3a��d�d_U�P�"�/��y�1z�ҬYs�܆��_�2}泟�K.��n����v���A�4�[��x�a�5w.�	���K�̥��]t�Ygѳ�Dw��G:d�2ԕ�+^��&t�8��u�}4��)-}���%�I���Ĝ�t�4�<�.��q \gB]q���Iښ��!�.(W�|ǩrF���&�h`W$��2C��]����F��?�3Ϯ@8����'�d����Z�~}�џp�	t��ߢ#�ZN�֭���=�x�b.G���Mg�}6�z�t��)S�˿F�f9s�jSB��7�L���?km����aMz��A{�k���ѸI;���~����玦��1�~{]�)h!k��]|)s̱tÍ7�W��U���n��=��l������A�HR�m��}�_��N�@/����������˖��<ʙ���-���N��F��,��� u���hy������@?�M�o�����YY��w�6J����&(s������8�K	���a~��i�D�����ҵ�W�Zæ��~��4�B��.]������h$��q-��?8�AX���;�<z��G�w<��9��Ң����߸�r&��	~�_�7�\Guu\i��E�h�kk9��sn�����Aj����hvvT����9������u)ކ����iA��~p�剓X�eì#���4�]���Mۗ���*ڲu;["�L�J�_=͞;�����j냺��'O[6m���q��իi���7m��x��Gih`�s�'�o���tݵ�`�{vh������9sf�%kUW[������ �z�(
4�&H@v́�w��(��K�R�J����\���!�s�Y��g6�����!J���D���:����FM��1��D��!�z\c�Ҷ7Rg�.jhP$������ͻ�:���]�_�ΞE6l�u���s�:�s�QZ�G?�Q̱_����q��Ս�!N�Q��{;--�_��*�Jh���%�N���uI�\>G=�}��ߦs�9�~��+�K_�k�s������͜9�ρ+`p����L������Fh��sm޸	�p������{*M�:M	)�R]U5�w��F6��T�qQn�S[�c�&���ݘ�]d���ߌ��B悲���\�y�)0Ir��'l��#�̤���ܚ�ҁv��A�[n����|�{?�ǫc��Ii�m�;��u<����;،;AwC]�c565RMc-5��smr�t��uk���ϟ�4�^�W��{7mؼ�|0g���p<z��ЄmZ��jj��~�A�;�h�+���.
J�T��-��k�N=恡|��o𜯻�:Z�v-�q�mt��>���M��?��	{h���q��L'��9�w�7��OK�-�t�):�S���f��k�L���1�����	�Л��yC 0�^���[�xm�)�&;͏����\P�B�+P).׸�4��8�������@����o骫���Ͽ�N~�{���ESg̠��qJs�C�t5+������.Z|�"�4+�o����8�-ZD�=�4i�$����XkϤ��ϡ7^{����K/qmx�W��9j��������">l;J�v)$���6Ap�v�a�y$� ��a���w|ۯ��&�-�0���W7ҏ~�#vM�����g�N�r�������7^er�2��k�������rJ��:Ϛ5�K���~��SO�u[['r�x�Ց{><�K=]=�z�J:h��6���4���L!p�F��x��o87n�V���hSX]P�B�)���a���1�}2�ۤ�=�S~-]z��&Y�.ҧv��A�u54�aB�3�@�D�NWs��֖V��wӤ}&���-��Q7��]��;��)n0��ôq�z�ZO<��4e�D��v�5WS��@����,$�斪CC�]��S����<�C]�Q�#%d��Y�xx{���G���H��G�Z1i�d��c
��a��ԧ>E����t���<�5�\��.E��|���WSW�VZ�z=��
jQ���)����z��{hB�$ʎQks��f���R����d�ܭ���hS�`mt�Zt�3n���[�r?��s�71
��&��4"��e!tA��E�Z&���$}%+7�*��|��\{�r����?��;���$����[���E�@omo��-K�n�B���`�ڶm��2[i��멣��N<�D�������E3f|�Z��hӦ���SO���9�������X���u�Uݿېh:md��S4︶�d��g*lź�k�!m�3�D�Jxx�?������s�wT߃y����N?�t>�V(� �|�:�(��e�p��7�(��G���sU���;�kJ�~�	J����ݝ��C�L�64�F3O9�lM�p-��0��'B+��]P�B�)E��t�DL�]PF���Z�l�p
�y�6��6>��\��r���Y����O�]��E��v��S�ءe��V<���-Y�ĵ���v�j甶i�����m{���|'W*�����3��R$~��7�o���j�Ny�I�?Fc4��՝�r�Q^i���R�5>;A@��ƌ�iT.K��X���ߑ��o�����9TSU�Ƭ4W�I����]��Ӵ�gbŉ[����M��~�rW�짖qM�A	5�W?}���T�z�x1u���jr/��CC#�t5/J�Θ�����}�+A�e\�Z���s��Q��_mO�8�}�[�v�ߢ��>���g�B$��B;���}ccF���mU���YAp�h5�~7��әt�O (C����:'3�1O��$��ύ�������曊Djh��m���fE���Z�iR;��`/4�����%C;�m���-|,R���<E)|���?p�ܧ����+h|�8�Oi��m�b�Wd=44��ȎD��֦`�+����]�71q�zb�6���9�ގ�#k��)\M*.,��>%!��A��U\|�3Π�^}�U��OQ$�8���V�o��q��zDH�;l�!��ֵ(��kp傪u8�衞`�u������* ��a�p��X ��`b�\�f6Nq�	��B���0ݏ�}&���2���L�G����u,��y�t饗rA�6�?��2�0������NP:�� �z�U�|e5
"�1�o}�[�U����6�SB ����f��@X�����e@_w�r��t'����d�NLr_ď�<����>��0q2����#���9�VO��u�Qgw��J�G��Y���  �jz/�����Ӷ�;8�}�������K/>��x�v�&�3��(;��'W�q0��0V�>���Q��x�X='6�S������\��cDkB�)���&F���r�\�#��ut	;Ui��{.͛��{v�{�~]Ŋ/s�Z*��NEF�v^���J��v2G4T�C�7���?��ښzT�QZe/��M��/��M�ոvl��
PK��}�)[�:��v��I�瞸���t��ﾜg�żw+!i��	l^G!�ޢ>|舊߱��cZZ���W��1z��cwg724uh�pIຸ>H���&�s��o��u��/Ƅ�Ca&6~��Y)�۲xHaA�C]P��{6d��T��?|b'i�IDŵ�<�s���.j �"���V.U
Rho�E�4w�l�Q����V$4��::��g��u��Ns��c-uժU\�DI�h�b:���~{�����T_�|�3�"��������J��]��mj�'E���k=�?�>��"�
`���d�x�n�M5R�����4����)����[�c�.�g�tn�
q�?�<_����ɼ������* �8�n��6.	{�O~��gK7���|c+o�	9@/S4��:[P�̻�X_4tA�C]P�p�h�10�C:,"b����;�Q�>���Ѡ"��q�L �j8?��s�١�#@�Tr��0���
��8h� t�ʛ"����.�;��#���
E|�RZd=M�89�ٞ
	݌3�'^j��o� cײ�_���d���x���n��M�>��<�H����д}��/�o�9 S<���p;�Ď�#��0��3E�9�EpL�r�w�G�n��������ߥ���Ў�iٲel�G�7��ϲ���"���Ot}̼mB��A]P�p���O�̈́��"��TF��L0�6�{�������7PUM5�h����h�
�7��m���7�З,Y�%����-�hɢ��'�dV~��W��/��vP��J	0�:��-�#I���|�v'6c�7�y�'���V������p���g�\����CxA������\@O��i�����W��}/�sm��Y�d����υd��- ����8���~@7��M]~�����?�y�����&OO����d�5je����uZ�L��a	)��AA8���!�.(W�:3��,��؄��6�fh������~�}���ϟ?�q��v�Ls��������h�	m�e�]�>��DO<�8�{F�����}��&M����fϚ�%ams�����T ncr7p,<R�%f�-ح�v��?߳����#�Qҵ�����x=>�ϰ�~q��Wk ���d-��z�)��g?ǂ*�A�?��9W���ϧm۷pa��������Ju�}���y:#Rd^�U��֭s�)X?�R��8N�B�c�t�s!H=wAyC]P��7��B�qr�{.��~� 8���s�D~k���_ �K/��}����tv�Vx�%�v��׹�\�h@N(�r���
s0�T�>e�IԱ���}�Y��T)-}�����)�D�}�V.FsЂ�z�N���j)��&�t
�]9~!=���AD\����$ܰ��n��4X����&�&:�#�b*%R�쵍������g�\ٮa\}����ϯ������o�Qˏ�?��O����ߍ��u�=4Ч����}M�8�	�q�;R�~~�U�q��=�ͣM6�E\H�(� �>�%�������������3sdW��)��~D�6�nv|N�B�5��e
���ݱt�_�%Dm��j@��,���lE�g��L����Na�=�]��oRo_�V��͍��m;���}���k賟�g��Hg��t�̙�l	R�^�k����ϙK�[[��r�>�J@����0ڤ6��텙���Q�3keF���B�F�:"���1��zǑ����9��֭}��.]���O>�$�y�����+G�#M�]:������7��:�}�=���N���{�'%t���:n�Z]�a���'~���##=`@�~]o���#�'T�sI]P�B�%ԃ5��#�Q�i`N�����ƅ�<?��ɀ�T ����kW;�z�{�F���&�gby��8��������?�ڱc�_�z%~�4<�O�Z��1G-��o�I��}�"�i�{O�����w����p҉T]�s���ka�������!�F��n�h�E�ē����UUTzu5Z�ꔽ�==��O�w�A�<�{�ٴj�j�޽�]?����?Gx mx�mj������~�z�q�3��>�쫗њU�p�뮻�V*	��?x�8���PϚ� I�mi(n`S����;B���F]P�B�+\.7�'z�H�g���2��NS����������L�Ą����>������[����~z�\�����R$���8�p.{���un����c�n����5���N�ҦHc�w�i�7���׉��痴,��w�������w������S�%�H�R���8ns�;97�����ؾ��/��1	w�u����&�7l��￟����Q���=b\���.��":M�굣�KUƥ��Zi���^}|��:ޠ�R1Mmt��|� ä�q��_P�@P�B�+�v���f�c.hUn�m���u����2��
cH�:Ei�L'?O�c��g����վe�f������n��N;��ܐ��~�}&yE���w��H~��=��,^D�w�`m�:���k7H��6��=Z��X�B���D���w��zդ�ip�]j���M�[���y1�{�}���;���Y:餓薛n���:��������uj=sԳ����	�O��1��]|�EJK���G?�/�Kt��ҥ�9%�*�a�H7Z���+��mz/����E�B(]P�B�)�GM�1:P�s�;xv�ʅT7�a�����q��Ft:��q�?y=���p�B�������@ ��կ�C:�r�s�"!��L�2�Z��u�x:����e���c�� @K�Ҥ�Fn�kG���4�͔>����p�$f��պ����Pv����3���O|�:� ������ﾛ��h����/�y��+�QsK�<�l�DkW�����/���c�;�^��������� ӱ.Y�䞄�k��JD�AAYB]P��kG0ˢ�[q��N�]B��;�%�Js�6�(�Fi�H�z��ǩ����l�H�����E֛�m�Nj�/]��6�_O���f�����Id�똔�u}���|3T�D�F����������G�RD��X69&�mk�v���eiЋD��ݸ~-�?�;�t�{N� C����{{����:h����/���7q���y�i��z�*%T}R��C��귨���K��cYX׵�{���]�s|��	��B�rF�T��Ñ/VJ�rV(4���xAsq��dqa��s�E�/ZHs����?��Y|!U��m�z�;�]T_W��B��5� �<a"�͜ٳ�G���Ñ��/WDmԤ1񡥩�O$\�e�4G���
o����m���s�Ɩ�(��UUU�k����CGP"4u�AA�Gz��S���o��-_~$��w�ĉ��#�����h��O�Q��]�����_��F���*!)���bJ�/��q-`�N^]P�B�+��u�P������[�j���`w@f87�߹����5�b<lWg�����]���J�θiz���t*C=��O|��Ա���LHA1�]�mt���h��B�=��ή�<�Lu��9��g%�t*��󊄼 �,�����@J)��6*�qK�p|z]0�jun6?BF���RJP���~�\�=�M�q/���s\Q��ب�������S>�s�Ӯ�vy`<n�5�ג���U맅�4KK�."5:��㙜׬^I��z
}����j#�a����,l����L�P��i���sB�����f��:I����rZ�D��B��DP ����rT*"[����V��}�G�n�55E���<7��0O�2���P2d�����cF���#�n�YF̽1u� �Be4�;�).71���XZ�i��l]Z��3�흎D����^�k8����j�j�1(��ώ�`N�=7-P�����B�۷#��������dM�I$u��|!sA�C]P�p(!g��\����:E;���~�8lڛ����h��!��#Z��8 �s�o��[t߼o���>�Jkݎ�ן��X�rM	�@�HX ���~d����ln6$k���/h��w��T�����uz>k�.�i�	���!	��86��u�!$a�p���V-vwg0z���d�	�C�/���,�t]�]�KDө�>�+)��~�ۑ� r���"�ض��mC̥*������iA�P~o�o����Ņkb�����W����1���R9d4eL�c�6��s\�kg,˂��7��K�_����8.E俠�nrP\�|�^�WL���,�s�Z��<b���r�m���Q'�߆>/��ͻ!I�x���$QHZ$�f�Ni񴩽"t�,iP�΅iZ}��|�7w����K깤��x)�@R���^X5�	<���6[3�d^�X�	�/֪:Vl����"��a�
�����N��a	nZ�j��M��A��̀�q6�%`��1�� �/�ﭔ(�A]P�pt�3�1x���v�͵���x[V�����7)Y�L���k����J؎fY�Gl��lC��xPf_{�k�v�ĵE���$
2H�FX��9.���m�� v ����_j�����fn/]ֶp~�:�B�rŘ�>�DTd.v�bE-F~�4 �Ґ�]��.�j���{4�ѭ��,�5<k_��
`:��.�����a��P��������ކ5��\?I;/-�|��BP��M�f_t�c��y���?���#��e
s�����j���1*zr14Q�nZ��(r��}m��X��$�|r���$M;�g6�Q�I����"�nP@ͷ{���(��7)h�����\Lv��tl��Х1��}����Ց��B育�҄9;Ԫ,����a�u!���Z�9v?tc�6��8��A�F;7$d����"�I�\_�qA�צ���rt��)�I�D��rG;�^���UU���ڟg�8��=��A��w݉���4p{}3&���b�$*,���F::��exS�����GK�3�� `���7��5�mL��7����H��t�p�@P�B�%؇�^F�t�h�p���S�Da��yh�������ln������Fh����!�T�:���1_�]��$
���h��~�9�:0c�����g8��R�4qA��ǖ
Ki���oR�F�@[8�Jv�a2
������^/�
���#�Ct^����Ni��@PB�%�'��m�b�y�cR��h	t2�K�Z�&��'Y�@�Ҏ~鱸��cGvC���HAb�����im�k�����W����A��m�422�����	�
������ه�y@��-��Ԋm9щj�b�CP������1�ed�0t��M#kg�^3m�7#^ԒsY�I8}�:�Y�r#����?�?B��D�9�&e�˺�M�~x��m��IAhI�ak�q��!��kD������oB�r��O{i���ܣ@�qm��g��v���gԨ�t]h(c�b�b"��<sߋeDL�N �D-��T*}-�~��*2ۖ��0���{�α����M(A�vxح%���!�.(S�� �*�/2�|����D�W���)�j�\5�$~��(��/��ſ7c��㪝9?E�r����	��>�e��S�K�1� k��GM�8&��;B�*B	U��@���e��3�Oŭ�A�x���)T�S#��Jo�(a�-��MO���\jƫ-Ź����Ok�Z�w��3ڷ��u>|�z������/���:0/��g�5�y)(k���,��݊y�ѝE�)E��Pm-��1�64S��m��ۥ}�溑��{@k�kǱy�$$��1h��u�L�h��	: ո�ߌ�������碪�I��f*�%Mi�A��}=�ej���m��Ag�u�}�Y;R	��4ћ`<'���clE���sy��G�-b��#���5�X�`��lx�-97嶫���@P�B�%'�U=SW)�����ϥ}]E��ʮy'Di�;o�����8���V<� )�(d6ZP]��n�ʹ BM@�\>���э��>��˃��R�����ݻ3�^i#� U�BͰ����"���RT����B�͍�qԶ)cj����>b��ƍ����o ��Uǃ�"� ԰_ߏ�P1��2�@A�l��mH�q�&��#��s�d�܇jkkw�@P�B�%jj�����==}+��[<��*b�R4�Q�ڔ�jS�!�Q��\�r=EX��Vt�q3)5���U�#l�.�|���v0g{�㫓�W�w}�����r�u����j/�n^=��qiuz��G�h�wS�gf���i��|\��E]��e]t<�ϩ{q�{:�˧q�9?�x9�,�uu55�t&�e��EB�H.�f�F�b�)�w�%5S������v0~Ŧ������:�shx�y㭷곹�RVSNX�E�V6��`P��r2�]�Q$�rԔݖ��tsKKS}mm�PV�bp0��1�p#�G���:2B�]"�F�V5�7��8(#�:J��Sݻ{�������JUg2~�K�|���h4-�1+�i��:�If��'ɥ���˨�|��J��]u5x���r���|*�"�)/���(_�?�L-$"��?-6��:��繍��}J�o�I׮nh����h育���,���ٯ{���JCT<���:i�#�5z����������0�^�簶��RC5DՃ����a������ju�A����ʧ��
��1(n�������)mW��e��U���M�C���T��*�/�dy?�K���pjxx$�U�8�v(?���|h�}}}�����AkU�J��S���n�j07T]��q�������^���̜3��䓏ڳv�.G��t�I����C遴�_+&��D���s��:��F��Xc>/�J;خ���cq��܈���r~~8���~]�H��#u~CCޯ��?������R�7�V?c��300���Nq�˕�]%�բP����v��w0��W��Z߯	��}����Y�C��ޫ�U���������\�1.�m�oe��������t���NA�C]P��� ����@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * B��@ T ���@ � ��@PB�� �.A@] �
��@  !t�@ * �K�U�'��4    IEND�B`�PK
     uK\z?�A�  �  /   images/a652ce68-b987-46e6-8408-d5645582d4d7.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  4IDATx��]i���U~�o����g�v�;q���&MBq�4�ԨiԪ�B%�����*!�?E��@�PA���NJ��8�K��Nl��5�Ş���[^�9��ݹ��_��f�}=��o��s޳<gy��MZW�)�uF�Yg�)�uF�Yg�)�uF�Yg�)�uF�Yg�)�uF�Yg�)�uF�dqaJi
��@O����8ؾ};�4A�$r̡�����T*�K�����!C�g��A���Pm������£G�����?@@绮G���G��bdd,W~�*���ETkc8}�MLo�3����b�5�;�~���C�){�n4[�Z���\�;JŎ���']�<�Q��D�m����</)���z1���H���b7)�I�!i�}׿X>�I�yS��<sׯ`tb�����4j:���p\guq��y:�ѩV��I��j�\ڢX:EJ�f��-
�K7HI�i�vj�R7���^B:͈����UՑ���曑jF贻�+�돑��9S�i��(J�'���Հ�6\��4���#MU�:�u��m��/����H8qDL֊$Rt<��y�L����Eӱ�L�x�J�Nwѱ�-�T'p��H�)���
�1FF0���',,y���H0�����\��as/y�����'�.�&mQ�!|=���d����I�
�''ۋ�n��f�b���c����U��&��iK%X�a �n����C�G��R�Y���ҍ%U0::*�\`�5���n��*�t��.����c�p��u�r�G��2��ׯcz|O�IP���"4�=�GB�ۿ��'&0;{�B���vᓏ>�(�\-�'2W�K�
�-��!����l�n�\����g�w�~4{=b��|�-��>}�ng;h��ڡp���W0La���4Ƨ��ڕk��}	{������[�*���G�
DQ�eL�J3���p֜w�l[<���	���+�1���&��Z dL��_����1<��c�5;x��+M\�|cS��RfjE�����w$
"6F0�(�s����E����k�nax��*��ؗ���Z�Šϊ�o���l�p��>tVZM\�p� @X�l�:|��ô���=��E��X-��1ONM�R.�҅hu��8;����)~�7~�"��Ce�|�DS0PQ4F�߻g��������hw0��yB�[q`�~�>������y��ѝ��P�K�'q��86��(�bl�����߇��e��]��x����ɇ?�{V+�,��/n�$&��K�
KK�x��c��4�{>��g�	�t���X�`�Lׁ��9�Ur2+�h�R\�!��{�݋P�7������pzC �B�������ÒЊA��|������X(��3P�i�X	�t�D��V��/���c��i�[���h�$��z]���G�ti��7���V����99>&]�ӕk�dcFZ$�;B�<(�loj��u�Ƈ�p8��iM .�8�r����]���)%�R^_Yt_(��℮'��Bp8��0 �(�R�;��bH�Y�$k]�XT���@-Z�Sm$���_eQZv;x����]QDR�t9���q��X��MR�
�Oid�H�U��3�!L�F�8t�׉f��1���2S�2����e�2+0N��	m~���<FG&��*������i��c���)�#�W�5�jǠ64��d��bɞ���~���ϗ{���o�zх��."O�U ;w��8��)pdp�YY3QEJ4��\v�L���S���	e �2u���$�H���[zȑrH��������}oVa�(d�1H�~� ~��k?���z�n���$�z�dȑr���c@H��1�3�TV7/pO�u��t�;4&�t�X��yfM���V��yY��%�8�q���|S'qj~�H�TGzy�X(��D]�0D�l"Zm��c���]�|wV�2�m�k�8�Z�A���uR�38�WC�I��ΏO`�{� &��^�>T7B�ǰ��e$��c���y�����`{[����Ze��֒�Ʊ K�ŒK%vSXC�[�A">�d�JO<�ґ��>��s~�wl��鳘<�I4�]�K�4�����B��:!-��_���1���U�Q�u$�Ļ�Ң(��~�s�7_�X�wn�}GM����'1��ǑD)�#���
/^2a܏��x���S�oz�&�MBG�� ����O�cX�׀��걦7��X�h�o��;U���)�|k�d$����D�� S�'����mw�V�v"굁r��=�N���g>��A.�1gɴ���J�����_��G���jY��`���ő
�T�]WϷ��ԓ���"g�~x�*��*�2b�d1�G�(V
R��:(�K��1._��ɉq,�,c׮�s��(�!��u��b��(1�q�&��%��u�7���ҟ#;�u(�q29�'wJ�g�a)YF�pJ�<�^����T�t���p��-6M�
dۄ�9�+�&��ǣd�v�e���ٳ�9���{�\"��;���"���o�&oiO���.����jR��:��Ą�����Y(��؍0斗��;�ro!n�8�m��������I�DrO.�a�K�喠�g~��{���zKm�߾���E:XZ^Ɛ&F��l�T*6�H�<�������~�u������~�
��!�8� �|(߮.6��� ƴ����~�ї~��R�����  ���4:i@����$wE�.GWQ"�����#�����Hc���#[�3
�&�����7n�WBR��$Bϧj��꧞�Ji�\�����Z099�ETl����0������W>�	b�"���UT��Z-G3-÷�CC��D�L���e;G"�RXJM+�X�<�ȹ/,.���d>D�2��o�� �I`i���Z�-��y���a�ڐ؞�& �?)g��������+k�\�Ţt22%Yu�N����)р4���~��&a�"�����ziJ��$3�6�d��}.����t�Tg���զ̌HWEE=�\t�&,e5T���R�&�*��&펏��H�NN9$T�9�B8��u�d/��Щ��G����Q�T�!��g+�?XC/�B��)�#ힴ�pQ+K�˹�����*|�
	��gz�,�7��A���@��G�w�a��e3v �NĤ�[�͉���;;;�}����˴#��h�����"�J%,..H�=���������������͇��v��a�a1i�@�i�9������C[^���3@�w�"h6��耵NK~;ZC�0���������#���N=r��L�f�Na~~�~%r��s��EM�s���c��x:�ۊ�M������P̏�������)�j��2�\�V�h���P�NG�Ukزm�`�[l��=ih���� t?�%\����@e )�;��eـUW�%�Ke{@�l���Egf�63��OML�����F�2���/��(�㑥^ `�O�ȸ�-�Ҽh��s�|5�����[��J�iKEI�[��nl��,(V����G=n���L�"`�fqґ��׀����R�&�/P����cき���C�l�8aX$SR���w�޿��F�l>�\<�N���	����
��/��Tޠ�\[/��D�������y5�1er��:}'%9uߎ#�ST��٧���^�,���=�(��<)���L�CLt���V�]@�ŗ�� ����U�@��kL{��dwcZ�K7�P��I8^�����F)�I�em(fB�ԪѮC�s�Ld��F	��#oɹ�'��]c�"tN���<�<a��6�����d�J�ٛ�{P=�+�KpI 9��a?�g`z+JQ(;}�'1�Č�y���o�'K�W�|��fsZ��L�_���pC�c'uen���j�	��V�B[?�R�����@���q�p �D2W�}n��v$��ӰS���C���'-l�-^���ʄ/r��SI�C�1q���Z<75��+�;�9;���BH������D"wD�P�F�+�r�l�!i���^1d�7��M�ч�Ut��!1г�|��&ELZTM�Ypq+V���,���p����� �d�ix����54V��5��K�E���ۗŌ���y&�!n���Wlr��;�Z��]T���<��HM�}W�2���'�G/F�LV�|�uE���>!36,�KQ�pJѵ�n(�̇r�|Fہ(BĔ���0��j��a�!,�����Kl�b��3��(�3��������|:7%���w()+I�;"�^�'�H�t��NBy�$g�e��������Q�;��4�9w�k�RfVR�n�py�4I��I ��CS�I&f�L��V���	q�lR�|��e����I��_Ed�TΛ��ԥc�u��_si	so�B��_�z�(m0��^�#1`�TF��%���_����G�P���7Ϝ�h���	�h�*,�4���D��,���C��^1M72R�8��q�gN���ob��w��P;���#���5�,���3��Nq��}AV�/WĔv&ıͽl��a!�����|��Q}�I���WWJ�j�T�
�P.!,u}iE�]�����Ey��U�O���}M�,��.�Yo;��$K�+��ٰ�v�K�#kI��h2q�(��f�}F��)���*�WI��<)W�Ð�t}aI�N��)��0�9s%M�̬��$*iRٟ��iG�U���
��J��\DBЍ�S�C-�E���~Y���Fu��tt���Q{��}��a�ӟH���d�C%�c�M�2	��Mw
g�����>9qN:J��8�,);I�[���G�'x��b��2YR%��j��|)�x[��3m�ʢم�\��X2�X�|�NHB(��e���yR���'9v)�B4=�92uA��Pa��L�y�(��].+�2��Bp�F�<�ڗH+ !�dS�<���h����A3�0��"]��Ou�C��#ЊM�=��}/�T��h�nÇ(
�2'f�\I"����E\_IcB���M#d=��q�pdE��R��+�&���R��L�����:�nb'E��mE�8�E�$Q��8�EHu����R	���\���V�Z-�m�mF�c�5�������GYy�DW�dMe�'�*=/�Z��\Wt�|��fv" LS�>��\V�f�70R�A�~h���/�LK��Ï>���9���s
�����i�L��c���Hɒ�S��Q��sN�T�­Z���f����O�T�}�kR*^Vλ�x�a#�NxŞz�M2�w	���67G'���'�c��v11��ݵ�) ��7���"�]q�Q�-��l�&F��-�r ���rU�ӵ����^�p6q����{K79�JCw�����=�	E�;e��5�JJ�FZ��Z�C�ּ�V�F�[b�ӧHNQtej#���^'�ju���E�eyR����p��31��c2�\��+|~��>*n��9w"��N��6�Sq�G�_
�f����x�F-�;B�M���Hqw
�}�I�@EL-d}� y8f�p�oRÝ�|΍�7(6M�sQ�f� 6}d�$|fa(O�kӴ�ި�T)�F�Ѣ�kn~ӓ��s����.���M���@���m(�&�'#�g�^�O�<�3g���]p��~�s�!\��.��Isf~"�=�t��l���E��?�ŋ��v�*����{#�!7�1�u���˧潫�P������n�l��6������1��{/�-�D��w���{���4\s+iJ��r�FO��)$�?���y���*T1������_��_�]�T�Q~P0m���rΔ�@��Lq��D��?y��;���A�2���y��X�C�܋N�����8�'Q_��q�z��3��3�}
{���r����e�x��z�2��G�S[aX�� �?ȟ��L�J��?��	D�󋋄\Hcc#��WWW���O�M(4��d���C�c6c�jf�c�V��cRb�EP�)��d��m���!�~�|)皺-u����W�DX����vW�}���*�u|⡇q׾a<7F8&��p�0��f��YB����Y����0�(ľ�{�Ν�d:�_A����Pܩs�jўgr�f�^n��C�jn�N�Cg_q��Y<����ѣ���u�ֱ�^��{62�x�O⇯���_}��p�<���G1ON]4C�]�oݯ<7��dI�B���l�e�<�<��C�,�F��)�CrN�=X�S�+ܱU��[���
x�3���G���jt���i!��Y(zm�0g�7ubG���d����	E��gbbLL�M�s+��;h���v�D8	�3z߶u��9�0�QID���wȋr���$��s����b��Lk�H�jO���|�DKi���O҇iS5��J��ֽ�ȁ���ZyQ;y�d1��=���Z;B��%�^�S�J�-��������x딞�[M�^_��nW�!�:��e�a��Պg�tj�͉E�z|/Gѹi/�R�9uT�u
����_,i6�[~ڥ�-��RV�5�j���y
�c���6Q�n�o�̙دSe-ILw�Z��0*_#=s<�-�M�G�=u�I�Ҧ@�m
d�Ѧ@�m
d�Ѧ@�m
d�Ѧ@�m
d�Ѧ@�m
d����О�щ�    IEND�B`�PK
     uK\�u`�) �) /   images/a27a8979-5023-407e-b6b7-e8628572ca80.png�PNG

   IHDR  '  '   CP��   	pHYs  �  ��+  ��IDATx��[�5�u���������?3�Cʶ��a"�;�DFd$D 'oɛ��ǀ� �ABbD�@#�DA �,&i�ER^�������u�ݗʺ�ꮮ����$�s��������u��Z_}kժ�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dɒ%K�,Y��dp�%K�,Y�d�R��I�,Y�dɒ�JI'Y�dɒ%K�+%�dy)qΙ��Ա]b��mi^����e������1�����s��_>���.���o������{�W࣏>�t<��O���{����gϞ��w��i���ǟ�$w�܁/^�۷o;���s9G��8��~����[�n����c��t���s���������\�1�v�����������X�}>G��L�`�A�٬��ϦE�(���,�KJ�V+ J�^�-�.�����5{{K�ǰ�,GߍY�ﵔ��ͦX�����v��v�1EUm
*l>_8,��']� <g�\Y�j̏��_k�י�lִ�k��`�7�l�@΋��'%����(����(,��t�a9��nk�XE���u}V�MY��k뺬���������f���w�tֹY�W��RZꛥt$�Uڇٷr/�'N���bw4�����0������H-wX>৿f���1מ���k������qz
pp����>��k�|�͖�hZ��� K��dp�e |�s1����ѧY|t~:��8/q�)��?��e�4�h[kZ�,QW���,�+U��qȦ\ʲ�����S����L�e�ӕP@cp���[��l��7�q�ee�VΖ8�7������m��jA�8����\���YI��Kg,���Ḉ�!��(�O߶R���S�t=_�'��k�`�H��/�	)KJ�Z�3vt]#�9����DQp�A�h.	(/�!��QFxS�n��b!|;��l����0=]�J��GREHK�r]K���BjA'��{Yh����e��Qi����Q�D�:.������^,��]�Q��)KCn�u��N2��P�7̍��u\��`�q��E��p�֖xEm��%��YK��t�}��@�uv�B,�Yn%�O�`'8��E� ��Rj,��H��=��b�jh����ͦ�k|o���Ƙ�k����V�����`]��`����;��Z�x?׶��'T��-��q]�Fi�u=k�,���(����Rx������SN{Ce~���'��=༁�7.����\[�=������'�  ��P#�[�mMhj���|�B��,��Y���?C0��w�_|�Gg�n��͒�%��,Hp�~���������������Ϗ�nVk�B��y�\�%�9�^%)E[��J�?����GJȦhQyS
�9�(�,`�@�1^���u8Z#�O6`XA�^�����c1���56)QR4�Vh�]H�t���p�t��z�c�D�8J��}��!R�F}G�`� �N��EB9Pf�c����Z��r^-��	KH]�P�fE��!
he�9>H���]bǊ�lYg��JP嘥P��\{@�i�Y���ȽQ�Vɧ�`�6:*�9�C�Xd`����9W�PF��Mw��x���Q��`@h��~�0����5R ���D+�V-�j�W$s�q�l��'7��Ք�s�<E�3�#��"}[ɏ��oˍc���k쿖�Չ�$pu�z@����^|�!`��+-��R�בPu+/���?�|Ӹ~Tv���N�%ʺ��K���<��@>U��`���O���Ni���sL�ޗG����w������{�<���۷o�DSeF�c/�|��7�7����������o����JU����j�s���'..V���^��X�����Ғ�am��֢��R�x���L��y&o����"1��0<�;�%n��zM�*@�1�����:�#��약\ϬD8q렌�
�r��x�ω����=��zX_��"�cXW���֗)�v�W5��qZx$�v�ԅ�����.4]L�ϰ�r�!zk�Ǩ��
�����������CG�f�g�Pa�^�k�I-�38�W�]��u�Ű��Ԑ3���6�v=���D�u��������{�5,#�v\�i��kݵ��3��i��F^Tl����g��Y����b����������/g�����+�|�y��R>�����LH����[�O�����+�����38|���O>�U��|z��	u� A6e8<<b�Al��[���J��  f
㕲��y�[�a ��3�<+���` ��		��=��l����h�="J��5� �8L�����W`B�z�*��F����0!�����u]����a,f򸁴"�����Tۆ
�`��+�P�����gN�I��+}/��y �l�N ���az׃��ׯ(l��m�.�7I��
 ��L�kw*�fK��v�Ee'hL L�(�����{L,�A�����΋ǟ��y6+����NOO����_|�����{�篿���d���N28�	�/|�#��|��w��w���W���o���������`��ge�f��p�$�'��L��v�L�M�P��;����{��jD8�HYo	�3�x�Iz+F�<SJ�;8�%M�[� #� ���g�2;w} ;E���m��;�D�=ˢ�q��0�d|�=���Ax���ʉ�J:�& �4@$���R���`���{ �DUC�*e6�پ���M �� M���2���<�d<b�D�c�g >�ڰ��}}�	o����cp`�:k����.�[�]����j��ɇ<g��wG�I6���p��!Hy���g�����/��W����������N����P>^����DȞ��������ַ��Ͼ�o�*��p�\'ͬ�ɐAE�p�釠��H�j�<v���*����U�`�y��������Gㆃ�����i���̘6�gu�ih�+��U0e�+�)�?�馔e<���C��_�*d�77`hP�C�o�O�ϲEB*nOx|�_��G��m�}>
ԇEsw�0Vʸ��u3�'ÚVg��YF�e.:�l���� i0��}f�6�3�y�����m�,������;f~�go
��]���# 9d޺� ��sx���ג[����e�[�>�@<lMz�O���"��'O�����~e>���������g����<� ��#�|�h����W��/��׾�_�O�����z���4+-TV�Q�>y+�E Rb��W�����u�A|�dЊ)0u����QCI�+Xd&���OҊR(�#Z9U��+W�&������҅}��=O͎|����}Lߋ�4~�k��� �O)-V3��!f:R�G,q?���b��%���� .d���h%W�M]�E)*0��s�g�����0](q�a�´1���χe����l&�ߡ)'�.~��\اa�����',C˧����JC����Y���qʗ��}�(-�;�3D�;�O��?~�w���GG��O��n!X�?���F���p���c ���������~�o�����D徤��@�ۣy�jǤ��37���lA�[��`�4��BA|S��4��?@��,p���~F&���wBe�6Cj��vj{ �. ��C恋U���7�ao^!*�I�h���o@��A����h�g1sKЎ ��+i�P��<�3�\��zE����^a�5�5�g���,;=�<�y����,�ޡ�T3���l�Ww�6}����Mu����3T� =ň)�#}� XFC�0�*f*?=���Oc�G�n��$�ӣ�^)�Ji(�K؆��BPWW-�8��E+�����LOX6�F�Y�.ְZ��x�����&�=��w�������������|������K_��'����o��gϞ��f]����L~8x�����L�V|�p�T�.׷�~�������y��z� �6u�o������E���m��R��q0𚴃i�7Rz������)P���.�,b�:�Ǭ��I�>fiR�^9��~6q[��01S�����S����KfP5�ȇ'̷�c��+'Q�T�!xH�ݘ��� �9(,#�_�N��1�+�:�2Ŝ�ҥ҄���(���>|@��!��t����ϡZU]7V(��# ���,l}�[�z�o�����k���f���FK'7T�Ŷ_��?������~�7p������FL1A�h@R�ql����*w���Ե��3^N��;��@~˿�w3x�tx��_?�qC�zAPU�¨xe���J�r]]ϘSB������,�=��&�)%�lE��q0����SNWJ��3}�(%�#���2 d���u:�y��晞覀�T=�<��%�?���IPR��R�p�;�˟��г߳8j�� p^���.!��c����[�ۆuW��ϗ�i�{���@�@|Ȳ�}3.��P�MS@8dWBvM���Gs�J��"��)�!0O,�$ʾ����S*��l�#X��{�����o���}�ۿ�3?�wL�A�����,�/}�K����;���>�w����W���^>�.U���3,��ϺY�-�`����<�A,V>����zm�-�����PQM��8���\:nKxmX�X8�ݞGJ�����Y�e�0����O����1#�ka�8ͶzH�0�y�=��D�� M��R����ަ`��0IԿg�ѹ�>K��������qS}�ZI�"&ڴ�QxM|�c!0�5m)��QX����lP������(����A���;T�\\�Y����Q^�W?��G}����~���_�#<�=�c��H���	1&�����}��_��o������]C�$���vK�����
D����4�*�P󿒆�ᬳ�g"�S(�`�A/<~v�M�|_�/����B�g��3zЩYƊP�#,#U��Y(x��D{(�5i�3�Tn��m}1��R���W�����㴱ҝ1s棌C
�(K!!k��{R���T�� ���v��'�0���AG����������<�7�u�Άi���>��$EMAϞ=�1������OY2�и�N���4GC�_����w��;���������>�;�X@�'�� !`�����o���ŗ���j}k6�Yu��P�+�+��э��陔���r,x�᠘Rr��8rJ��C�F &R
K��u}�>�g�ö�Q�0I,ͧ�����ee�2��J��xuP��c\�)p������?q��F��,y_C ��k��g��=8��,�?�W���uqF1dO��g�uߓ8��T_������g`{gꚸN1${G�Y&Wh\:99a�bR�U!p�a��,t�m\;G���?��?�ۇ�{�{��{����>��,7J28�A��[o������������ǿpppP�r?]���G��i�P����ٚ�����m�! 1@���]���Շg9X
Q��ਫ,  ��5@B��_����fӚOz�?mK�b��ǃu8��~VL[�K�����TNIN`�۞�9��n�c�ze*|�͢�R&N?)�-�,tLȰ��j3Z;�Ϯ��a�cP�/v���>���<��(�'=�5���O����q*�>�vOL2���S��2��oߴ36�KB����U��.g&����ȶa����?|�׾��ǿ�K���./1�q����=_��W?��;o�ڷ���_����m�,#B9��@�X,�K��d�P�%��5�'��<�LD�{edM?(��o8s��͐��K�zE�MR@$T�S����S���w��6��t���m{�h����M�cl*V"���2%�2f�3�FZݧ�4Y T�k{`�@�H��}����6V��6N�s�hö��S ��~�g� d;8�����(�0"�<�Su2G��z��i�w�:�N�����&����M:]>�� m<����_��7��>���}�_���1d�1������ٟ�����������o�u׶Kz�ufW�����Wt|���3�~�󠲩(M�g��g��q��%4�+�����$������PyN�WP�%<��;�~4������w(24)/y~7�ii#�ҧ��P	�/�}�5�O_��{��5�}�n�5�.���c<$�_����8�<;�,���m�.���cadsF�wQk@� ^c��1��A�ϙĚ��:PS �7�)�n{�z��xٮ!�2��>�C������)�3p�>��0�o}�����5�1)�Gߟ<y���H4@��z�)p2����ݿS���8A;���>�ٓ"����?���ӳ�_����bQX���^d)4`pdGh�X �%<x�*�?�j��t��Y���w~����%����Ht�$�ʦ����1�ݩX�0{��<4$\b������=�Ȯ�ƛ�l�G		����ë{� �z�H�w0��e�uv��/L~ۀև����A}>z0`��~l��k9M�<(�L(������L�N˓M!0Qt�ތ�m��������}JG�Y�����)�GY3�0��I�������rR�ҚqH�p/I��8^M3d����l@n
�i;x&�k�M��?��a��|�yMM)�&�?q�x7�f�C�����?��tw�܁O|�M�����5�'2��2��F����ʯ}������+�b&'��FH'7@���o�7?����]�g��,����i� Y��p���so����	�3w�^��h?LQ����/��~�	�w3�Ā��g�_�p*M�*�ʟ��0O�}�N�pt�����?�wx��9y�%����S����iIB�=ٮĽk����u���6���딞k{f+�/e�	��0��v��+�q�j�G���5 ���D����ꫛS�/Y�]�j۶g|[?��ϥ��$�a=����֭[��|� P��G��g8�����}���_�g��_�Nn�dpr��qد�k��ů����?�Ju6"dE0�6����k�O/?��B[iر�Q��ʘV��,�[v��|�:��Hq�^�&u͎��� >\Ù�X��Rh��n��1��[�w�5�����P��cj�S�H�^�2��bbf!V���س�9-+��K~a�'�L)�1���d[�R �2ύN@4a�7��ˮ2��i�O<�=t�%�X�qB�+���� +㘤��W��W�x��?;����/~����� ˵�N��̿����b����o��_ny���d�����Ç�7��%|�ⓝ�f)=�ؽ�����L*� >�����m
��R�^�k���|���:�+�[:2�@MmJ!ɵ�1��R�!x��H�D��/�v�G�_\f�\t���r.�<Z3\J�T����ܥ�w��]`L��np�W�@`��T��@Ӕl�����&"�0��N�B�ы/�I��)ڔT��ʣc���Iֿqv���&���,�^28��r|���7�ٳ���������Z�ᲭgX4#!ք��?~��m�%ǦS���m��0}o#����s�4��g���v�͏CR�̔B�R�<?��H	��5S�D�3vt��.5���2��)�@�O�[)�d�]H�0�]m���b���N�Qj?�6�R��f��Q�w���e�������]����&��@JA�.-VpB쮀�>�?�Y�~<�wI~������d����H'�\>���Ϟ=_�;ƈY&��J[���-~��W�����d�^xJ��qЭP�A�2��p�J��(��{n� %�Ц��:$۸�B��*T�����:iSFJ����u1���B��8mx.T>m~�Ec�&���y�l����w���x�Z��
x0I=a0¸n.j�K�g�|��T^�d��JwYI���F��{�}E ����x���#)�O��F7���������o#Hq�1yϝk/�\s��w�z��ׯVU=�@S&����`�| *|�e'ք"2RZbXh�B��ҏ�S�JD%�����XI&g�mRߘ��vJA�(�d�5]Y�&���8\�\�뗺���~j]������$%SJ3,7g$v�_�m�@A"���z������������|�����B�f;8�����ۮO�=��q_h��.ƺA"��P��޽�>r�r���
�yy��A 󓧧o���]@�k-�\s�ַ�}���=맩��A1���mx�-z�	���$x�9/Q���Ү�<h�N�ݑ͛6c3�J�����l���r��?�~G�0_Ovl-��/�G���y!U�������S��6�E��I�{�ۦ0��	��~e�;�6���־��I�#~Sm�Vv*��_����>!q���s��k|�T�:���b@�cU���"U�KN��G�8�J����>��zu?�x���!dpr�%��k.���ݺ�ni$XhY�l&3�\'v����e{����4ӃMjF��O���mj��f��7�v����1S!�b���2�����$��yX��^N3I��S`�2
�D�&ݴq߸���=I �q��8�3�/䔺6�_a�T���M�Y
�M}NM
������޶?oc�T�y�:�K��w�����z�MՔo���qަ����W>��[��1d�֒��5|9���{�խ�i�8%�`T���K]������Ù^4��ɰ��������ݑ�r�.A��xPV�7�_d��-=#ֺ�7�h
��J
L�
��y�(A�z۽毬��Iu�'Ð��v�J7��f��7�o�7�M<K)簝)�S��T~a�� c7�
��4���I��]X�]�p�o?!���2���y��a����ocaB ��9E���D�������v� ��ێ����N� ˵�N�����栩����\<��5���S1,~(�`J\Z���v;3%�u�Y}�O���@�^��w�P�aSr7u���N�CxyFg[}���5)��u���[�0��c`�����������D���T�/BR��J7�g��Z��.�nj�~��S��7v����n׳7��( V�cA~��gNl]7{���s�r�%��k,_�������4�R::�u�X����<=�g{��w�e�hj�9�=5�N��!ƛS�)�x���>��&˄������ݠ.�fϣ<�y�z�u�ٶs�~[�����1Sm��u}�k��aXV�1�����ނe�-H�P�����Ux}xM��!ʳMN�u��8�<L�W�L�k\�]��T[Re�@(�O\��̰��.�mGS�V���!�c�Me��[28��rx��]���=ytb��������D���>���Ǎm�ױq����T?��z���u��΍�*�
R}i���xF*���'5�Ӆiu��3�o��}�'媫;�z��+�_M?#�����gj�R��)�7�|��0�!��]v����M��5��q <��3�S�ϸ�cfS'ή��}Ɣ�_�dpr�����ՙ�Mp@�|���@��ZS�����/;�t/?>tlW�����M�10hu(xiI)�9Ѳx�<99��Vr}`�.��{J�nS��dj?G�gmX��Ǳ1L��?�b'�����]湙��U��}�Q��|����W_�p�w�~
p�e�zR`.��yX'��*��)U���MҞ&4esbq\�FXY��dpr��i��ў���	k���=��*�E��I�E~XI���v�� Jj�2uM+��&�m��ƈ��?'�t�&u��+��1#�g�y�*��tL���;uS�-���,;Vt� �14BŚ� %\��=Ry�:?��Եa=����Y�)�f*�<�3�I�O���7���?d��<-��N����18(���z,�3�	_��L��QA�0��6�Թ�@w���uJ=�(o��t�R� fM�0� �$[?l����?ɲ����,�?K�,L2l���c!s�#�����p��eL�1@�a ^X�XY��)hRP���;6���Q�2b�Y��N���b�Ri��ҧ T��w�E1{C��|������rU$��k,�jc�CݹF����r,��jJ�ƚm��Ԡ6�O��nIQջ�^��e�k.7��)_`������+�[9߱6jJ����)8��Zr�t����ͤ��
f����}-:���*D�y��u}(���zkS�G��yk�B5�
V0Q�w��Ϥv������$��}94#���p�o�{[G{��Ho&���N����v�%9,�>�v�g����W�v�Pރ�<@�Y�)`:��w��a��;�j[�ΐQ��`k\g���0��;;��xfQY��J'�XNȶj��l�����R����R;��e䆃��>��}L�~�
�r|ɱb�,��`�+�Ԑ�2t���#�fF�\���� Ř!�@��I��n�1��J�5�j�tTߖ�p��x��㝢o{5KJ��$�A�랁�Q��z�ϛ(0��6�P����w5�Aj�Æ������f���HZJ]j�w�K<iZ��>��Pd�03�G����x������Ɨ�J�S�P=0��@�79_y S��p�\4����F������P|�f�!=�c�F�1�1��O�:�^��w�2)%10��0}ƀo�� 7��àN
��fA���eYَI�~�1
č�vl��[��Nn�dpr�gǦ���ݤ������+d ��;p��'���~ 飾ҟ��NS��)�C��~�o����TL��,,u>��ƃ�إ�rF����Jΐ�$%�����M��bo+ih�f�G�\a�	N�r/�� ,�u���|�uJ`�̬��g�3 �hOJ�XO�
��ۀ��jb��3/�+1�9V�z�R��E�#¾e�P�@�%�B)���	�$Z��Z��َӠ����-�P��
�XP��AZ��%��
^O�F�"eM��&T����[����b���H�J9���d*��4��}����x�����X�B�!e�<���"��j����j9��u)�O(}��SK?�~��m�f.�Um:�,�J28��B�;����)\�pP
m��pЁ�f8�������*�����rw�/�?d�B�)� ų��<bi=P��(	�� J֙�I�1�'�Jf+xgiN����<�|���J�f�4{�0�rzU�x��j+`A�#2�xe�g�Dg���o�o� �#afA}d\/�gV�7_ul�O�2@��m�u"�S0�l�N��|�U�� aG@�mM�gӺ�
C���;S���^s/y��|�	�#M� ����HyN:����� J�M�q�/���{�KB��2�L�<�7�����S���{�a�w�&	�g�(�a���!�hK������� �� �e���3�){���pD�-�l����2�U�^��)����������0(fTy�k��nÀ�f�	�'�$��U)��x��l�����������t�� ��+7�f���* V��� �58���Zo~j�G�^�L��pR����	��j�(�o2����f�t����`��t%��쌀����
f3�J	��㒾a`栴���eF�R_�}@H�\����j=P
42Л�<�o��P0OAN�dm�MdL[�l�ޝX�+���<� b���c��w�D�����8���3ՆT�c�E��5 '�8�A'7@28��b��؝i��21��m@�ϩ�`<�N�J��I�$P�Sץ�2LtЅ� E�>>���K���
e�GQ~fi�����Jp�/�9�FN�����yv�(��,�aQ���l��g�����N���0�o˦&n?��Px�o�%��bzS�����X.�e��!�j�9�y�����dfy�l�o�c7c+>.��Ƶ�-��6K�V@J�SH�q�c�C�@�f���G
չ�똙r|m���XP0~�b�#fO�ύ�%���0��gx��떒�v�����T���γq�a�u�w�&b\�P�CV(mB����ZJ'+�A��HR��HS�SiR�����6k�̬,�������tڟK+�!�*ߠ�# �z@`Ya�S�&�W!&�ͨ�5^	R�B�
�&A	��T��i�z@u+̅�g��V@D�_��4�j�_��=^�M4~H0�D�Bq��('_Ã$
ĉ<;FF�ƻ��/	�$F���!����V�Dq�F�5��A�M�~q%�H�W6�q_�ܔ�a�0��_ �),����!��0���ʞP{Z�&&����O���:����4�m�r4�Z�*�S��#�� ��R@!E�5S������I��	߇0�N�.	Fm������)�����fH'7L.�H��1+�sq�mi4]H�N��lۻL;>���]Tpp���&�'?�È�fEmd`m�	�z3�8a��pL�(��K�ء��!�(�e%,�5#6�=�ς�� ~��#�B��{��~���b��x�P2�1k{F9
";(���L
w�f�r���zv�;��f�n7L��T�F��ہ��ι�����<,�厼_�pG;6Լ*�PA& Μ�.0
��X������փB�
�L��󠶕�Ĵ���\��`6d�R "�l霂��)IMRLF�,tY`��|���\c�K\���nXo�K��q��x3��F�����H'�X�[����LX'�p?ȥ"1� �e@IJ�(��	/;�{�l)U��Ǹ\��A~XOL��;5�3^�Z��If�G�T,t�-���s	��y��J����R�e�b�a��@K�e����i��￬��+k�aP��ot�K�`���*'���%�5���Ds}��%�M|i�dc@bYoӵ�..���FV$Ic=8`��d��J�o�s��HU�34�C+z�!?�+�p���55�4��%l�Y�L˒�c�Q� �W=;Yy�˨�>��
MC���_�؟����v{ς*S5���$���Z��	�B蒬��3|&�OM&a���3�7�[��ǐ���̴���x0Ѧ�Y3��ˌMY��dpr��e�5��6p��]�58�Ҧ@A*m�&^v�ɟu��)�kʬ3�_<��_W�8�@x`�kI�yvE��θJB�N�gt������R;��,r��v���Rd+p�0�ƈ/	�%++c�!}�f�һ�8�Qy����aPAf�R�$j�MNr��c=d����;pN�]ʢ���l��O�7��fo��Cj����Z���E@U��d�PI&/&���v�9��b�k��FV�PZ_NZo�Ƅ@��y��4�g�����PZ�ai�ƳZ���J�DJ:�Y�My�L��b/.�������J�.)�#f~��cv)�'�cj�����%H�,W\28�Ʋ\�J�JT�@��۔sj@ܶiLѦ6�igݘ-5�(cr�fO��la��lj����ˮ�s[$�H�5Y�*��4�ȭ� )X��*H��fT�3X�c���_}���yM��έ�i�XZ����S��
�{a6���P���v����b;��3��(稈�9"а>e�d��t	f惎�-ףuƯDj`F�ŉ��q���ο�~Q�U9��0����mJ|F,�� ",=/%�ô�lSz���"�5^��)�E)�̰?��,���h̠T�3ǖ�,������%ݛV�����b�&1S�7�q�R��o:kň���gA��<� Je�ϖ8��|�oG�{�?�w#|.�V���5m��e^b�j�׀��	�M�Cq{z�gl2s�^G�q�,�^28��rqqA���d�.c���.�SH,�hکYa�_�����$�Cxݥ(_���St�м$�X�-|XZ�K>V9� E;��}߮� )+~��W�-��3QĨ�e3ZalI��T���XƲ�aӮ���x�++VT���7qN�졂?1���H)��gQ��X�g0[,a����%���$�+��Q3��9/en�m��:1q8�X��a������ljf8~K+&�V�l8������4�+��Y8Z.�NI~$5<:;��]�����h����W1�\ 0:��y�`����f���g-��J�����ۇ�����\��9�ό@E�f��FY,R�)@߃1�#j:�M��9>����U�~^Ɣ+�̄S`!9a�a}���c�.g���h���D'\�l�v���xy���'˵�N����'a���_Τ�w�x�e{S�E����5�]��T�+m��@��-��^Z�_��ߣFVt���p�4C?,*xu��]2���ܠ�$e�l�F��A��bf��`��J� ����(P/�q0��s�=� и3oᖭ�l��źDP`���[�pqZ�`��A+X�&���w�>y�>'���k�{pv�
}հ�&�	�q�bR���w��>��i�-�4_3��;��ߖO701�h 4b��,l��!	���ѝEw��rO��v����!��h����p���%����V�}w�����z���<>��	���ý��ò�8�-��?X�O[8��h&%׶�����z�S�9ň�X�������]u�fJ���,���1U�.���.�1țl�3Mc20����5��b�y�g��C��S��6&!+�C]<N�"&)�b?.�Ӳ�a.�&���~��[��ȇ�_��
���P��C��
���]"0��V�Dp&��%*�G'n߁����iUm`Y.���[�e���ܛ݁e��s��&�G-�pQ��z��^y ���z�F�ʺ(<���/�]8x��j�Ϋ^��Oq�1��h樴gl�*m�N��44d*��Y�v۲�/�F��F�l��?��90k�!_G>x-��0�WC��2���n.��� ���OBA�`s��1ܺWL;~��e������3�EnY�}k=��@p�&1�#��W�T�������J����nN�g|�� �)���χ�`; R�)_��=�ߙK3z0~�����m�O�=���+gB�V��e��~����!i)B�y02�q{�7�	�)�y)�M�N�������NS��΀U���gU2��5�<vp�?���)I���1�vr!�MRg\�<�P�p���y��#,ʺ���3x��=�ώ`qt^y�M3����^�������Ã%�zt�j8��[.���9���@�R����=�><>~� b�����k���lY�a��A}G���V��x�usfs��/P��Hq^�pJ��4�a=��h��8��a�Ni�0~.l#+h�����QSS���!���ұ���=/�4��x�]l�A�q����{�`���9��ϱ.�`�}�"�����@s'���þ*�-��ڙ���|)��ɋ�C�@���+�V#G[bYZ+��o.`��s^j3���,iHq�B�+}>�)�Oyn��'�oѳ��s?�q4�]�e,����8�N�6M�(1k�!ܞ��q]��!io3'RG��d��?4˕�N���~�p���f��F�E''��K�fH�D�}8²STvw>��6�泭��.��DQ�U^v*A��.Bf�W�P̐�g�sp�=T�V� �9���������AB��"sT�����n�~���5��!�Q��;��ʓ�3�;����N؀B~-sb����)�CPs�C���G��b� � �IsR��/� ��5��lm�{Ϗx��{�ph*6U���7%<:]����+GK�_.`U;(�'�gx�����?[ � *�bw<=z��>y�^�p��ZVְ�-���e?!���V�`��!�٫g0��P"�r�%%B�%�>���GL�����>��x��,��z��iQ# *9���(��ԑ�~$��D�5���5�x����p:�~�X��s���J�˄�S�3f��������#d,���Ӹ1�
��lR�_^F� N��Y��dpr�����;���z����p���I;��o.*�.��'�M��n13��� �`NR�+Lq>=#��r���C�M�=�}�¦�R_2K��UZ���y>G�JΘ��⏸ִ����Z0�KR�8>[�k����@�R��^�d��]Z�5o�jk8^� k��V�k����%,�^��wggpn���
�9��R��p���{����]�褁%���%�=z����(=�#Z�m�WR���U���7�*�s��~�u�@0R�W��;�����.�lPIn�p���.����^9��3�2ܓ�f�����V(
�+S�P�"P+��l;4�v��!<{�}z*!�i�O0������:cf>H�]��-H�;x��Nljِ�������	��\�&��G#fc�X�0���^ە�~*���
���e����6����� 0)�]�o�dpr�e�l]!��v6X��#^�ҫ?I8�Jf����6I����b�x�l/N�hp�v�����`�;�),����d`jVF.��=�P1S�۳
�a�h���|-�7p���+h��( Ha�k�3ҬDlN�-�pR����� 몆gk�� ��-6e�)h������;`3�[_��'5��h*��a���1�bV�o���,��f׫T�5��R�Y	�JΧ-��>j��=�T��\ �Z��ݵd��ZWlʢ�8���x������[����q�@�"� �B`1��.%�/.��|��(@�5�)�3A�=��ϱN��9�N6#?8i�v�W}o�ރ;1N�!�ۇ_�Y�AX����\]/��1ؿ���I����⾤�l�W"��{���D��5ݳ浶<���?����'� �
�#q���M-S@>�W�o�vhVv&N?%a��z��O3S}�d�����5R $���Q@���$��6�8XS&bz��?c�����0�Cj�J��צּ8�0Y��7��h�����n��G?n��*%�9���hX�E�hY9�/r�<X���"EqO�V�����r����p�lZ^�B>"�j���U�f��]�sT��!8Z8[U����Q	G�l��x�⌙�"���r+fk�*q����M}�����;9������]y+�WX����%�^U�~���5���;��U�l^9]�L�Y�aү��~<�����m�"(�vn�W*���#�ϲҧ��d&B�Lm1��9��a���[�NE�@�>��^6pﰀ#r�?g�x�r{����#�Ξ3cD��4�ͬ�A�0O�z�Y���,j^~]5~wcv��A��Y�/O������[�s���$I�a]�]%*��w��e�n���#fOv��=���!d,�7��@(������A2�����d����A���q�
���:H'�Z�h6�Z	� �"�$T�����iB���-63&+�7��%���t�	�1~��*P\��c`�
�B���LB�2+���X���n�i�K�����fe�=s~~�Jxfe�[ޏ�	�~�����Fc^H�4"���U��8�zA��@|@��dV��=���G+V�U��p�c���S̫`��Zكf��s^.��t�P9ZJ\�O�&�����7�fGK8[[Rܒ��YU3�K�I&����){���|�~���A�X�igv^lj�8F`�
{FKhh��L1�5������[Ρ^,�6+nMO��m���vŀ������z�)�E����G�}q���i�V���R�82������v�f'�&�ЂW5DGXǓg�JX�C6���;���=�wp�a��04����d�4������0g'�� ��#�ڂ�5��f�a�"A�Hƃ�J�;P�Db�,�����4�ښ~�]�-���'�^4M�ip4y/t�ٿ�� v�V���� [�6~'��o~HN�m��zЀC��w��Z��ٜ�Ā%ܝX�B ֏3�@f����Y�H'�XP�:Z=�?x�>��0�U��9��կ#�ųJ��owdK��q9���f���p�\�g�2z���b	/����}�{���S�}���O�ܽsW|0Y��x%!3c�>}ݽ?��G۵�~�wO���򢥳z�9�,J������%<m���%��{p�`a�"&
��0H~ 5��;c���c~+ p�IN����V�,��^��ɳ����Z�\XZ˲���zv /��~����|�����)���h簠ȵ�b�3��**h
l���h��K(��TG�%ݵ���%*�2	a߬k��b{Kl��"%�w��{�9�92�<q0����7� �~����0ܹ{��g��r���GĶ�aU����5��I��-7ng0Gpu�u]!�B��+o���s8�(38�%L>�9�x��2�� �Q��ρ��e��~�)o�<�m�9�>|�C�+��{*����揱��w��ƹ~RC�8�Z�WU6P���>*n���r?��6c������bV%IY��dpr��|N���`0c�m����vڱ�Z�fL�N�b.SN����t2��|���� `��������o��-�p�bo)J����}G��R�� �����tŽ�S�S0�����%��+��ji�93&L�"�n�̲ɑ�bu��ܿw������˶�v����=���<��Qxf�-20[�p����f��v�噮���p��8F0��������)<|��=�����pA���{0���s8�p�{sؠ����9���-�mĬP�W�Glm@@������,ˑj��V����}0��=��ضr�gܧ��GmX���m3�\�2����C��o7�ȃ@ϝ�>X��>�Ƕ�i
CO��6U���(f0�Kx����;�#����l��7X�Za�4�/y�KEϓ-�CD�(��J=Z��P�
�����d���`�lЗ2y�M$��E�UX�2;z-��/�Q��;2c3�]�2#���};�Lʰ����&H'�X�ܞn��� 8^q�����\gq)[�p�Lۈc[tJv��󩈔�G�@6��!�:�|��[�\�IL�ӧO�q�ᛟ`�A��P,�7���)��1]���Jl�Ј��0�~'`#1"���_�G.�6��p��?1 ��e�#QRI߾8_����.��촪����7��i�b���\��{ǨtOJ�C��cu� ����ye_��Z�ˁ�l5G%^m�w�@���3�ˀk�ǝ%pD�j� ����7���O����6���f#�g{Д���8�`�Py,V�R��S�4�[��^�i52�=Y����n�3������;�$JkC����ǘ��ᅃ��G�E ��.��0�+��/P᭛��@UB��f���v�[���y��Zc?�7\P�~�gxhB��"[[	@�?S�W)�-���|��=�?�3%)02dL�w���1$��،2�����	�2e��ۭ�Lj�OML����A*˵�N�����ɇt1���J����䦛~�9�����fn�ǨL�� �1h����V���~�m{�q��6�1�x��n߿��kFo�W��6�cB��z�U��o<M��Ċk��+���)������Ȍ��`]����~ü�0l�#��8�by�9x]-�4-^S!PxRU�'@��zN�5�d��F��D���?dr�%�-��d��`�{ܷ/�7�����p{��sE����3���c�ݠ�oW�a�U#��i��
�bY�����W.�����cV�n7pV��]nN�&B���<6EU�,3ͦ���;ڼObƬ��3��R��9���F�NմG�:��jT�N#�MdΌMS��kb��5^��bË����L�g���΄# �1�͑!��=>�MCCsD�^���ޫ�;��߷��2�{& E�'��F��М�I�)�qʬ�j��#�Ӿ%����B���!��P��yV�-L��{>�lj���iI�=e������
70_q�VbR�Y��|ؠ���?�+2��N�\�����r6�)׀���=eX�����̦k"�)60߄E�Ϭ<�ox�?L�7�#����.A���~�;��9��6>��q�m14��(̍��m+���N���'�Ƕ�v*6%�D��&}� ��x����,���[0�kUm�+pJ��u�8Ce�����`=� ����v��I!U���v�7�"x$C�͆��31����K2�����˕�υ��켣�لүtO����y��{��~l� ���4e�M�|����~�N���Yq=V�M;�LOA��7��E�.��s�;�̘=h��!,��1`
�qN�����J�#�Q�U
Z�7 �7#5�	�F��4�uK�ܦq�,7E28���X�)�8��� F�FM�{v�����LɶY�63T�ݩ/���!�5bj	�eQ�Ҏ�sgٯݻ���~#�i��zv���rXr*�_g�R�?#�C@J7���F����4�^�|dh�aSB|6���)� Z�c����+>h�9*����kg����p���3YiK��Zar����>�h���f*�wA���� ���u�� ?^5� d^��ϥ��E,����lf��ocɬO%�������Ғjb��U0%�:\�zڏV��
���|Vd�����l1��e���~{ny
��H�h%�fa������(��̪Z�(�[����2��t ����N��� @�;\����7~������R��$#�W��mf�]��)���+)6%�cJ�k���9�H'�X�v����|7Y�b!@�/{8���z�sI0"Sf���@	�M]��Ùi?0�����i�Q�E�i�`iy��j�i�$�T��I݂L0�07��m�xPKyV|4j6'X��;��C�)�l��y��������B���?�9�U����G�:>>&�	s�/�@�,=�[Z�R�>5ċ�цNrз��fK�T����|���o��)�´��d�z��({Z���]z�n[_r 8�GI%�f�(�4��bm�ȟ�B�S��R�i�F�	�Kf�j�@q�՜V���bP�t-��e��0Gjrd�"�fs6m�éY���;���o��!�2��VO�ɉ��#̣(��ٜA��K�5�y�o�ݡ��Kf����h��+m��(|�b3h���dfB�E�u�l�*�=u��l4`���v�Ѥ�:M1������DI�M��m�*���9�r�%��&!�H��S��m��x �ΰ�5� ��'F�N���l4���lrq|=9)6�z�d#
��W��Z���X& J����0GeO{�P 0�"�P���!Χ�"���JaKe�7(@�@ku�MG�������B�L3�j؜`9�)���b��F%>��i}9�+*R���B=c�t&���`�t���}b�s�8�X����������8�CR$Uɣo/ա�+V����%t-������= �C� B6��ʿ��>�O}�9L_��#�H���m��=�fĈ%[�l:B��yXq��Zf��6�h4=�l!}I׶M،�7�]�ו���W�n�����]����J�������R����J��p�b5��j��m�9+�gx��9w�|Yl~�Oìa������N�������Y\5���d[Aϼ��e��x�rB�z�o8Ȅ,��7hR3��:$���n�!e�:���*�	�_�'^��f ��K�Q��2�@S�h?X�������,���dUU��-
�1BN,4��G��0&�߆�
9��?L���eJ��S�k&�[бFB�,i9�G�Q;�5��8����Ⱥ G��f�hE�Mこ�(�`ʎ�V0��FV)QZ��A���!�݊���mdՓ�`[r���2Pt���@aY������/��%PcM&��o� \NI���C�y��F{���{�Y*2���c��[�vto�()�h���`G]ʓ��[��x%�Ԝ4r.���9����ƛ���&���3������u��1��S�Z�*o ��MOF����:��$�(N����
�Rz,|��s
n�q!����L���F������p�������&H'�X��q�k���	�X���;���Ejy`�/�*�p N͎�����7E9�3(=V h���މB3��A3iRV�9*�M-��AQaY�a2졲���N�`�J�8�EI>�r�d�T��ό�H����b�@}�+t�J��4_�6ˀ�g��K���g�+G�z^8��"ֈ��2��{��F����H�݄P��>'>f�1����.�F�s4���\KA�\-�"�րW�F�VF|zԼ���{Nt�r7��MG�W�{N�H�YJW���tF'����,1�9Q�Vo�g͸.~&ι�}j���,3E��w���YV�b��O�?�"��k�R�w^��m̊����jG
²�|F���+:��0m|�;��٬s$��k,{{{��Md'3F��kPej M���IW����T)T����E=�ʠ�8��߀8�Ғ��5��oӲ�d����3���W������B��k��_6i�	R�Ӹ>8���׭�H'�_����*i'�X�fр�sX�~��3���A�S�N2������39�����jD_4���+��i� V��~6����<�+��^�.G
�S��Kp�����Y�DH`:^�ӭ�(�'�G�����ߘ�"�e��5f���6����7��}�p�K߹�k���xh��
���1��z�]�}.RϷJ�s��	G%qbe�0Ϙ�H��3e���jb�46�����If35 e�V���5���MK��i����W������КVχ�]>�i�؍�=x���xV����.�G"����V��G�f���)F��o?�EbS֕��t���Ş�H��hي��5�ۡ}���s6e`�(���8��x�ŧ�%���+a}��?FWyO���~�#l	�$�:E���iq0@�v��Z��Z�l�����6A��$6���Bi21�j&�uS�uP�HKn%W�w�`���f��j�o�W�WJ7�Դ~�#�{�{K�"_"��q�9 ���x%��/Z>~� �P9������X�:b�K�H�������@"6�\���NvKI��L��!�#�q}v���Yn�dpr���m�����%�8'N���G�O"ivcx>5p\f �3��\C��w^�6N���RV
��J紖��M�o�%�,+sx�6p�p���9-��e����)���4�(���<�v����AC��%���4B���H)�j��J	k�?�����`�^��à����pc���O�be�?Bַ�W�,�UnC��>x�H�����c<$��94��Li_9��a���;����@	sB���\��)���CӁ�Xh 1�x� tKû{���\�o�Lۊ�k���b=������ۙ�䷖�fh��v̎��>Lô}�rl���_��
���l+��xR33�-���s�r$��k,���<�Zz����x4�c-���i�!h��Á'NӺ)y3R\�^�Jdx��?q���ժ��@�=�.�G[��g����?���Z8�m�9��h�^4�t�'�.�G�H���^��N��u����\�B�f�g����;�P���d���Fo�(i������ zu��Io�0�Q
�y��J�jH2X�gҴ����r���FL7�/^6����������_%�qiZ�M2r��i=��J���{|WqP�X]Ќ�� jy�ȬN�˲e�ݦ+��o"��J��{ߙ[����0]Z���L)ߍД�b8S����N'3� 	C�G5�$��:�I�Mܮ1���?^~\�r5%��k,8X��5�u.z%�/hL���:ɩ�95Ì�</K��8h��\�*�^/I���/!+����IRe-}'S���nvOiZ޽�r�T>�8�mDy9m��l�)8^��Z�4)��֛8�|b�]���[�T�Z��}�N�� '�J �2F>���ه� ��������ϊ=(�ܱB��n�q<�q!/�s�4����\""�OL��J�Zud�ְC�1D|�|OI;�x�u}|g���ٿ��M�a��R@�eh�hi��N�Ԇ��FL����?/�]��¬��4�˚3�ӱ�նk4īvv��|�VV���,J�9�7�Sh�E���f
�-�,7_28��rr���V����7�Zp8��%�� %��WJR f�lpT�	�u7:�A�z�ϊ���,d*`�v�,XI��t�Ψe�����"ٝ�y�ځ	_Ϝ�H�)�rW�§a�a��8?S櫌�>we@�t���8h��?B��I��u��;�����β-x��{l1C1�Њ�@�k�!�|K�z$��rlUZ�ld�Q������A���˅[e��֛m<��`Ċ醁\#��з�U_�֯�RE眏꫎���j"k%�`�0�b���BK�5*�:�V�����R��H�ܕ�A�����o��<����)?���m�]��)�J��y��35ai�����D�e�u��Lɱ"c���dpr#%�?��_�8cj���?�AR�u�7,sz��^v��"a���p<�G�-��:YU��p�f��[�08��b"�!����q *�
)p�=�cl#���7��&�
�xp �%���������z�����0�B�NIw��-��wb��FU�����͖��Z]�#�Q��W)ye����q���C��?�3��U�ؠ����bs�lp�=+�<	��V���P��c<W�k@���G��o>/�$o���z�$a��>:��(P��Ű	��7ey6>F�MM�bS��،2=��2����^����,�}��Sy�c
��Nn�dpr���Ȥ8Z�,���δ�`S����fELt�E�@E�ԥ���(ǴNf�6���3�0�Cl9��j#R5,g3�w����W���fx�V�PYJ��i���|�,ʦn�-���J��,�%3�HTW�=���xeU�B�;Z�*�x������b%傳ΛW�S��+�_��s�t�i �-�fuf%�.(�3K���7KY^Y��+q�6���ȑ����A��	7ś�?�zV��Tr�	u��Fc�}R� �Z{<��B1MZ��AY�p<�r�4�JMc͘zh)>�T�u�G�U3��>�=��7�"�~�!#����L�I<1�GB�#<�	��']�G���'~���aa��i����WӌC��L<1 ��Z'Ӂ6�����uYȾ�s�A��YO�+/�\c988PG��eTE��%�DC�L(��zC����y�fG!�!�A/��|�).3��h��E�X�-�]�Pn����G��z������So�	O���B ���ࢪ6@ci?�[�������/a����s^��0�og{p���B�V3IE6���5��iGD���	j�
?���ߪ�t*Q(�ԕ��4��������i���M�;NDX!A��]4��hƃ _��.�c�0�*4�هnVܭ2��`Q����l�G�U����w�x�J<72�p�Z�3&=�1���W�=�V�� pG�-<8��	��d�{��EoEۦGCl��ø�L!)6�e$e^��<n�x���3�W�~�y�d�����5�/^�^t:aKҶ*��*����b����i�����/{\��ğa���_٬Q�/�އWރ��S8;y�y�ux��]�{pfNfnu��3�z�ެ6k�6��� ��Oa�jp����!�X���9,�ȬSye�Z���>6�Pi�n������b�+�@���;~���T)�[ B���3��,��
+A#&#k$�j��;�4a�Ɏ���2���u��M��-�<�у6�����J ϣ xsT��A������uTI�<�Z/%�����b�]M�Y%��~��\Y��7`�&&ɘj<���k�h\���e�)'.�Y3���̓����xa�>n�g�����־laY��dpr����L:��)3�)G�(�;e��t*��y�e��1��4��,+,s���h�G{KX@'/���p����/G=X�!`�r�W�вW��c����_p����� �Y�Y���X�i�Z]��l�$D��ֲD�z�-��z�������K"�ׅ��8��U�n<?��z.�.6-�g�E�X�Ԭ�υ�T� �7����Y���t�~48�� ���ꜩ�m
��>���I[���ޫ)��b�c��)��6p0Ś��Gү����[ah���fW����q;��)z��\���N��:��vzV��9�{�L�WbIQ�s��^��ˊ�����[f��*��簿�fs�^��G��(�)�b�QL�ď�<�v��0G��h����!����v�{�̼9���1���~M��o����]������q�[դ� �?>H[Ȁ���[��_~+ԇ7�xc��>�H����r�/�U�a����h�2{���`����5.0����wyS�pH����Wxl�I���;f�S Q�k��̨u��׽U�ſw!�Ҵ&�7m��U��=��
���e�%�2������b|������@�eA��'�\cy����&ݎ�8� h&�>�CUd�ή��\��M��\d��Yّ1�s�;H2c �a %�ܤ���K2�<��_��޶;;��/ס�	�+�sO*k��R	�e�z��!�>�O�� _q�#�����||��g8�1���^d�� s��Н�ˉ����������y�?����������@~Q �wɾ;HJ�����R
��\E¬�p�'m0DM�1]��>E��I��Z�a�XvC�'���Ϝ�!ȝyl�+J=��&��0���(��bp��9rb'��Ƙ�4n��D�(���(߽�n���1-��+���SE�c3ʛ9Q@�2T�rs�'�{�I{L����� ��^�6TKeӱ�#oטr�-�܍n�6pr����'����̔Lޛ���ߺ���E����a���RA/�t������{t�uZ��?��;����1�8��N���`x_&^:�[6bB[��w��9�H�dp��m`L`���!#�CGac[���ӷҹ:ѓȑ�u�����¾�5H��!1xbH
������b�� �����_�k P�3i�� 7&�
�˾K
C���$G*w�Rv�\@�+yW.b����B��(ٻ���xC~��SP ��k퐝���}~ذ[R-����,����5����z��{��$�Ym�F�G8�u*��]�Lz܏�$��\ڞ�Ԓ�[�ʵ&��]�i���޹�/ ���;�G|���#��G^4�Ey�����!��=���$����:�/�����	���3;?��vQ+5f)�R��o�(����Gaɐ�j��z@���I`&�R��Ģ�-%�[��ʉĘ���-h$,����(����C֬�Q��t� j�ۋ���U_��TS��k��*�)�H˜��Ż�>��vR���}�ٱH^v����L�xu�D���['tyZZ�0�Ә�wmڀʽ�Nn�f:�0����v��,��d�}��$1�<������p����\�@�/Юv"o�#��G�J�+�n2d�1]2��*#
��v���G��e���H�.��r.�������o�����/ &��|{0�����,�s��{�bN}�$�d�%r� &O�R���d;ȨY?���#�d�ү�Q4)�t�W��5")dҤ��eE�h����[��IU�0!-1���'&�Ҹ�&#mI~|4���z�s���g'v�������O�y�>_8�q��~�� ��<==���[
ģ.c��e���a�[��%mE+=׮����AJKk����d�{������Nn�~������<�#d��#{�Lx�FZ�Jlޅ~�v�'��*��"���4�ˀ�� �#)y:�d�@�H�̫����, �#5����бޱ|�qHi#H������tt�ޏ�p�p��3�#�W�%ILÎ8ߔ��
x������+pRI��X���C'r���	3V���g�
��M���V�c��q,�/�-�@Ț�
Vb��?f]��t�OFd�T��R	;$� ړPZ� ����f�'x�}��	��d�g���|��~������~���209.������KŘ������a%<�sCߙ�����������V�CZ��6(��b��� �� U]�u���ׯ�n�6pr��/~�����Id-i�.�-�ˏRIS<:��[�@ˢW�Hw������QS�z��2`�R���*]�ԍ��Ek��g�pX����?���eaL#|;��=��-@��m�;�p<�B{�h�Fn��cN�D��{��N�|���v�$FN�#���#�&�È��:~�'Rr����(5rQS��BV9i���1�٩��y+m��Z+"�d���+�Q��I%w�ʆ1����Ӊ�a� ���� ��կh��j����e�+BrN��rT�F0xsP.�z�1_�-a�ωl-��� �i54����w��Ӕxu�$��r�]���ۦ���n�ۥ��:��Z��[�z�om�xq�t�N�o�z)\��ٲ(1����iK��Є�t�x��)��pK����"�?�����~��NL}����<�.�KE��BZ��8d	�*
��В.��w�a>�ĳkM3\��:&��=���ϕ�?�(6�`��g��[�	~F��PS'n�b�*;ڂ� 'GV�u��_ҩ+9�#��Jk?�l�0$ݖ�vbS�H�	���B�<$�(Z gN@__���_Y@�R�N�[���N���|||���J��i�1֎�y&B�P����8���ԞCI��������=i�a�#����z>ۓa�<2O��&kГ�ߜ��	m��Ʃ�٘�2��n�
�w_\�[n1���%� fz��P�pQ�q�'2'�-�=d�Q��41/�]��(#��0���n?.f��;|����������㯟���=|��>�DR2z��E�T�k�kc��3� �E������:E�������1����Bc�v�~�ϰ����^"��/����_�����F��}��P�n��T7�� ���@��ɭ�#*˶�l)�{x�!oYa{��G��
����~&'� Vj�N��#0���<>=,���|{���w@;$�����t�OW�LE{����ʥ~G�-ekv�m��˛�zn{��y[���.������w��zV_f8��F�ˮ��9a����Ħ���A��k���T��ݳ'鑷�\���h��^�����B�i!FL+&�EG��=��M9I�b��*�1I�S���o�ay�� �?f�P��D����G��o~��>���N��������XZE�ӜꝘ$&�m\����ErL�����Ƅ���Z��m��\�鬋�u�V�a3"�a�� b��T�ԾtBI�!����f�CU���d2&]G��P�1$6�LQ�ANQsG2�FpB�K�x_���De'����&M҆��BP)� �[\�Ɗ=A�ǽ)��P�S.��Z|� ����+�����vH�W�O����:�U^�u�ލ�6pr�Q����0��,dZ�FK��,��So]�l~6�.�[�(�T)(��L���lbqp&�%�M�l�9�g,�' Cw�L�v<�����N����|�]�#Py����'x|~$��b�cHL/Ƥm"��(��CB��ĴIث��4�ᖴR���Jd鿜�) H�=����@q�2v�DK�ȶk�X��V
m� ����!��������O�raѨ-������e5FX{�l��ꟙa���J�!$Z�Y�m�f��C������6N�"P8��3�+Amg���Yi��얇֐�6��7�Bϡ��g;���^�i稀$��M�jP�v�|��
`�5\��� ^c�6m�x��?�d�^���jb�����,��hQZ��s_R�!���3h�PfeC!��O7��T���ѶyuM���;�\�~��Tyzxbϲh�:�aF�&p��a��\=^�	�n`�6L�O�H�W*S��lRl#:t�%�0�9 #�І�n9�˱�J�������@��'�uT�R�FE�z ��"$����뚜�C0��Q��h�0�l�J�oȥ����h(���R����0��j��3�q�Y��4x��P㜶dFԐϤ=��|��rR��l3�O��!��hDd��-U�N�C�;�E$WO��,�>?1�l1깔�_G�&��]�hg����Z C�ɚ@�X��+�F�O8�a��o�n�9+�3�ohb,����E��J5B���y6�w%A;a,���bb6�<�I�K4�)�1��vc�Wۦ�4��9�{bN�|��L ��k	x��b��.�d[���^�0iP�*K�EIpV�v 16��K.�h����9�@����5~OF���%��E#�I3���߆��(��x�O���9' 1���]PP�"�4��0�#�U��:����+e/�m�l���!�T��~W�`�����ӽ;خd �ői�%��T�рy+P���f���{�椵�b���R�j�T�	�B����P���n�0��68��<m���w���J���0̪dgu#�V�^�q�������N��{�1���Eb�_PqH�����d$�@I�/�� ��|2x�\
W�F�I>a�C��03����N�������Р�Ӷ�YR��� q�O[L��3�;:�7��"��7�ݑ(�11iH��"��K�p��-(
#�LbSl#�R� �!�&0![.�u9�Bv�1B5H+���`�!� �����>�)c�r�%Ȑ49 �:&��B`�:r���u�?I��x$=Z��0伪퐬:cH�8M�|�8��ͪ�jHߖ�b�j2X`cZ�Ŷ�3���2����ۇJ��h��נp͂�cP�����xƠ��n�6pr�������CQ<CX+N�Ĉ�X��>�,��z҇Jb�4����,�|0R���%l��>,�&�d �<F_�=C�9o�#-�@r����hf���/�O�GXf�t�O��*�f��,sb8,��b�@��TH;x>�����,��H�rTi7��&����%+���S%Z�S��69Z�B-8ww�)9%G*�U�4�2*���_Ʊ>ͥ�_�����0�YO���V��KC[U8�B+s�ǲ�� �H��7m#ڨҷ��FѰ��H˄�LZiZ��<6�v��iV�3H�-���(�n�(mP�޶w�6prô��e^�q� |B "'��FXm� YFa��E�C�`FH3'�@��Ŀ��yRC0ș�C�Weӫ,����DtL!�����T�¬=�a
���!T��k�Wm��S9�Q���m�ی��bkw��,�[Fo�yv	v��-o���\�[1��nIC���x��T&:F1d��-v��nM���6����ϭ������t0�����Czk�[v�ր:u���cC*w@8�����X-V�]�M|�,�������Ϭ�t�ԖM��T����Jadk+�(��=C`'v�hk8������n��$?�/,y �h ��̎�]������X�p�;P�r{cG���yӋc���}��������#ȶ{Ε����^=m��z�p�6�Ľ���y��X6�x뱷v��	'�:�ry�;Oack�A[/�:c&-�Lp��G�P-����~[��R�zW���4 �� %]�>�<- Z�Ҋi�$��xg
5���z,X-̶N?����kfT��-��$[��<җG
��_��Z���q<���O�?˶�h1�q�Hr-�����h|��U����KsΛ�Y��5��zu� �.K^�����;< d��Z?[o��i��0�m��n�6p�wB�𴤨s�Ҫ���J�-i�Z��/n��t�aV��ϼp��6�F��M�DﲗN���y���Z���=a�2.��܆m��zڙ'�zi�;�M�fB�0Tm���2/�hm�<�@�p��ɚ��<��B�Y,�� `�7�zz}r	�����H�X�d�;�u�e��l�M����LK�!�X�ӶΞW[['�L�.^�YO6���ɍS��ꙩ8�$%�~��%��I��B��b�A1�V/-OʼT�N�	@:f��ލ��'�5����)I�|�,ޖW� ֖��\_p�"��I��r���v�$T?/�i�x�ך�z H����G{�2��G=&�c�ň{c��� ����oߞP $���>�«y��!���s�#;n-��	-���׫����]����z|_����6h'7L�����Jcr_MxY�.Q���W�#��,i��%)�+GN�</V�*�1�Ku��J�Ȱ���qҒ�V-�d����O��;�{&��.�6�T���:-� re>_lזS����~�O��8i`0�G�5m-�0�68L��0 EkQ��8Ψ�kJa}-�W_$< ^49�����\�֥w�Η�KۓV5s��+$�-�8%L]w$�����X_I�:���^}{ j�����0���+N�śŊZұ�ِ��if�V���ޱcKV�$ּ���fY�a���Ӣ,1�p�<Vm�=<<�z>��p1���≢���H6�<y� �h�Ke����+��?����Gu� ���� ��l=�؞�g�]4�@�� 8�ى�i�I[`��k��!iM�:�HGX�w��?�M�V����@��y��C�y[9Zx�w�h���N!�-�봇�'m����韢�֌����H�p��ت��DR󀍍�1?�n+Y���s�w�P�]~�c���\�A�9��
�ҡ�aۍi[Lr��-�ւ���mcG���<����P3��\�/��=��_�`��9?����L�.��zc����p4�֮ڵ6G򗾫����c��t�N�$F�C�v����zjmZ�۪N�|V;�Y	'�9�Y�l�-a�{�.�NO+�O9���������㻱ux����5�F�O8����X"���y�8I·�&� �o��@�sO���_�QUқ��N����I�T֊�p�&��j�A��:�|��ܶ�5��[�-�,�Y�)�m�ZcRN����T���޸Ҁ�Ǡ~D�`�-��_o7��U�U|�L�U���3Q�F����P<I���k���U��ɵm>�^z�v��]�r����
D�>:�V���Rr��]�m��i=a׶F'=I�2%��{�2�>yoK� ė����ڲZ�^ա�4@kk��
N����u�:Z	�[�u�=�b��w��z�d%c����N#����<{$��6���ڵ�Me�x��̾~���~{�f�o;��J}턍���m�ysP4S��-����Fx�u1��s��D�ue��n�6pr��/��/8���
ó�	D�6l�f1��FT�g-�~�c����-�-�����{�_R�L�֞�ާ�h����>hy�/=k��Z�ڋӪSk�x^�������;��x�D���>P�������H�����{m(w<]�':�K�4X��6�ޚa��Ҿ��8F���6����Nn�����y�qHw�򀂧��$����e =	\�A3+������[�z`�&����}v�4�D��N2�i0@��
�Ufy�bp-�W�.k�֧<��Zk`��)���B�����+���Z�����e��!��:O����>���!Ϡ~�j�@7��Ĕ���y�V�K��De� �l|��\�;���M�WZ%_�I��y��}�Nn��Δ���.z���k�!zRc+M�>�~�Y̪�	HxwpH����g^H+&[��7�;���E�k'i)�.�w�ŌZLV��o����n��Ʈ�M&���r���>�{�%>��j�R���M�6��i?_r��5��NV{Ҋ��gHh��x�O+�VݿH�w<-Ho,x�{B��v�lw��m���)��f-�z뻝���?{^G�����=�1c��'�<�gV���s���$5�{���@l06���3Em�֞�a�~m�^��� O��u[X���utYe� ٓ4�3������ǡ�̰4[yy��+OOk���v-�ZTfI�� TP'ʬd���l���md��%�b�֦����>���%�������:�q�G���:�@8�q��i{�07�y�F��x��^�Z��%&d��e���s�yC�*�M�Ev+!��.�8J��.�Hs�#X����B�g��/r|-�Z�X��ƴ�^�����6_��cm�0�}����6_�4�o��A���4ze��̷���!��Њ��l�R.{�w�잱�7�,p�e�ei@;><P��V�Z�1�5����N��0%_�@�f�\���I@z�Y��['�PN�C��;�(V���k�����WV�ND�1$Gpu޹��4;iˁ�I0`�u�$ڲ���eM=`����)���$}����ÂJ=nl_�qժ�5�@��t�{g���;��`�qk[�_�W�@�'�<����ݮ�-�o��h�ŞG{r���|��A�Z�@?�~���s	���=!C�/=��vI���^�}����:�@8�q��.��k ��/ӕ3�&@���-��)1��b����f�^�� �k��4M�.v�,�3�+z��B�u n�Q��LG�/�� !n,�.�$��^�GJC��▾�әPC��A��3���u�XI'}�l̑]�c8v��k��Z@@?C��äC��m5H�.�6�ӧ�ܥ�k#}���(�4�R)��[����q��r�Y͇����j�>9���L�bz�� ���@Gn�P���=��~Ü��K�>̥Xci[�2�=* /;?<��H��������Z�ig��wZ@ŧ:r�:CKe$�3נE�#e�6�y� E� ='%-q�oj�dNKk�M�P5~�����ף���HRO�5#'M���@a�{R���$�ՊX��&O���j�������g,k���B\i0�Ʊ>Q���7YY�C(���>ِ3���qBb襜=��nG�\V�P��zL�R�ԗͭ�&V�֌L�Y�/�T��<-o�9�S��y�w\?�DAP(v!�����[�M��F�)��0	�����@K�������48o�K�d]�'�tU��|����[�Z �
-�>��/cx�O�m��iYO���~�H�T�F2��֑���<k{��6�|�f+-�I���\�dX�����Ŏ�����=�����6Ҋ)f�;(
I �����V�G��mO������2+�C���q��^�	�����>~7��e��W����-X��^_K�s�o�m���XWy��) �u��8.;��r��W�0���������,���.�����A)�znt���['��1���~>؅>Ml'�MͰjc���I�=`���-��X˘,��$y��^�-��!�N�#�MP����z��է�ak��rl^�~�M�=��)vM�4l�-��7��~�J7��i�u�L��N�p��<�8��m�4���:2v��:��Q��li"t�q}8%��m`A�ݾ��ڶD�9;>[s׎]���5p֑��H�m��H$�2Q�M�PT��V"%�H6=��П6OJ���s���9��Ԧ����@j
���-�b��yje���=eq��l��jO��v���,s)���V�.g�,���j�%��YǷ���:L��Z��J�:�%��W�
�b��/Ш�\?}�k�"�/-s��ԝ1T��P�{�B¶.i�1`��ӭ�
8�uK���F�G8�q
c��1���G<+)����v��Љ�#�0���i�a�~�i٥�Te�*k��U�~:2���X�gi�)W�%w���I����\=@(���\��
grN�����f>%?/�K�@Ҹ�z`Mk,<���]2��C%Ş�!KG@ǌ���Hk\�h�z��
 ]���]������$�[c��6o��mÞ��� �h���n��;���6�0��N֋��'!��y���.ʭ��S��cǗ�S�Ϊt=f��l�0��6�y��R��,|��h�Ȣ*��"TN⴦��{]�R'����x	���H�"I �TaͰlL�7���u:2~t������OO�.�C��k���K�!]�s��p���5���r�p�۴ЭFHo��0�Ě�V���N�t\�ׯ�>H�V�j��'������==�"�������8�aNbsa�R��p���Ҿ���OO#i�l|[N�0��x#i	�O^�œ�n�v���Ŕ�ɛB����Ĉ4d��1�!�W~���Dݖ�J~��(���c��!�����extZ�l��_���=����~k1>g'���l�bX�����y�m� �U���1T��#5��7�,s���ڛ�5��@�|�1k�Վ-�i��<�g��i�T)�R��_6tr���;#-	ۉ��J(�,��.35�y��9� �0vk1$$mà�D>�Bk�Ӏ�2ЪnZ���\|��yH�4�,�"���O쐇���-�����v���^v��G�-��V�in��ԌS�,��X9��7��<Bu�;�#��ES�Cut^��DkU-==�ܪ]�5L��R��v�Ć�]��ZsQ�_e(��H�Ej�Io��Pl<��ڽ�����븭�O�C>紃�ok��vi'7N#��Y���n��$$$��vЋ���o��޳֋�u��O x�gzA�o��[/�����u��iq��AJ��Q4<<<��|J�a�e��E���	'G=)1Wv��N����k�xk�OjhfQT�<C��̕��n�ϦU�k��>EQ��rs��R�ʑd��ʱזv�~K>XO�?5j���.�q�m�bW$�R��c��S�����a�pf�ĴzS�1�e���ã����S-�~Q4��cC ��p��S���z�����p����"o�� �rJ��L�9�ˀq7��@8�m�$7F�� �Nz\5�ϋY(aZ��d5y���'��$@O�ҋ�,���ś�-��FK R73��y.kZ�e=��]r�5�?�A��:B�����y�&Ү<ӟ)�깧R���ѓb�Ln]����e�c`^ �wמ�k;W<�&<A��^\+ �P]��˾�3Z�a����D�ׯ�l�x�ϼv��Z;/��Dkk��=]�O^�^�ot{���[�r����<��m)�BW0L�\�5al�ނ�JI�ȶ�M4��Hk#Z�fF�Beۦ,��V��ů�nh)/ �y7���o�.����BY�垔I��z{�Ӕ����k�.�<	[�%�[PkǑf�6�8V�1��p�2�p+����>9�3}c�ƀZ�j ;�īW+��c/L~��y����{@�k;/!�S��j�L�lt󴁓;�������/��]���.�6}��5���񀋼ӌ�jMl����E��+wɔ<s]E�P��缥1��P0�6��R~�>#o1D����n=��i30�,����oICk4�ek���G+,�Y��Ά��q��c�t]��8�!@���e��-�Ćp��[�����X��ʟ=	��׸����e�� X��?��osM+a����T	`�vu�6pr�䖹����aߒ��3�X������.R�[/NL��$�,�i3�u�\��'N����<�lQ8�D_K�u��U����W=&i�g�S�Ml�<�ڼt�{����EuXi�٫��m4��[���Z��඙�X��nI�6V����'�$}�1u��cm||������m��P��e��Y{��s��J���K�KZs��}�Nn��x!Lf~�� ��u:-�o���K�[N���b.��Kߋk����TЅ�1Kr�X;���[��䈭�f�=*q7�%탧I��ö�  �I�]�1�f�L>C�i*l���o+��u�����뭸�'Z��c�� �g�봴��${<�W_	/iٱ��*�+^:(m���k�'r2ț�����i'�M�:��D$��⯧���^��[͆��6$mO�i�e �IS� ����r����Q�K#�2�����)n�'��=�!G"S�\�U��>������ϟ���{��ǔ{��'�{�<j�YO�o�i�O;��z<�ǹ֖@)��ú)m]v�ux.t�^��:�44���@\�شJ��Z��=���Î&@m�n�7�[���jM������q����?Cޢ�-��)��ӟ���B�'���kjkQ+@)�t�����\b����9҉�M��Ü�)����4���S�E�hU-A_[Z�=l}���p)����i�#��h�����b��ӂ�VZ)�*�l��xf
y����H'p�	��1kLli= ��oA\�����)����Gk^�2��+��a�X�Zm����Nn������HI�d|7$)H�[c�k��(��0�K�'�y�ު.j��ʫ��qt�t��7^�������O<6�����`?��*��f�W��^��k����8m����+A�Ћ�*]~�a�^��on�:��.���)��u@:�<������蠂ܕvC�[�P���"��K����\�ݘ����8�9}�UΪ�CvQ�9	��vK`F њ�����~����OQ���dS%m=�\(���B=T'�r�����/���:�8=a6���ɝP��qqM��y�i=���Cr�+���Ug{��C��^(�ٕА�_+�Y�}����0x���%_�[�}Pp��Đ�<��d$m�j'��:H�9N���~(��u��S�y��fLs>M��l%o�T[�S�X�\nm Y�#�r�B���*W��� �Y�o�����q8-}W������&E:�@
sj(��j{'�W`t���}�B6�������\m۹'~x�?<��K'mę ��Ҧx8W�Yi7d;&{S���7�tٵ�q��*--����h'�NI�QKۖɟu¦���4$:N�,r^x�^����ŷ%�k���W�m��(��]5-b��n���Gȋ8׵v�e�LthkBl�Z����L$�9��ζ� �_, ���8� ��j�qᑧI����u��fL� �hs��E�j���&@�kb+RҶ�b�h0��%�;Ï���O�I<�.�Y�������#H�_�}$ߎ��Q���tk��:&\_��/�C�^���� m�����8-ƼL��"��IoA�%�`<W�	h)Nǵa[yz����r�f�)�ω��U2_`1��;�t���AW��\�C[e-���'�5CV;���~g�׆�n�{�n�{���ٓtm�5Cl�O��1����(q��c��v���<vV�@�4O���Dt�|W�;��N���r倞w�[����o�)y! ���jPWo�ȕ�~���N���w݇Z�)�Z㡷��ѽ�N�XI�R�<����^�[QȪu=F#�����,��<=�4,-�ӽ�%-v�3/�quJ�%c���D��ޖ8'���ø�n�4;��@�M���߄[����I-gY:?�͖ٖ۞~�������Km`�>���u�1����l|����S�]����j1巾�����ޑ0r�׎Oy&`I�e�{�h+=����H��H�D�'wO8�;"�<F�i[�4��N��Ȓ������f=�7���K FH;��9}�����9EJi�8y���#�>�
@��f�1V��� =)��Я�W�����c�l�- �`I���=+u���J��v�����Z�V�X��![��U��42v4�u�3�U �o����"�����Co��x�p`�J�O�&�{Z��=�oڶ�}(�G�l�m��E8�q
a��
��M��5��1F*t��
k>O�ӿ/�ͦqI;�ctv��~�����(c����<�0���б����)�	��� �Lt��$M���/�{�`�[�p-���<�����c/ϖf���i�o7
HS�qV2~�mU��SCT{�"����6M�[-��Z{��w_�'��v�sۛ�V#�*+��[cޒwgҺ����m���iT{�5���$�㴞!y�,��R�6�2�T��P3N�V��
�[|�"n�E}��L��)�/]��I��؞����K��� Q�B�x��}w)��D���JǶ�u:6_;Ze�a��)����򧜢���<`�6��[Q��9�(��&��=��mN4H�'�lz6Oכ�|��mӿ��>�:�� ��9��s/���[��^\���ZB�0����c2������M�u�W��٬踲5�ݣbӽD^��+��*^2ԋ�t麟/����1O��� ;D���2��
��l]���5m���_jo;Nl<O*o��˥zxLN�Gƚ���s��Gx����@o���
�
�0�o,s�v�g��j��k�
��D?���|�sW��	�VkCg�'0x�3�Bh���m���)��h%�ؖD+ԓ,[�[�_/t-&�I�=I�y�c�v)/vkvbW-����I^y���6��N;�\`��e��x�	���� ���[R�6���e��R���� b'I]8�J�Aw5B�R�3��<ɟJf���_t�9�0���Wn�dc��y�D-K�u�L��u= pͼ��/��Ec��- Y���YoK���:�צ����y�.�`����8���Qo-쭲��h�d%0/�}�:�b��J#a/�}�ۺ��<�@���$=9��F�W��!f��"�J�d�G���mS��1u���\��S�c��cm���s�V���5$�">0a��g�b�@�	rX�J� ��T�A�Q�IV�l�pc�)��؛A��p��>��UT�3�� `�@u^�FH�!az��=��k��8zLۓ;�?��&��V�޲����J�JѺ��N��^i:4��H3��4Ԣ^��YO����Rk���q���l=���p�	�ve����/�yز{[�=�I�*��BuBƦa��eF�~��K����^�B�i\�9��O�$4����QM����@��3�ðj_��#�ۦ�.��l�YA�7�z[kz����;��%thj��:��Z9�J��n�6pr/�&�l3x�M���D{	�x��sI�����[����j���̂?���a��;�L]O:MoV��R�g��d��Ե�|����3��& k���s�Q��+K��2��vG`}�\��w([�m8Ծ��o����᭍Ks��$y��ݖxL���4�۝�ҾX;1���dX����m=�߭�/��6��}�N���s�.��x���Xz�/ZZ��$n�i1"���|�{�����������[ߵ'�F}<pL�2��-��QZ�WL�N�g� �V��hqt=�6�M�TO�{�Y�Iܽ�~*��~���SƸ>J���چ[U<�-�f��R%�[�}V �cL��ZK�h���k��ߧ���F7N8�yJ{Π����.vz��fQ�䩚��B-�]���E���N�e��Z��2m֜�4����AɛmT����[�*��l���<׋���u}��w	�H֑^�Ay��b�td�4�t����x�є�������,��D�f�IB壤.�����o��씿{
,km�|��m=t}5�j9-�^�Y�cmPG6�s��ђ��<�U�=�d�uJ`����8�]��җ��sLgѲ��TX�h��2��{�k#@�4%�]��k%��L!١�a�>9�D��^p� �n�w�>��|�xql�h����@��S�\(^[ۭ�`{���0���V����B9�S�O���Ig'���V�9��ߥ:X��5�ǳ���������*�6\�A�y�2@�Af�1�e� ���=�N�0d y���|�E���y��/�ݓ�-y��R���{��fE�6e���:#Ћ���=E����W��Li;h�7�����'�2^:�������w{.R˕�����i:��+�J[p�t�W�^�ʏ�d?������i{m*�j��V�6�@ݻBBߛ㵯'�������X_3�:r9�gB��[C6�}��ɍS�Cs��%qk-��Ԯ����]�'	����A���j%Ȗ��ӮO�2�������6��^�x[d�u:��皅ٶ�gO����5�i�t~���k��� e�졾R �{,�1����
� �	���x��p���4p;�찯j��t31��`ǁw1��.Y����;��m ۦ�(�=9e�R�+e�p��K��}_~��v]ڀ���Nn���J�5�@5ive�����+�Z��Y�c�����2P�ᵞ{���4Mh�XC��I�D{�#8��~BF(�����.E��7����w�@qG�q�$uɲ����D���k����\�Kl�I?��KN�r�H�0�;l񙘷���R�e���Q��Q��/(f
\D壆�^�K��=Dx-� ���4Ւ�.�"Wk�r�t����
/u�K�R\a�qJ��%m�\���ҾbS]Ҡ��B�O����z�_k���4O�x-m��^��Z��qC���A�fsr���;"4xL�6~��xi�$h�� xҕ��d�ӱi˧gз����PTƢe��X�gP�o���uJ�lI:s,ࡄ�5��>Ea���ו"c�·�`΋����$�V��"��Μo~����X�hF)8�S��K�Pkn��)�9�����7DҎ�c�!��q��PD����4�!׌�oS�g��8f{��+�J�h=7���ǔ7~�q���o�m��V�z�� �D��k���߱�M�N�z�B/�����]s����4 �pZ���cӴ��׷'5wbzє�f�e���o�-�����ߵ�Z��s��|���/JNy�f`�.U ɕ��5���k�]k� Ä�˒�h%$�X���4�*�H;De�qbJ~�R�!L�5*�ڪ�����,��i��H�x1Gf�rm/m�͑��e,��Zaz�z����l\���z\S��nt�������bS/̨�����]��a����]�et)�~gc�̣��K]��V�Je��纠͉��;[�/t���k�[�����:,33N#��t�f�MD����R��_�����wV3U�����&@!���ο+�b�b2��R.��v%UC=��~!���1��D�f�t"�JJ�hR�����e,Tڏ�'!���m�줭6��c�h,�v%��H�a�ω7_�y��l��t���ڰ-д�����8-4����ia�ki�ǔ~d��Ŭ���K�sW�ŵe��d/�:���v�_�n��3ߧBL�7J��X ��O�R^U���K���TW�q�V�R/O��{v�zyj�����U���u�G�@<��o����C� I��[
XH��&�9�5)#7>� �gU̅d�5u�pEm�q!��2v����{m�jۿ>�v�/l|o\]���X7���^:�uE�+�6�;���u&�,(�i����.��òһ}��`�4+��=�I��iZ[�*���{�$ �.9��=Ǽ���V6'-��'��l����*\ױ���Jן��[��x������$NY��%�e�����e[�B��Pk���A�����)�jM�؝@̉�~���1�q e��])��,u�M���۴^�-���p�_4�ռ�
�r�4�s_�����>h'wFy�Ldխc��'M��vQ���n����Ꙟ[`cU�<M�!owa�M�}إ�8m���4B:te;��I�l=͍�뫤�V;��v�Ӆ�< �fخ�Z�O�c�c4��:��_$�K�*���nb.u��U�Y]N/�<��6-��VF��� T}_���kFC��]�������P�BJ��v�W�WEhbo�k �y��iB�d�m���iJJ�����`�3�x�^PZNͼ��R��f�6��ۻA,�i��,�m"!1��= R;~����4��x��<�xؑ�$A��K������*?4�+@�nh�-m�_ޭ�Br<����z�&&�x�[��'T����q�\H�f:�I��'��:�����Y��&��" =�Tz �M1��P�� m��@1ֆ̭z��4����x��5�l����?V�l�mU�9;���i�e����Nn��q�!�;�׌<V���)� �&O�n1Roa��p�-^��Y�����~�JC����#�C�ř���(*�9j)s� ��z�{V��mu��Y�%,�h�'�����U�Y��ҼT�Ro�5C�i�1���k�Z���gD֎�<��+��[�]v�v-�B�|�uu�,��3���'-�ꥡ��]�B��������mt�UBۭ��A8�q�i1M��L�m�G,��7Z��5Zix��]��iY{V�hO��˂(�J��O
��{v,#��[^�k� ��-a��v�}8�N[0������;�P_~f.T߇��S�J�M�G ��,��F�d�@��T������@/cfLF���X�!���"ȡX�#�C�f _���N����Xu&�cʟf9O��ti�>l�\Fu�C}�\��H��u	��%(̎���k��g˨������Dy�����h���t��)��։��</U���C���
]$�f�!dڼ�ܓ��/�J��^�g�^KN��j�ZL-�6?'wB8�*J����M�t�I�6��)�R�Vb�R�.���<�
O·�M��ՠ�*G�^@,鈖%$C�0(o�鏵+�v�+���c�=�8���r�9V�7�A����9��g��k�z��U[:���)�^Q�A��xUmbڎ�[Aj�$�ߦ�uE<��́�����A�䜁W͹i�����7:�[&��z��WO	�����f�R���P%��6�����	]3g�-@���ق��hl����݂�㵤[[>/?[�P����5HaSC�CPL�k-�h]V-ͫ�ҳ�W�F�ˋ#��C����[�κ�붓���z�͖�Y�%ۙpۄ��M�8&��Kj[���� qT�I���/:ͼC�gz�]S��o(���~E�̩x2F�pT�Ҷ�04��a��b�`���̻"bP"����V��+J3��ҧP�k��ɍ�0$qL�iS{__&���C��ȓ�tz6�'�t)�Zǚ��C~�$K-��2y̳\XVSH����>O�l�r^����4�h��D)L�H�u]| P�S^�)�p���m(Ͻ���8�����<���1�[{�p��i���~bn@aa��5:E��ʼ�:�^lAif� ؒT)Ę������պ_=@(at�4����{
\�� �6L����3�o�9�<m0�<��mt#���[�����v������8Si��[��u�^z��+�W���jqVy���za7��t>�~�'�5CaxF�b�c�"�̚��J���~���������v댅�#�Q��YDٞ%��b1�?ŊE@N�H���8_]n��Ӛ���#�C�W�͸z_ R�e���N���W��Y�~��AO�饇�1o����΃�tJ��鍡u���W�f=nt���[�1Ѽ"hK�{	lHx�Z���6���{��rp��4��R�W~4�ړ6ƴ�P���nO�
����F��6^����-�0ډ�5�B��v�����NCk��wK��k���bm 9TҰR�n%ߡ�r躖�ز�����y�ZD�%�1����sۊ�hu��5����w��M������3N�q� ��빥�R�S.s=F�`��j-0�$��B�y;�s���; ��,��˚
� '=&��8=F�%��V�b�-�^�3�Bf@:,K�S�RR��\��Qg RJ���aT�7]�� �^��cjm�Y�8��2���IMP��4t]3�56�YC Hƿ11~Vr(�Xo�ym�1�k���X���ΠR�+�R71��6�2l�y���ӆ����NC�ڪ��7�{�����_��-���gvotߴ��;��2y�I���:��m���6�,Tr�FےX��.���.�ZBV�ʣ�nJX-�Q�K�oJ�:��%��T�S��'3�
H��q�,�����_�BZ�k�4k�d�B�(B�Y�Řm;���%�I�M^E9����·� �-���`�u�B|x �k�U�y�f�IG�i{D��Pk�j��Xpo��)�d��=��?��րY��'|ڂ�u�����m���)���u���	���,��-�sl-f^Y��A��*�m���u=�օ�i�UZ��,���W&�� ,Cqd�Z���wv�vZB>�!��J��)�ϴ�

?^D;�����#��%h��M7sE\e�nE��h3J'��҈t������� �ua�W�>#����6!c.&�k\B��0M���I9Y�z�!�P1���	��u_�1�O�������V�H�V[)�I���VnNF��Y�R��v�=#b}�(�"�����)\��m� �S߇�-��X�/�X��=XB�ʁ*ɪ~u�u8\7��=�Nn���x�l�������	�c�?a���K�Z"�t�A�}.��K�i���4�[~�.����rb�i*Κ�.2��Y�%"�-��$}5d?�G 'Y�b.��N�('rȶ��v�O�,i�dP˰�d�X��R�R6Ța�$����~,<.�v�!��@�MsesCb:��1ݥT�Li�K��Y�~���
�F��,:(Fɫj��K3��0�� �?/!Ό����<���0���+�eÊ���)���g���'䊎Ԉ�����Ҹ�Ӎ�S���z=	�tF���Dn�)��̜x��������w�`�oi*�����p�dp\=��i9y���Ԯ��;����8��᜘7Ҭ�l#�<�Sc�3�ۍkf.�<
�n.��(S�X�:�b�停�U@[)��!9���qf���40�7,��|���s�u�4�u:�ѝ�Nn�"�v��3q-i��U?��K�B��8����d/o�޲�U�Zb�K��K[Dw�$C�/�*Rӟi�$�0<ųv�3���6)p#�.�9��:'�	� sBf��,���°>�Y��������&�����8f�7�U�����&kx 1'ڽ
&0Cfaf�O`f&�-� `��;ld�9�	Ld����ط�D@��z˃� ��6G�I�Ŏ|�@Ҟ$�^�$�T(�3����8�va\Ӊ=c��Q�����V��K����	@�K��?z����5�sBƲvK���ߊ}��a<�'W�[7<��[�s�uTi�Bmg�����h'7N�<n�߅q��8��GEA!��W�������xR���e��k�I�6��[/¼��Z��!kna~��(�n���ȄN�31+��ւ��S`	��7$��6d�,y�&���V �ML8o)�m��%��/ ɺ�A g�Li�Hڦ4��I��~��`I%ĴK�[@ɈU��YbG��J����SI�"��Hi��e�v!-������Qm`ȅd-&&�W*P�E9%#m�P{�%�P ����4*��|o�h�X�D`zF-
���h���@{ f���ND8�[�v�kf����� �^�kg}B:�K��-��O6,@�au;x|�2�ύ�6pr��{$�$������ѿ�	�ڲ�w�2��1I�:^O[sM�V��Y�,���,~�p��LZ��5�\(��%�@̊�,�N��M��([+r�*�;���0��B�B(Y7𶺔Wl[ԝ6	<@�C'Ů�`Ұ���RTi �'Y�$U?p�X�ꙹ�/a���I��|�X;��z�]d���*sF�~�mR�$������1�]�j%�4� w��0�H��UC	��*�~_Ƹs'�8��O�D�d.�Th�����i$��N��y� �hNd�1��Y��@�WK�Pk Z�ڂon��v�]����/��N{��m�50�t���6�}��ɍSX9�U�VC���z��,��jW<mHI%�z��e�Ro;��z��<�p�:[~��T⢭��ۑ�
]�H�d��Hc��4���y�L��Y���VR�03��r��
G59.#[��,P������e���XS¨)� �+mT#NMW0�DC�u�;'�!��;)����`vb�X
�o���`�x�NI[��a���m'r[���Ę�X	�_,�5CXm�Oq�o�Qs��Cb�I��z뉀���_����?-�_a>Gx؟���m��p8<,�_�\h��v~X�2%��cm(� �%$X����E�y�Җ��)�6���ɛ�ٞ�hM��c�ۥ��:��d�Cꁈ�d���4��v�$QS���nIq-��z������/8{yyY�Ѵ0�wx?���m8��fbYT�=�,�p�g�N�R��0b��H�vNZ�"駲3cJ�̆��K�;=0��ISs��xX�YÂ�6pӖI�.[*��9/Lp�Nf�u���V�*hK���NS�˸��F���<����
jQ�N�7�&4v���>���4�E�����CL 8Q'�T[�����M��� H�i��T�%�rZ��nA��i��Rv(���.��@�߿O���-`�l�P�0��nvǼ��Ksӛ�-&�Rn�"���6�֜��d�{�]Z6�P�6pr�4C5�=��m�X���vA���Z�޶KI��H��5h�Լ?B�F�+�X£����k*�Y|x�D��~�����/�˗oHA����$��VCj�9����I�RQ���'i�ђک0eP�8iJ���Ck2L�m���v
k?�̃g��a��Zf�34�(.d2�M�K��F�[�;�=m}��2,�B�&{'s*w�\��ڒ�˜ۊO�H!#����aCҀЩ�0��(� �Zr��n�r���ݒ������Qd��q��#�(!�=���>|'٧�p����i� pI�)a1�4;�V���d��4����^�������b��x���������]���e�)�4���s�f��m~�3m���$�!���b�j�c���Moo����#-����e���|طH:6<�H�!-慖��O(aC�>ˬ���C�II#�J ��!j;d��D-N}(�PcBCte�X}b ��&�1\��~y��m,�H��9��:o'�	��f`
zΐ�L�\\L����}��~w,�87�H�lϢ�I:�$ ��Ff�Fc�Pf���! �����*w���<*� ��O��y�v>���'�Q�|�A�񤵅�mL��֧tZۧy87�P����[�������@�MG�.�Z��J�J?��m��n��`�&V��m���[�Z[)=j�tm�-�qo[G?o�p�wV����;�$	3}>==�����#)Ga�33K���k*ȸ�0��+�K�!҆1�t7�|�'��!8�,fHL�>�B�4��1m�9u�L������e ��!i'`2�\֐���Rhxd�a*/���͖��sH�c��"T�1=簁��,��HZ�@RS��b{�b +�tY�3��u��>�,�q�d�6I7�Y��!�|���8����X�=ˊ_}<���>�d���v��M���(��<տ�2z���G��u%�>����*@�P����6pr�4���0�V8OX3i=0 ��Dz�y+�x���`M/��soy�o]�.4��9Zz�����v�i����"5��|�������5���R�Aկ�0�sE[�Rb�����:��U�t�V �˞]I���	�~y���Vd�㱬��v���q%�Ac����t���yIw&��霘���1������:YKv$X�=���N"��;��i��'mB9�+�Y�YkN�}\ G�w�d�s���@:'��Q�(N���^�E`�ǉ0ft�&�%c]��y �jK�ة�5��E�gc��K\��i��M߫�lYtX]7Wʁ���P��^<j���:���Nn�a�'f�IK-�E��÷T����{���o[�gW�ձ|Z�p�]K�C�� �9���R2����үx���i�`2mS�k��J�!��X�n���L�QN5��\�'�O*)bҬ,���[Jt�&��U�v��
�-�����#���Ҟ�E/`oG)�	��l9v�@fNɻ(zW�sr�_T��Ϳ����,�4H`��X��=C@6	��4��Yo$��z���i�[//˔�ς����u��~[����a�����Ŕt�\�+V��C��xkj�9���ɍ�n� ��[d���j'DzG���-|��P8�PZ��{f9O+$�~楧�8�x|�C$�r,��Ȝ��-k�͌z�� $-��E@EU/��^�9-�䏚��x"��)�d�����,6��m����m�7mﰚ�B��=�3�4�̠øa��w�����ә6��ݸ�A�&*Δ�~|Z�<�i�t^�.�e$\��X':4���a#�9�^J�3���< Z��Ѱ�ۯ�k�<��ˌr�jn1��?*\i�k��zc�c�ܞ�k�V�V0��hǾ���,�!æ�1�����7����=�
uPz�b��2م���{�x�{�x峋�e�zX/xZ�lտ,��&��C�aꩱ-��防��6��g`�f���C��@Z
�^�.h;��7�Ɓ���	���g�Pp�S8��v�@9-���k�阴��M"��"&���%��L�Wxh�79/`d���>�U3/�a���������������
p����4�-t�	4�q~�1�$~K� [�q�1eF&p��O(F�k#o��~���H�%}�-��1�lYz�Ƿm�KZ����ڑ��֊�K���ތ�ׂ��n�6pr�4�=�ˢ�,�4Y¿B�jI�^���۳XI��+mo���I(��'+F���^�<j�|�e�$I�:�!B�& &gt0�}��>J*װ1h�W�Vm9����m|7�gU��	p8"{V`O������\��`6��g���� ˻i�#^XG6$h�(�	O �w��~" ����Z/ Ǘ%��'��.iO�.e	{>�;�� ���>P9���K��%�+<.@e��} [T����<���x.�o?��̷'J}!�_�V�t+H�����$�ZԨ�J��1|�_�� �G���M2�7���|�����Vze����A�=�Nn�����&vц��JI��PޯA��^���G4�`��idy`g�驤0��S�JB� �|�){Ͳ󏲝C�0�8$|�2X�h�F	�� n��	���Bp�>��:f:��`��N�H-�y�0�|$ ���w�|[����<�z��}^R�Nt�w��	��=���~y���t�a�@���?>��D�3����	ޏ'���ߎx��������~���>/P�q��}� ���������3��� p�M���	�Y���=nKB�n�#Ӄ:�#�HX��д��%9�S��h	��(���6���Ӫ��B��ys4��z�Њm��Nh'�@A��IK1-ú�V��>�Il@(a��e^8� ����s�~��6C��H<OR�����i��QBy�U�CΔ�|u]=�R(�����d?�`?�. �};8,`�m_�� ��6ؙV{\�Ǉ�~�0Ñ.4dM�c�
�����#����F�_�ﾛ�pOpX���ox�f?���Ϗg����i������ڂo����zy��	5�d�0�����v|yy�/񼤷�����=���d{���$���, ھ3�@��U�B��I�6GQ��N
��UZQiM�1_l�����o]������hbZ�G�m��߽�E'�m��z����Io]���i'7Nޔv�d���.��|J�G8�[�k&[KH�*��!��r]Cz/ۋ[�#
�D��֢�,�ZGcf^�]��0�y`�p�)�+�%m�㴲��D��v�|�?���.����0����:N<N�a�<.�d���e	�H�I�%�s�|����W8�Gx�����|z���a����gƸ�����m-��{��q�����㸇��+���߾�A����%�����O{8���|����;���.��#ײ3���09N��CB�6���z˥i;Q��v�zi��V�h��g/���P���r���N��l;��g��mֲ�P\��!�^h'w@<_L����Yg�QH^^��t��x�BrQm�EQ�)�|d�.'d��+8���D�4v���vn���*�z�Z�?�Rk����cHL!���:%g �5*�@�}' y���B�7sf��8�~� ���^ v�p�=�3X� <M�!�7˻a��0M�:��XL0�O���>��m\�||���>����^�1]$;D=���>÷w��y>�3��f��~_ ��y���i��󼼟�'x"`��S�_�����.�l'���T���A>Cig���;3�-�mP�)����M�\�����>@�lR�g��%���LzBBK�鵀^Vot�ޖq+NY+��ܭCsB	R�o��m���i�?��h�/�2�*�f�l(),M|j�?��q�%AxXu�@o��ҡ,N�v�SC�n��EU�hhm�p�
�@Q�i��TuT��q°Z<���
,m%���`���s�p��xHL�*��Њ��hH:<�y�qz���>�_���o���m?�������#�g8�_� �� �	�x����*����T������i����{rY�'��Z?�/���~"p󸀞�t���|���K����R���0-��m���� ��\=�x��vK@�4l�R����X}�����@Dp�2�-�[KIb�J��H�D�Wl�X�>��y��iR�2w��bۦ�U��+����Z�6�T/��i	'�0{5�F�C8�q�t���6�����%LK��e��pA���;�ȶ��Z�0�y��֎�)ϻ-���>Rl���9e�i��j^ؓ�*r]d�1��mO��;�j7��/0�>��]��ׇ�f?���7���|N��$w
�p������-!�U<��JAb��?�0������ �������\����q�3��q��1b�p\ �;�dOG�g���k��6�ϼ~�}��N�S��Z��뿖6D�ho���`P��S6��_Z��jO�X�A�o]\����mt봁��=�ǐ����KI��9a�Ö�ʳKL]�KR\��j�n��{n~������O��� ��n��:Y&'��m���~z2�{y�z� �&������>E^�w���~�!���B)�'T���D�f#ރ�{���ՆH�a7����>�EY���H6'�n�yz���>��ے�	�y��R���|�:F8=~��x��~�(��p�ze���,��b��w��D��[��녹����ͩk�W�<���W>�\SM�mW=���8&ş��itYP��׍n�6prD7�^؊��n����8�zL��J�:�V<Q�Z�-X=vO��Ьf���ގ�.�V�m�K��}��8�0�	������� <-`����� �ఀ�O��}���grw^b�#ڣ��p~���+|8�_�'؅	~�x�O�H.�_Α�hI`���~Z�˷ӟ`<��ܯ�����^fԣ�������ʎ���"������q[�\ϯ�趰��� ��-��#ֳ��}����� J��V���ݏ�}	\Q�k �x�*��Y�xu�6�M���͓���'��:�W�F������v��zV�j4<� ��UM�ɰ�$�+6oF���ҵ��ҳV���꧁o�E�AGj	ņD A;��]�ȟ�}<��m�|{���g8�i��o�3<,o�7����?��9!^F<������o��<¼{&F3�/ ��+�_��w�w����	�Ѵ����wx{x��B�i6ć��0`���ŉ6x�����k�[3}��V���j�qk|���ƥ���1k? ^<�^SC���496|OP��n�[��-�"�SŞ� ��N�(���Z�6�Y���]�ei\��IK�t��$����oO�ԋ�'���#��2������;�oB�i��T�Mzmt��ג�=x����>=_��~7N�9!c�৏�<��/��|���� ��<������#�^����~�������	���i�;�����={�W����~ �S� o�����W���#�?Cس;��<����o7����$������8��O+�v(��x�Z��r)�WN/^�x�B�3]O{O�%����z���7�m�\;�a�{���<�6iN����k�"ԓh��yi��1��4h�̣^��Q���:x�n1��LƗr��^�3���7#�GS҉�#�@�S�ޏ��#��i���7�yw�?��F�|č�����,M�'x]R��ix}�/��v��}:Ӵ�9�8�m�@'��n@����_v���?�/�OpF��K�^�'x�/ �������O�:��ͨ��/˛��Yk��Ö6�C^[�g�);v�E�^�V9����ix�[�����emk����4=)����y�j���G��Uo�9���;�k�LZ�vK���/1@�����E̞D���5�k)G:Z�H_-��j@L>=�fߕ2G��dA�Ǥ~(<N��"��a�Ȩ}ٜ<������o��� ��i"������oР5�A����Dm��!��� ���:×��𾀋��-=�NL��"=O������k�e�ݒ�N�w�ƥl�=]8��_wh���$���`2E�T3jU�W��Ü���n�P�X�ڳ��8��[ZDox�ye�J��`O���A�-wD�0��kaA��>��/E���	^�7�_��ɍ�0�I>ewL�x*��Le�������]D{�]��V'mL(�v������}��+���ƶ���:��Ā �j����D�Ջ��y��G�!�g�W��lvdO��\�������0��˗� ~x����m�_l슶&Ӏ[8��얈����yx��4<�?�8��z���} M��1�04Щ!�ir^✇N^�� ��b(���;=�mx}L\kz���0x�U�պ�[�cY��q>�n��U�7Ͻ|{s�������s�)V��vE�����6�r/���'{zk��"�Y�{�UO������Z;�� �����
X,���Z�p1��6�E�/�fx= �뇺���d����l6���یਜ਼�������@��B>/���0�������0�>.��0���a{�=�	�Ӆ��(��� !.4�H��ж���'8�a��yy���t7�4'�K=P�vt[�q�^�����E���
���M�:mR+\k�zm���?��U@�=�i�,(�my����|���j9Z�5��e�����Cⵧ�A�[�}�h@���6���ɍ�"1E��J��s����OK� B�t3����z��1r{�+��|J޵ A���0=P�������[����O�w���]��#i#^���ny�_�p��x~�a7�޿�q�i�b�u��2��@[/��x���uA��9�N�`�#n� K�LNK�/�%^x�c�<4��&�A��(���
��9�ץ��;�"�VHM��1�u�r=�� ��n�����j�������liR�\�s��۩l��-1/oD�|�.�@���
PU��.�F�G8���/0���5C_
�ԥ�\,M����ڏ~�-�a]�^ZͲ���~��0�5x����˥z�V��ŝ�� �?�g�y&�@�]�у�#|��
���� ��
��m�4?��ߗg�3��3��^�eA
��_��!p���q�;t"9k��>�MK��g��_N�/HhB>Q4��)$wk�a&����s�cؒ'�靨��KT�Ʒ�����֋� ����<�x^=D��i4��_S�V�k��u����߭�í*��=;j�3�ao��i'7N�.b�j���Ҏ7W��%�|�Bi���2���jq,yZ�Ka�̧!�z�YI�./��E�c�l��0��D��xMDW��4M龛_�p<�A8/��?/�`�^ޗ�O� �LOp�F��-e�䢞�r�_��yx��mA�/쀎�f���\~@��{u���xz] ��/@�<p��m
- ��8- h&����3���^�DNx����8���\?��9:�~�Q ��/����S�ؼ�� j.������O�q�yP4>ghn+�����;��O��պ�|�����8�\���B�f�=p�c���^h���I��<q�jB�^dN�&���^xK{�#*䵊r�x��[�+=-�G1��f'v�t�,���1�e���q�}��� ����)��	�����y��Hr'�@^/�QwU��W���fF��)�>��/Iߌbm)͸�h�c�l�Ԏfȹ�>���>^�;�� ��W6��~��@ ��@�/~����x�����j��'@#�_����i�I�I�Y��y�ԟ��D#���@W�H�0%�]�;p2�6�!��Vމ\����2(�up;��D��MW6Bc�prj(���B�6��)��t=�R�S�.u�I�0r�!\}ڋ��o����p�U�� �K_���JN�\p͉��6�Ӏ�FqK�:Nkdhyؔ�h�w������F�<l�xi���T�|)����F���{ɔtl'�O+�����Qg�p}P8��ā�ٍ��>��E2:��U�#x@@��ū�C�O�Q8�&�� �ﺀ�8��tR׺����=4V��H����ˁ�4�C�[�j�g%#X���mqj׶����MR/���%7�Y[
k�{Au-�����ڬ��jC!u��&��&����3�]!6Cn�WC�P:��{��O�v�mӪ�+�qX�m�z�N����E����th����4���L��~�]3�o)Y�8�d�7��p���m�]�[n�杽�y��-�Y�����9�<������b�_}$E�3_z�t��ʯ�@�����Ұ���(����r�ٞ��<��GVX,x�睑��=c�_��3@����:����)�)@.������Y۸�,�,O�bY�^5���m�+1�D��|w���=ͱ���qf��Q��B��eDeL�H ş���س%_��ɮH�ut����#&.m�]P��)\ޡj@��~�[7�&��\P�?���ƀ�̿�,�IR�Z<�}��&�R�z�^�C���Ӝv�|H���7��2�AR��R�+N�xf�X[�Z��!{2B�jh��AA�ï	ι�>NϤ�Ap�Z������%�e�#l
E�.%�rm*D7~_+;>r���D���3֦�@f�K��sZ\1����xĜ�x�~��g7��'�
��dN�q��oN�q ������d�%MǮ/OKb$�Eu`R7~�y�7H�����s�Y�(�&r4�ia�'tj��a{p�򺞾���lIҔv�~T���P9�?`:I�= ��	28���xلbO����0�aɩ��sE�Q�c�Q�b����S�曤���%a�"�/���Evޔe�����|��p��`�wR��^�i��O��ű
YV蒆2
T���{~0�m}� XA�O��M��I|��|{�*IsGI�iY�K*.�G�������lhIVD�R϶�%hSi�I9l��g�w^�����d���������\�~��{>��h���s����/�K������߆;w�{�R/��<4�Z�a�@���e[� �^vGzp�咦ip�	�3�V�ׯW��I��k�j���'I*ﲛ�4���3�M����z�$�K��S p�UR�n���h@���'5#R������3Ww8P�.޽�N
��
��	�0� v@d@E�~��.��N�w�|�~��K־n�ʗ,�[��h���oSa�a�ʥ�A��u�������^b,�kݗm&ֆ$Ƨ�d���,#Mp�OgV���]�uS����`���tϞ?���7p�����|�'{�=������C������w�����s��%��ӛ��47��!i�Rx?�����z����4(nv]��}��=��e�r�ʙk�z�_N��2�Y�����i�^Lgi�by����L�����9�̋�aڦ�ӯ#��7���I�M��SD�8?�ۍ�ȁ�zR��2�� ����,�+-OQ�y-O8���nlH����"�ῥ�R�-�
d��崌&l�O�}�uU�Yq�p��_�����dܾ}�˥oC�����v���+�����ǃ�����oԣZ�Z偯I	�u�����^vCzp��l|�{��K�u�t���&���bQhj�K>L�r�%��3V8>bm�O�-�|�w�B;HZ�(g��'��u��srW�;nVĞ��?x�da�eX�1�����╜�˷��Ԉ�I3�t]��h C>� �:��m������~��)~�bU��4��u>�����6���=�����r�r�f���w����`2���ׯ�O>�����0�Nk�b�d9�K�Xߐey{��˟���d�%O�ݨ���w~M2_%sҘ�0��;�nL�
��rh�`�	c��c��i4b�!��-���5#:սb�)	S0H��C;�X.`~>/F�s� ��@�<{�'>^ ��&tp/������U�R��Kd�ZM������m,~�b��5_�l��6��a<�|���������,���u��� ����s �.�|���o�=z/^�a��$i�,��z��#�r�������l��yX��10�Z�dU���H�ts�H�X�nS�����j�l�
i�IuO�� ��utd4���bEܛ�ג�K����������K��g����ү���c��;pFk
��#�݈�����,~�t��`�M,#n�ZqP�ځ�PX�X�Z�ʔXiR���vх�i2��;�ul ƌ��O*��z4�k�����������ٓ������ ���:���~�z����N�>�Q��Π� ��d�4������S�W�0gu(�u�Y�4	���l"�H��ms��\ �q�A�[�y����p����p|���gpz|
���{y��أ��Q�Q�Z����x���gL��8����W���w�·O�p����B���îu��hXqZ�����N�rV��u�n�%ˠ1kVYHF��3��,4ꈀ�"�b1���h�6Y����c@�I�|�w?`�u%e������l�>?U*Gly��>N�v�ꐿe�ؕhM/$�j|bF���b����:�+��u��۰Ґ�X�ܦ�B��hY+�{���<�=}��i	�.�;�W/]�;o`��U�^a�J6��<�g/�Ãǟ���?�'O^����<���O�qC�%ۥ<lc�J�Me%�h$ ���Q��E�����a	��z���c����:������9��'�\�= �w��������y� NOO˶vvv�ϒwغ������Mr!w/�'=8�!ig�.�����5���\��#;U>�C=����O�bL��H���L`i�"����� �� ��צ���{R��ʉ�g7�~p7��Ǐ�����\�r�{�>\�|��\g��A+�������do��܆[��E�m��_�>��#x�����í[�<@!�5񲬶���, ���%K�}^F��A��k#��Hݚ�����^�L���u���,����t��p����Ͻ��k���Me�S:�Gʤ,�e��]�vK���^�[zp��2�*��l�{ <Y�m}(|D-;TN����� e||�%��<u�ޡ�l�n.��:�ܻ]'p��myծi�Mx�M��������x%-/A/_?z�
� `�!4�T�|Z@�ǯ	�� �~����?��?���1|�߃�ל"��>x�����������x��eG��g ������;o�?���෿���Ձ�*q2\�@g��w�^(���a�5�E��$�����4�Q�qq�g�hm��nMWK��Զ.k M�X+ˁO���V^�G��7IK˼�������G�p��W�{>��x
ׯ]����CF�t�@G���y�U�����~c�l���d�e��gJdt%��E�࿍�A�#ɈXm�4e�����4�6�/כ~s}-``�ʤ�]�Z����g$ �n�O\���А~G����3x��1ܸq���O [����y;����|	����{�~/����
A
��z���x��}��������}��%���w�c.C�b�O��J��@if9K@[������R~�h��x�buj�#ӳ��#۱�F�XM��x$���s4���`�xϯ4�s��x�w};°4���x���j-X�ɋ���邺��d��=҃�]�$��[�c/�5r��^=��mMOcSP�~}�w����UVS�33\�Qf%����e���zIJN2m�k��\���I�S��
�SNR74:D��V����7��G��˗�a�O�N6?�<�ӌ�<��l&.N�Ix���s8�ǰH�>�`��z��!����ߟ�7��M���������r+12^�)3��<��^dx�~5��ů����@%��k�����V��]D{w�q�`�M�y��a�����t�@�6��Ӟ��z�����l���C�xE���ށZ �$�)K*���:���G�x�&[b�����/u��4r���g�1l3��>��Kg����oS�����t�wU 0A���������s���Zq��z�������Zz
�M`�d���V�,�X�9�{6�kq;��Y�w�ܿߧ�k0���{����BSj��1����XY ��R��	�o;�N������cm��SO��*�^95�]ϛl'�C0K�a��? ל���9��'O���FӅ�y� 6(���[zp��Bx�N�/����s�xG�GH�t��\�m���u=�v�c�u�1 VD�ZPR������E�{2i���/�n���?l�T��N���������\�r��h��A�w� ��M2������p�p��`��f3fR�;��Lǰ�C��p�q�7N��dPp�,z�s�N霋�v�h��"��b����[�1��߳��[H]�q����ʀގ�a}MMʶ�#�����Sx�����	��~!51]�I�K�Ӂ�H�>�;�у�����dDt�f'&��\�W�;�p=m��T4
Y��:N%`c�)f��{��]�As�I|_���X��,�CO�>���Gp��UX,W$��n�\����BX {�<��p�.��	��\��ޜ����̇��>��?�����C�p�$�������{(.��3Xh���(�O���w�i凗��|�`P�
�:lbh5`o�������Wޓ�^�K 崎�6\��z��?� d�@� Ԧuh�+}��o�SV,����_/�-=8�1i{o9(�Q�m�hlʀ�;g$>���� bYn�՘;����6�l�еt9`�&>�.�ԐD�~H�֕�?r���h�������0텧��1]�����8�^ý���_����xR�d���xv
�l�tfkL����B��:H�߾}ۯ=���}�(�;(���S����m��Ӧ�fd\�<�r�Dc��w4t5�ڻ��?#�2v���`��dA���m渆�	�#2a�v�/�=��n������)�w��������te�z�^���.H��Z6���3(cc�j� �qX�G�TN�KڣB�'E�Mm�$�&r����5�?-�K���e�1�F�Mp�ɏ�col<��))�=ȇ�wf�0^��˃������3�fg0�~�Ν�!<^����S8�W0��ɓq���^-!w�-W+����������z��d�_l�x�&)v��2�~��)��m���J(��I�v[;��8W�S���2�5������������C/�8w����K�|;�g,��ʀ/��������҃�����p��
8sQu����H4�a�N�X�2�*H\�:�@�Ƿ��k!,(a��e���Ҙ�M;��.��ZUT��_.��%0'��	�6�S.�y�9䡢�\9c�\�tq�3�����0�O`�;В�a�����޹�{��x����� ��ā<�/Ls����{���ٳ����wa�X�u*x����IyǦ��)����X2��+�!߁:B,@LC
�8T�1�!�W�	�28�a�@�{�0Y�v�x!s(����A���Eώ �����$\#��˗/�LV�{廆@�9��@w�i�����d�e<N�e�e'�Q�$@�7��@�?_��t4���i�t�I�)�j��J�}��y;%z��m����������k M�^�{�H��;n��<\�řz2�9�J����	Ź4e�e�ɿT���*�yI�?��o>::��?��$�8:x�Fg0Ha+�[����|�� .^�x}�¯q�+�,����4�������C5p
���B��ɧS�e��}�q�O�{��&<�=ۊ�X�H�%yXǐU#���>ݫfz�5T�F��uS�8� {R�kH��x��x}
���l���v�q���w����O�%Z��a�G`�����upo?;;��|�z��N���ŋg~�Y���D--�d�.�9����ez����9�ݜ���dG�w��amj٢�y'ƍ�4�i��3�5+Rٙ�F�� [y��QW��1/C+}	f4�F���e����ϿKP���;w�]q��5�cAۧG�^83Y��(�_������(_@�6w�d�S1X90qk�ݣ5�����kp�Fש0�G�P aY������_�1��ۃ�j���� ayx�5L�O8�˟����O��i�7�Y�8�i�g�D��J�W2�4�rh���qџ6UR�y��x:7+�������x4��������~z�������M�>�9�K�����u�TjM��{�;!=8�rY���Q�zO봚j�,	 �hϰXk�x:�A����ѝ>�]mE�~DV��������t�.�.�����j#�����Ũ�pa�B�^���ܛ���Kc� s�k	6�e!�����M����<s�d�_�,q�7N<�lP��A����]������ ��8�Kq`)��]���
��C�Y�mM�w}��Q&&��:U�US:z{� T֧L�2<o���[�Y��Vx+������+qmc:��kN���.��?��k8!��ųx[��~���8*i2�I�-t�e��'[.��:Mc(�k�#�S��Ϸ���0�AЌ:�Q����p?�h��~[���Ҁ�v"�'�M�=��TzU��}:��GQ�!�a� �$;��p�]�:x�9�.�:�O�,��ו�s8-��tw�rx�<���ˀ�I�r,�48�6vu��F��z��]��5Nu�i�D�+^��z���r���2mk��2��|,p"�k�'��:I�����q10L����uN����#8;?�|��t��S_t
1�/
mP��	̕d�h�11%��nbWb�{�n��ɶ���/h|�ѼV������}9��≥M��jW�'7����FA����e�=��2��RH�C��L��7Y�:@��u2N\��r�S����{��/��tN�1�*Ew�h/��(œ��{l�/M�ӧo�9��|
n�y�C$M2��--lU`�p�INs$(�.tb�畗�4��k�(����&h[����2,��i�G}]��.V�6ۀ2ם�v��(�h��1��]8�w���7+��Y�`�\�|6�d�I�� ��Q�;��������z�~���.H��}\�Y�	ݓa���P�vc\4����QI� \�p-vF�赼i�%�#;����O-�|ǃ��SEW�T�iq�����gBF�.&g���.��>w�d�D��:��A��~��3wyw�����
�/�[B6��Z~Z��j1�O3.|e$+�K��%������;�6UP,9ȗ&f$���uJ�W8�������t'���  ��IDAT�0��m�/=OM��� P��'X�a2��<����C����w��͛�ͮW��L��5���Jm��;%`ڰ��e��'_#����6&]�ŀN�����hs�ag�>��t��p��F��Q���I�/f�%8i���ϻAW�v+�ӆp 3������9 �1���)�7Ҟ���b��t���ģ��_��t~��
rws��:A�k7\:/_��ã�V��Ip�1��)�$���=�mp#��bPkR7���H��A c�$�����"����R�5	�~pW����?�v��X����T%��/��!h
����zZힼ�j�&k�U/�!=8�r	s�|aX��mv���F�Z�Ј�=�G���7;kͨh�A{�����K�]K���Y�|Β��,Sm1�>v_�_>+�w��˿��7���Ւ!8}s4�Ý#�K�%����-,d�Qؚ���}�d��������������g0�}X���������O����|�EGo�e��2�p�J��@�T��V K)��N+V�f��� �o��������:��7��5�he%��~7� äI�6�:�O��r�J��q�d�7��$Q;�>
�ʼ�)J��EU�% ������^vWzp���^��h��%��6���ڢ9ٱw9̬m��;k�ii�4�/��H�yv����Ƅ����c�FWI���.���N��3=�#߷�z���яxѰ�1A��"Sru�����x@2t�b
8.^�*�ʍ�3L�ۋ��%˰��}[���� �]ڃ�^�
C?�A����x����
#V0&�t��� y�M�������5�X�� 4/��t�@�����J�hX�ʊ�Y~@��xSX�u�����{�`6;���38<����U����I�~R������ڡ���V%�"��;҃�-�6	�Ԫ����ЈJvB�嶶�Ō����������;���j�O��Nͨ˴c#�6#��Q��5:�w֒��ұ �,�P.����A�_��>���~;���Ňۇ�)\>�B:X�l��,F�>M�@��^>�S;Y���8]�����<���#��Y�0ڟ@r>�@f�Fة��ɓ�0s �3p'g��%A�&��'��a;IKǂ���ʵY���Sˌv�G�}8d��r�wRk���v���5V��qk;�\k�*�#�0!�0��:�u�z��p~v�w����s5v�(L� Нϗ�X:qzv>+O���v�˄;#�X�8Z��)�/�
:{�>����H�|�c/�!6��_���H1���pO�}k䫱*u]t���Z:���F�\K'�W1��K(�N (���ׯ_��ds�ұ	<���`������3������$A��%�$ΐ�a�&�����rvϫ�M�%p�n�����w�7��C_�qm��q�Ѕ}qnRz]mnö�0Vo����jq�/㶘��,V��?+��Z읶jͼTkk\�_��Ϟ���ߵ�Sq��,��|������O`�X�Ӯ<x�A
z"�)D~��V���O7ke���IN�\�|�djǅ�uv�\$�{�����p�Q�`(z��u��`����m#O���G���g�|����Pǟ����_��_{o�~�:�8��g�gp|6�#-'0
��,�*�Q-r��P��`��a���tx?v���!g�`����L��gO��G?�7�}0Nk�.W�/ف�g��oSN��kL�uЗ�����c�����-�,cW����>�|H�.�@�� �Q���߫ |L�9d1p��O�S���W�\��܁�l����g���s���O����� ���_�?������a�0��>�8Q��E����������dGĳ�IBS��ѹi�Jb����0��۝9l$ZG��i(�#�;5#�M���2�<~�X�s�Z�W��wL�>t���Q/
�7n��[����я~��@vezf�>��S�f��!9�����`�Ң.V.�� �Ma�a�Z�,]y�N`���8t���ａ{�w�ŋW�>�83 ���C�E�3cm����l��i���l�ug`z�[�}�wH;ꀧ��c���e��6h���Jˋp��O�-q�4N��0���~�X��-a^ƣ����}pp�_�.�k���T�7M��o�=�z�dץ'; 	��T��9�A��p���'�"P��@4Pc�y_m�Y����v�����s�����"�GMgnt-���I�4)LV��	�����>��#���0��c[�S$C��_or��"�i��&��ك���}�fy (���f�������6O��x�������|ۯ[���)�S?��Ȃnaf�外�w�Xe��,  ݘ4	���t�ξ���0��zB`r4�@��ص����x3َ)��_l'''��\�|�}?��o����CFC��G��Hl�H _�pɯq"���<�8uD;�x����^vGzp�R[sQ�.�1��aR���d	b�5FE>�u�������S���$�ɪxd��t�Ia��N1�E�S�/��h�H��  C��g�����/�K�νwކ�x�ד���%+��:ۈq�j��:�?��{u-�DZL7�E���|��d4��ӏ?�O<�{w��������$���>�|U��;,�|1{�yQNy� �S]�k{hv�^���+����f/yKC�jJ-�����zk����2ٶ���	��H<��p7o��;�p+12'����C �ru�>Q0�,Ă�Ow����>�>]��nJN�\���$��K�E�{�n^ơ���j�;k�����L/|��˟��_��ROC21Z���eD����-�Ca�G�)Ь.�EA���� <��~ܹ{��}L�~��2_ �!A����5��8�n�r����`.�Pٓ��|��?��GO���K.�w`��E�9Lx��
�Np-K� (-�IB�h�����H��}uj�"��x�~�rEoL��Kڰ�v�.m��u�j<�IR9���!^r՟�� c2�<��8C���]:�n���`Y7\-��Y#�B��T�ݐ��$eO��: Ѐ��^,G����|�9,]K�9�c�����O��ҏܷK}��t�:"�f|,�"ӎy���&4����n��N�ړ������7�¥KW`4�z���@�哼���G�Hɣ�ywO����9<��cx��A�v�'�TY��X��ne�&~�g�W�$5C$�,(�2�r ��~�(C�np�J@���H}����5�����Ә+�G��R~Wْ���n��6��S��|��,P���'Xv8U��Ӫv��ˍ�.�O��!�3�������d��;aK�$6����G�,|��	�Hp����.��%$�����Fx�rT.)�QQ�bD��Qd�[Oљf��Z�k�?|ɯ��%<����*��H��Je������+����՘��lZzT�;��?r�vc,=%��M�܋/�������/�6Ѓ�.��eXg��]	e��Í����'��O�³�O���5\�xnݺ�Gҋ�*@��9�2��Z��9P	 i�ح��֯%	�# ?��ήU,/u��ʓ�}��5k5�sm��c۳�i��� 1m�򖳩-l�����|�Y����r|��c�|�P霔�-����v��j�� ��?]��ɖ�`0Ƀ��b�@q	��8� ��IZ�ya�����2�/��d��:��cGeD�Q^�J�B�;�ʘ�A��E�ْ����n4���4r��+�sB�ƹ5�H3Ijɠ(�$�
�%a�똃^�����E�r��m"p��˗�����.�]�qpQ��AA ��חd�tk6�3�����pW�ހ�ox&�{�<$pk�	����My�rq���k��Q�TN���m��HF�^����vR�##Q{%iӰƀO_�z��Ƥ�w��̣�J�vyNiȝg�t�2̪�c�$���~"�gt��u���1��l���d'$m�9ʌ�>d�&��e�c�F5ݬ����S��y>��ͧB��z؊��Z�ۆ1���T��5]��`ȃ!��S���ǥK�����D�9<z��O� h	'�Nʵ��d_��Gc�g����.����^p�U�1	.��u\M�Y��o��������5���t���ڮ�j7$|���ی�|���Bks`�@��OC�+~OT��>4���҃���?��θA�o�㏇���^a��c--�C���[���/�����?��X--뾦���(;ƒ�(+#��C�/� \Ј���bYtK�^?�Y����@��\�x���t�AH�?<p�pR����@ڔIsbF,�@+Y6#(�[�T�m�I[V��QVzܭ@�xy��;�']�铎İ4}����D�l���d�%�9�{i���$m�%m`G!v1*1��VS?͈4���2
�F�R�룅�"����k���ͫu)V�1�~#����P����˞!�`-�G��F|PdJ��U�H�5�{�֧R���Z`�O�~h̆UV�~�uO�U{�$�֘rjmʆ>�T�g���a��qQ|<��n�����c,�E�U�<��.HN�\r|��{X�ɥ��*���c���fx-m�P�Ӕ�s�6���Z�K�����rG������a���zK�L@�$�֣ ���+R��B���o��`i��Ik��\"���Xi5'����/M?���p �}ߤ=w�u�ݦk��wZ�]ǙMG-�i��l���d�e0��7֩��FQ���?ޱP	`��(l�s���4�<N�t�/��<�{2��H[���9҅▋	e<�	��լs}
��:Ѣ�x������?βT �2}�r���ڦ�nx�h��떷�6� N4gy�����$2��#�����i6Y6<~���=yĀ�g��V����ddh��e��iKNvL�АH@��l6e�b$6�lQ�F��C�i���a���N�{9�B�.��L��d�y'��O�>���J�*'��{�>���la�V��S���A ���p�q��|��3,�2�4A�BQ(�5b�����ΩP�l������L;V�M�t�$��c�š={�-�#J�]I�%�>�@��+����w�S=0�m��ɖKz�rAl�S�t\�P�V�ïi�α�����-���D�^�����ڲ��HY���ʓ��������s���{����!��+���x	X�����H�_A�r(|ufJ}�	 ��ؕF��hc�L�6*G�16@�n-.��v ��֍�0R�.�Xޓy�?k*X{��`��;��5M��0����HNvD����^^ޡHJ���j�-j��S)��s�S����K9�Fs���� ��������k�9���� ����(�x�X+m�A>����y"�(����X��8�Z�r���Q��SQ�+Iu���m!0)kS�ңneڼ|� �ߚ�՘띰|�P<|g�F8��ΐSN���qsР�Ʌ�ˁ	�ֳ�Xi���!���,�����vz���҃�-��p�SW_��c&�3���K�/��8c�BlT��Yi��gx�4�ޱ��qpf���K���V�<�p?8��F�<]�sT�N��A��D��B,�kc�!����!��f޵tQ��>m 5��v*�o{���@˻��ԙ�UV�h˿��Ɂ�,A�Jb�{>V.1 ����҃�m�%x��m4�O-�ˈ����,�:϶�k� �/��bE���\/��*�@�:�Q(������, �RF�Ӄ��.?����|�6��f<���~����(;�~7)�$�.ƶ-Lp7����v]c�8�A��&�x�[�S��ma^o��`��%zYV�����d�%���:�bu�l��j�������Ml�$�ϛ��7�׌[����	������Sw-���H�!�����r�� ��u=�3��V�3���Ϯ�P�����3����~|�<4�Z�� �J�ߋ�.i{�����k�-@n��Ұ@z�6��+�X|��NHN�\��a�m��:j�uTS|����Vǥ=���d�1u��/����N������&Hk�Չ�+��k�a�:�z8)�J����4�e8e�ǀg�N�n\�� ]ڡ�f e�h�7�w��5�ß�֥X�!ô�~��ńhi�]�������2A�*n�^{�����@b���0�N�άitک���L��]GsF>rn�	��a��Q[g�pk`DOWө���x����}^����%A��˶r�F���[L�!��Tk;�;k[��,�e�M�lH�t�]��̅/pF������aL��s����nIN�\�9z�������x@��k:c�I`"��k3,ݬQ�������]�XG,�4`V��V�V�G������`��	_�mZƴ����@���d�,`*���O;�\Q���;����a�������V�W�x�+�֮�m��s����^�_zp��2�Hg��wcB�kи��w�84O�1ce�!�C�j��0�qH�m�P�F�U���	ʚ�T��直�4&�<)����D1@ [��X�<i�[�S_3�@i��AD�F8N,֢-�.��r���۔�?jS�X��@��m�>b`M��^d%���n�)���X�}���^vGzp�����m�Sl3�3m %�4������&�-�As`�Zwj�z����l�z���aK#L#JN,C�)��4t�YT^!H����C�ٕ��up�&ۊ�i�G[mO}��;�쎃�莿�<�|�2w���I�3�R��!�F����|��K����O��V_�ұ�˞A�]��ɖ�t:,N%�#u��7�<��w�R4#�u�1#���p)/�>�Qp -��YP���������̰�O��:0f��Cy'Gd��G�� �ŷ��H����Ի����l*C���jx����4�z(��|U�y�RX������,9��S�\�>��<_�����:{"��l���K������(�<�冕�"�K~M�h9��kB���g�� �_ֻ.��h<�,%��#�.L�+ğ���?o׽���d�w�� "��Q	�T�ҤI1��B�X��x�+?%9�V+;F+�����:G��ޤ�)>J�t��7R ���V���7��d�����4��v� ��"��L��D�Vz�د����n1Vڈ^�Xyhu�Y����/����@L��7}W�r� ��������	>��G'�"=8�rYҬ3@mI˨XN��s!|�P�b�������RA�>�:�f� h����YԀ���c����{�OK�M!u�y+����e���w�&ۀI�t��2Қ�m �z�:�$x����x��ck��@�����n���� &ɉ�l�I�l[���vHNvX���8�\U�1��N�{'��G�1l P1��!�����z����6��w�*���>k��Ȑ_慎��ĥu��kC��hm���m�t+@k�#�b��>+�Ʈ�t�x5@c�e�{Ǭ�x�q� ���l�-mMbqX�6����j�^vGzp��2�b����e	J$�j�.���ؐ�\��]�6�oh�-��&m̍f��]�z��&ݫ���t�⍉6�*m�6&��.]|�h�wաn@�����.iX@#�Iل=��C��&YK����.J���X�M ���ŔXqЀ�#�-=8�r�����ͦ8ԗ��'�*uy�ca����ϗʆ��4�2^(�`0�3ԍn��ԯ�v8��y}�\��7���u�Z]X��b'b:P\��9-��u��EX�����X����9����0+=���ћ�E��kV�m�H��]�ү�w��c���^vGzp��2m0|`�����[�D,=���Gh�ʨ��5M���C�����A<[7
] ����&�o�&o3����z�,]�����M c��fie1 ��iL��^yY��c�]�ĀG�oK�-X�)��dȲ��igO/�-=8�r��X�7GO�t׎��L����j
E�:��/��k�H�ɚh�rk��cF���&��h���:���|�OyÅ�|km[�eZ<=�~3l{�ҀH;�ԝ���Z���%�օlm�B#�i]p�|�ҷ8��	oo16�p�e��'[/�]')z�xH�Q�ۇ7�a�w�3��ˎ�+{`uı�\ꫥ��|%�����k���	��"ipc����4��IT��������|>��c��c����ph:�ڗՎ�LR8Ȓ�:���:�s�i��vj�>��i])2�ls\G����m[;���uP��vJN�^F�����Ԯ7,³#}G'G��EN	TF�S��S�0N�H#&Ok�`�S��r��hy�i�02w�3B���'OY�A��h�x�h���y��z�F#��f>��t�?с��Q���܎�c�s�<~�NNN
�oU~0N�C	q�e^H7�X:�L`�ZE������0��U�=����겍���Yi��A3� j�ȴ�}��7�g�Pyȝ`Tw��{/ư�M�c��1��)]�`R�%��uQ�~Vg7�'[.�=ߌ3VD3\m=���2��Uhc�5y�2$<��x�^iz�G���s�a������W��dgO���b�h�O�F��G���ϟ?����\���e�^�
�/_L�@C��a�{{{e�������H<V>�$` ��Q��t$@�@Z����	�?�"�.�R'��_��<]�y������ߣ)?4T�m� HS�����e�e��';"�yYK�y/�6�2�J�kF�����`�x^�tc����� ����zH��˄�d��-&��	̬��a����ğ�Q1|�L>���]y��!<}��
4N�w��%oxH����/^��g����޺	�o߮�ֹ�B[�Xս>5���@[k#u�t��I'���/�^�o������Q|s6��8�#bA8�Dl]�	}���z�O>M�V>� ť�'��˟���d$�U�	�U�Kl0 �C�X������ߦ�IY�A�e��qt14։�2�"�K屶q�+%���2���L-|�Lp���ק� �@�q��u6��a�!!C��Ǹ�	AЁ����'���?t��-�2|Yӿj��uˈ�����d�j�\�*ӑ��tI�<tMG���ii����sh��� [9�����%��ڮՖ���M�4z���҃����ƜX�[cN�69ʱhi�fnվ�#L��x������#V��^���ճ�v�����6���`��X�����Ξ<}�<����p��E��7��ץ ��?Z���.����C��ի���9�����}�iӺ��B,�ȣ���(4&Cc$�J۹WrJF˷�$���($Ğ����XxKF�����+�Լ��S�^�\zp��e����.c�ب%6�`M�g-`��]-�Y��~��iMG(��i�H�AOܠ��#٣X�1J^3�����
'��x�;�&>��w���lɕ+W<�kdp�C6ҍ�~bW�m988� ����<@�)!M/�8u�9]�]`k{F�[����XF���1�c�Y��w��j~��Yb��BW�s���V����]����bu{���ɖ�x�od�	�h/>7hVg�Fo:��B9�pZ'^��������ȋ ?��bo4�u��5M?��j����/b���ТV4(8����������1����A �7Jd�h=B��������˧�~�A
�C��i���3��3����-=�~״)�4]� ��F�bﺰDZ���h*���P� PJ
�j���Q<]�Ե+��e{�'; a�����ىQ�"_xi(+×��#E�Oq�^�/Ӄ�:���_����+nƠi��r�t��C�X4��Ɨ�,�_�-&��"PA@�~��'����������iQ�_��$�e^'�_k�g�<�l\#��]>�%��#�y�_H�����:C7��xٚ�b˵e�fuaAd۳����l�M	��(]��M,&��#�� �����:יv���׿� �ƍ�� g:���;v�0a� �r�{���իW~zO.��� x�b�i�AQ/�%=8�)��0�g�s 2U�Cs��{�G�Ӧk�l�ig�;�c5���I���
JdR^)���l�WY�,/9��>��ZMqꌍ�Ā\W�7d��_0ܣGa6;�o}��~:g�@.�ERX�fa4�/����5Iq;�gh�\N�Ȫ$�Vx���#g\��[�o9@2�_��W���3��moܲ��\�[�Tm:��V��[K��ueִ�:7�O�b�3����^�iÐ�8�o%�|X�?�GcWQ�^&���9��׿�K��O��K 3�������}���z���w�?����QX�B��@zZ ��z���ɖ��Ↄ���0ᷘ��roh��Em��a����Ъ�
�!�h����#Uީ��*�F���U+�QO�:��1)�������ŕ��?
v���Q��4��P*E�y�_�%H!ݪ�WFW�(#wi0���RlV r7����� ���w��w��m���ԇbR���4n���U6���!n�����`F��8��¯= ɝ[���\���c�\�z>��7���������pt��K���b�<�	��X����]�{ ˀ�z��Ǝ�#���I5@H���m�ҧ����:��u,'y1fG�Q��X���JP���/�v�A�<���Sx��Sߎ�IY�]Xa��wvv��\[Y,g�����5�lVl ��μ�N����¶҃�-\s���^X�	bF���k1�|lj!&޸f�&<�J��<dZ�yR�+�)��΍[M�f����������%c���O�|��w���{�y@uvv�B
C���9�3H]�ϖ0�\D����kב�B��ـ��y���F��)���8���k~>��hn޸�F�7�����7�{6e���0� z]+4�a�9E�VG��׵�VY�i���&1�B��R�K��om�J�=L6��_��������`�������ז����"�~JS�h4 �£�7I�\���pz�z��ɖK����:jn�5�x<�'w�%NOqG��F����i��E14���}o����kɫqf�4DG���6u�Yw5�T��_��_zÂ[~W˅����L�/�`����U�ё#��hx=��Mr7bN�`��#�=��&Gk��;��*���3%�r�����u�]�������wn���a'PZ(�A���|Q0=U���x��@�̛,{j۲^M��¶�9�W����J�GKK3���׭�]O���p���������Wf��9��ׯ߀������������z����_�����=|�;߅K��xЛ$�"�z�X����pm�^�_zp�5�)��/bqp� �&����-@g�,��\���2�"��X%����!譁���OꍒB�Б���Jꭍ��i�kȚ��7��.�1����F�����ܽ<��W�a=_��E�W����5\�8�!R�X���-Vp�@���fo�t����r ����VȈ�����{7���˗����p��w��x2ϖ�w�x �!�I;�#�p�iӘk��i�o���������>ڀ!��|��Kϵk��Ot����-2I�������N�a����9:��ٔK�.��ɓlR�eӘ@�*q}H�f�88��`z�z��ɖN�$���1 �{]���[ƕƘ��G2<Xl��;X����*�9'e���n��܊�F�5�T�A�M���9��F��|��l*�e�d,�5��7�Y�"�ũN�(9��{K�se��{�ptx��1|�@��q�.�ِ��4�����b�dW����ԯS9sF��j�����ҹ+��)��[߁��_���>py��|-C};�p}��I�˫%s%ۆ�|و�mm���g�i�ؠ"&_f�G�$P��D�A��";��/�j^�:v�eW�\w�^���Ϝ�4N���iӲrP�l��<Z�g/�+=8���b�]�:��u ��1>Bo�(	@����S���	g�H_\7˽����z)�/<�HC�c`��ۚ�:1�{���Q-j��N�d���x��� _,��@ك�d���������ׯ`=B6ރc�/��d{	\��Kesxs�­/;�;9F^��b��܂���֖�n)����4YC���f��u���VNڈ���5$X ����7�m,�������5��� �����8����cx��YX��¿x�=z�hX;5vm���;0ʷ3Q����[��gQ�~��nHNv@p�e�k�A$��F����F�ʸu ���yK��vsꆀ��c�b�l%��ɠ�,
�'	�E��T[�����V9��:c�F�[��FJ� ,��h�\ʃ�54�A2�� �1�`�t�)�7oN�8���(�t9��Nf��2ۇ�,�}=�v��|��ڵ�Gǧ��zN���N��2�8f�d�$�;q�$�p�i�ٲ̍�s�hP]��muG�e[笚l7�3o�a��Z=����࡭mn
P��\3���x<�cq�>��a�=���p�#';vp����Dꭁ�[�z>����l��;�L�f�g��L[�؅����g�hv)m@���O]�Q�2=>Z���y�Qe�ő HH��_�Q�Y���F�plm�|��壕��[~���ܵC@%�c�l ����5�x���+xz���'�7q@�xo����2��p��q�)��gg���4N�)�8I&�۾OG|8����i[�I��<�_LP+��X���=�����r��c푀p��#��M�������>����B���&����6�^~�7:�N/���w�s=�K�b�!���jX �a��&������l�,�rʩ���Μ2ȼ��Ӗt���F�];�����b74�Cy�-�|Li<e\�s]�[�6���-�N��{+J9�������7+x�:��G0�N�ǯV�\-#�P���.�>�pz準��Y
�|>�%��܈z0�lp�?W8�㒘���v��%��v�!����ʀX�����嶩h�V�V�]�E������Ip#�ڔ=�q�<h�������S�]�_�x�ؕ���k�n:�r�<㤃��F�?0���ݐ�l��� �^VM���O�%�hm���Fn�)�:(���:j9=�Ӭ�J�Íu���F��ݑ,F���)�X3Fr��4.t���iއR?l���Q����1��=x3{��/���>\w#��N�^�ځ��3���f���d5���e� O2v $�B�e�v��C?\ӲZ�4R��p0�E>��	����|u+m�$��e�O�Ei[��ť鑀^�x�����n� _�, ��o�{v~��\����
h�w�J���@�J6�ڃ�]���l�JJ:�:̶sh��]��N��`4G��!�q��(�57�Rx^ێp'����X	��4e�,;fX,�ȟ��0�v���I� }�Z���7/¥�k8��^�����#h&��p��xsr
�O38O/���
��)d��#n2�@-�V�b����gK�˕?�e=s�@; s�l�m���� ��[Lb`T�.�#�##lF��%����n1	*���T�}��m���k]Oܵ���sx��$�[��AP��=B�[��)�<���gz�=��ɮH���N��u���D���*M�h���6�Q��y�hZ����_�vb���*Ya�ߖѠ��|�@�;�"$h`���tp�I��	��&0�}�we����#��4���g��ho�=��j����`캖�����<��|��� ��櫙���w��ho��g(��=�e��ݚ;В�mɒp8c)��0b4FM��T�V6a��	�ii�Zun1.����E�|(\�|X�J�H����LO�a���>���b|p���LBϰ</���a�Tg�������=҃�-�p�tzC}עо�6�O����G
96m�����YjI��L����A����.��e<������߅9�t��Ĕ���z������3�`˧Q,B�-W�����w�� I/�x�f	����#�8�����0�2����/����N�q�d1:�sp�N�t��w���Q�A�c:�o�����N�A�~k1vU��は� i�R�(�I�>��A,��-ȶ�8 �k2_�7g��Ca�t(���Ǫ@���ܕ������?e�x�l�ѰH�����@Q�g鶁 ��G����d����!:�M����PG�wX��F��0$�F3��!�
�q��h�+u���X��|�tT���1�bLڀ��,��b`�K���mS�=Ap��a��?�y�g�X���G���t~������C8Φ�L���fDL���w������2��z����|
s6�fsX���/@��}��
��ɣ�᭻o9�����<���Cl�&���_������ۘ��W[]��)�w�Ŧa$h� U�E����I0������\-���[!�����޽=�J��7�B�[�Ǔ�I8	���-zn�$X/�����҃�-�2z���e�D�iF��(�_���;!����X�F��5@@�!ob�Ph�c��ؒ6�����+����_�x���������/�����_��ۀWkdOpW͡?qx�Z@��ʁ�Yz��o�ެ�M�3׳L@; r 0ރ�_�]��=3u�&~{06ۣ��B	���������9,�F�Q����4�$-oeٗi�2��0hm��Ϫ�'�������3PKOX��%�����s�.V��;rp��^aQ^�>��������?�:D�M�� %\K؀(��$��dz��ݔ��tz]Y��4�>N���X�l�	|�U����u�ִN-|��~`X�h2�'���������S8�(�?�e:j^��������_��_�����s,�5�@��2w`c����܁� �h�/�\: s�Q�=_���i��V����y�	FC4V�y1]��g�_�b>��׮�����D�(kg�3l[����]�Dc�31�)Ӵ�C�/u�����@gc�1��ƞ�4֫�!�F�޽{������������	z�]�3x���@*F��.pkyN;y�rU�\�Nd_������d˥<��<���c
�NP���@Q�~[a�b`*U]ט+O���!��yG��d>bb�ry~�L��ã���N�h�t]��x��\�|��S�V��>m�#�!�IZl9F�c������p�t2�F.����e�[\:����N�&~�ɇ~�����a�$dשׂ���0���+���˿�I��_��(�C�}h�v����ӧ��M	���7O�F�jȔW���w� 8999���^:�>�=�<1'���E�>����"�f9���l������@�/yyͯ���|(����kܔ�)�"��l��.��OBG��"�2�s��(���I��&ŉ�yB}�D�WqLX^�
�reXʧ��d|�?7 |�חy��B;�������^���������WyL��@p�;v�l�������>{w���lz'�N���E���&�F��C���=�;j��<�ˋ:�uN�v�j�2��C<~�N�A��?�1�~}ⷡ��P���蘔2ߔ窬�dm���z�7�>/6d�ˤ�/�օ,��ÑO�CE/���C���}/�����gR���z�\���Ӭ�^�G�>�k< O����X=�ϰP6���{�}��^�>�ۀ��ݒ��H&��V����DiR��zG:��oe}h���fds�ι�Py�B֣��Ȕ�#g�J�pMW��~�c��qzA���S-<��E��35mMȲ�XzT�A{�����C|�.�Ez��͛~J��O�u׮]�uD#]�Ce��-�a�q��"�T�IYgشpj�x���������g�ܻ{ϵǡ3`3�΄�.�h�4�kc��w#���w�V��&^-����$*�`����i����+<��{R����z�|�p]��s��}��\�������;�?�?q�Ù;�� �����W�P��#V[��nIN�\�Cl�'�$�  �2~ ��:�M ����|V���c�A5���J�ƾ9Ҥ�5/�����Q����-F�[l�U��N�P���y����w����gx�ɧ0M�⅋� -�V�aZ��7���R5�������挜1C7��^�r�_��kp�KV�e!���(uc��mN��ŧե<���MV�M���W>����&m�b����^��g���/V��:����g~rA�+�&�Vp�,����,[���b���?�xG�'[.x&
��~�]v��0�A����!I��$F?�u�����4҉��1<��A�:Mi@�5��EKw���cF�7��8�>�^р�s�ڹ~�:|�;߅_��W��G�ݻw����8�C�Ne�i�S�(���1>��3�{����8�����D�̚eT����MF��3y��@)�R&��F����nMU�DU�}�
h*������	�������d�g�g��a,���u�;-_�{�4��z�z��ɖK8[��@C�f�L�EE�uteGPK�����X�Sxˠ��&���9��1���Dcf�x�`,��թ�$�V���TF-��	~"�x��w���o}~��_�o�[x��w�ҥKި�:L�z��g��Lwu|���>\��+�Dd���E��Ev���˰1� f�k��Tk9��n,P;���#	N�8�NL.֛�u<��ǣǏ�ѣϽ�X\o�[�_�z�u��������� Jf��C^�A����a*�.HNvD�n�bXl�R��gc�` �<a�:1��N3$\w��u�$��Fc��P�Y-nM_~�3_:�����oc��b|4��Q-m�DA��~�;P������A
���E������qWΓ'O���>�����s�3���F�P�i��C�}��%��S���B�{]�v]����%�W�8�y#��I�|6���cݍ�<8:�� /_Ë�/���׾N�>ƃ���I8 P?�O�_�]mn?��z����Hؒ�%\R�Se�*�΢~-�D3�]��6:���Y���yc�M@��n��X�K�p��L�ݛ�3�A���A	�A�E�hLp��A�i��O��Oރ,n9�r��rLj�4H(�~��ӧ~|}��s�!�*։���� D���e�=6�BS���� ��<v����OfH����"4з�?�r{��w���w���Pvx.R1��BN�P�oƩβ�~�^Z^{��� =8�r��I^,��,��K/��QSO�K=.�)[�Jy���f�c!�ј�����g�4$r��r	.�X7.r!s�i���2xR���l6� coo�o�D��;j���<�N��"V����'�x&�!����wrm�����Ha#���[o�SHh�0<��b���w���{c��iϻ�_ft�1��1�X1����3cg���ډ.���i ;��_k���F1Q>p�+?�	A
�Ú�ýw�vuy�/r�:��װ-�w\�d9{��k�K��j� �^�Gzp�CbuB�#��%�oGL�+o>�k�<i�3��O��n�N�M7ҥ7؆�3�s�:�T��FS�X�%�w��_xq���7�Z�H�Q�6^õ(x��t�����|��#/�׃��ֳ��=~G��KP�&]�T�g�m�3��Ѐ����9V����ku�wT��1 ��X�'}�g�Ti�j�o2u�7+Y>tO�e�Z�b�ăU���;w<���\d]�2僣*�s�ƻc�z�.��ɎIxYu�ۼ��s��I�)��A#�>?4cMN�*ˎG<����Q�5����NZ���e��Os���.��r��W�Q�m�Z~ �� tf�l�0�v���&2X�>����N�!�x���YBlU�q�y�⮌���X�UF6kL��z �� ���)5	eZ��$�=��� �%[�B����G��_��O�K\���<2	m���k3�ypއfA�b���l'�)<x�)��g?����Ç��?��/|�5GȜഏ�Z�4�}�δ>��.���(_!L*�HN�^f'l�h� c><dg�`R��<5m�"�4n̐3�D>O�4`c�6�4p�C�Q}3�u���8t�1%MOE[@Pq�Mj���ԍb;E���-󣕽�b5��6�¶����1#���R�ԧ3�4���'�^[�y���$H)�9���|6������كpzzϞ=� e4z'k��s��������J�ø�5�'��x�ƌ�th�MIK{�ٓ]��l�L&*q�Yt��Ռ���e�e��1��㬏����2uf'ׁqhv��F�)�46*m���z��c�:��7���u�4��x��K�a�ƍ�7椫���@� ��,e;�:k�,�Ɓp�M�jZ5]:dZk7�៼,�]�5�5��:Ï��|�
~�����t'���88��!���ys�@��Ǉ �pq5���:RZ��6i�I��Z/�҃���n{�������ykqP���JR_w"Ӕ�H�Ҭ�%k��A��1Pѵ��AwZg�5N2����\=��WEèIU��8� b�l�����3ڽn�Dg��S˗�%�S&2o����h���n社'��|J	\��+�tz ��1\�~ӯ9�np��(�a\L����H(��Q�ۯ�"Y�<cLW�z���ɮH�gcd�ҙkh"�l&��h�}jS(j��.b���6��~K�W��d��<��֨���v�t��JYq�5�-�^�Z]k����8H���C��!c��lBi�c�u_/�:�t� ��<��F�_ˁ�ܹs� J������b�5
m7'=2N�y�k{ha|�ꨗ��|��F*�!�Q�d��h\��G{F��m����`x���t��O�]��b9���I�~Fx-�.F���3>���"��e�g1�y9v��c�v�ޞW�m"}�w�Y��+�@�ZX�&��D,���Ud���<�S\++S�@���wzz���r4!�)K�y�Aקt�
2(�?�+�u=}m�I�o���������d�e6�V��83���}�y`fy���]�e�eMb �w�2n-~��s�|Ĩ��s��r�ʮ���Gc��ӛ��!�k�0m:��U�tm�Fzk�5�Y�o}a3�mc2���eҥ� ��+�������;s�%s��Y�Y��%uG���d"���y���Y�R���d~9�˟���d�%/�k��ѹ5B�=aXڧ	ʈg�h��x4�n� ;z�ũu¬c�:�5����6�GQ�<4G�uj=6����6A��iy؛�|k�d�Bl�8�i��(0i./+u��dXP�.bQhԿ�uǃ�&�@ɺ��~]c\bf	F j�."�������qg�=! 7O�����w;P�&�I�7y�lYHE:�$]�V鶁P�z�s�z�~��ɖ��ޞ{'Ӝ|T�&�z�B/;��`�!��F�t�[-\��NHC��S-m�m�66�?����}6�I���:��N��y<0������D�&���fY��G�fQ�~L�:U���K����]�ّ��9MG�<�>^���t`[1 ��:�dP,����y =k�x|Z���:�:�z��u���~>��
ay9��?��nn��:QçUK}��s����dd��@�c'@s�up�M@�g^�ߠ8=ԍ��Ď9��_i���4E��`Rv��j��L�w��4�g*��$Љu�Q#�S�׫Yw?0�Є�I�ګ��%����"���_���4����)c�T�f٪EZ���s�.hacЧY�մ:��|ik�1�/@^��-P�o޾h!'wZ&��|�E�Pn��i�m�g�M8;��(o<nk࠵_^NrZ4{v$-�RN�"�ح�������;Xǔ�"7އ�zUէ�������d��: ��4mD�T��^vAzp�SR�B�T�GB�W_4:L�qP�e����FX�=Z-�(;(̦#�6��9R��y	P�Q�#k�!�:Ic#�i�F ��R6��Y!�Ս��"�jk�Ƙ6Ko ��beh	���}�̬02]P4��d"�H�׺'�h�x>��&=+Ϭm.�1 KӋ��q�n�{8���m��l�L&u�3)�dMɡ9�/��ڱ~_���iD�kGL��TAZ:V#�ut��=#H�����3,_�h��)��Lܷ�[�JX�����I0�V�mm�� Y3Y�Z�4_C6�b 1��kV������m:j��'y�/c! ��z�~��ɶ��I�<M;ת���rx� �R괪=*�b���Q},��Q]<���m�K��6���ky�q�����X>czj�)���)����<�X4�vx=j�����6Ӊ����" B�h�k�E���0��
�$F2��}ȿ�5J��iJN�\6�I |��#��~����Y�S@��]<�\�)�`�hk+���GX
�5Ӱ�rZ�m�l[�,
����@��FlT����ڨp�!��m�͈ۤ���Tuj�wW��šwʷdش�r�Ҵ�bc����6tc/��KN�\��Mr���>����g=
��F�u]耺nT�ox��s3â��6"m3ښ�ծmʠlj�e�(�}������^uC�e������1Ԯ����H�q�勂��mp��}�/�S�%0뚇X��x�L��NziPv@zp�#ҭc�?�-���2B
��!S<a�A�N^�[��AR\�.��&�?�Yi �iI�k������1<���[II�5�Z|�`�Il
��Q��Ŧ(j�^Kz<�6檫t(P� ���:]��P�O�5����z^y<1}�;�E�?:ٺz.VG�4ϮHN�\���y2ok;@�|��uRu:P^���S����.�lK��jXL�(�Qv1v���~P8h�0�}�2}`�֦�a��,P�uJ�@�T�8,���l=O{;���\jrY�m�ዲ��<��e.�1��K���hqt����ʗa�z�ӗ�l����;	����b����gK�4�Q��ʀ����Q�(�ꄻ�ɦh��|�t�~�Y�M~C��U�¶�:k�����Z����O���Kc�������<-��sZ^�xb���qc����
<�?�޳�u\�< �\���<S]=������ϳ��TW=��0rt�c 	� �q3���ZȌ+��H�l�cccׅϿ�;,+�?C�k����Q=�����_�?n���W���ɔ�pf�Io��p57�åC�&EC�g��mp�D1��1.���$8��ﺳc��(�g�`ſ�M�1���(�8���c���^��1�?2�x_l-��-v��X��q	��J�ćV���C�;vm��������1c��ba�s���x����CQ\���q��3���]w��?s��!���~$�{�OM�����כ��䕧͆_TC����"n?[�ѮSV��퐶��L(��������1��*�� :����6�V�� 8����{��	댁��TJ����B�������V�c �G~�HM���!��a�����L=��x*��P[�>��狒c}�X��5}{���ן�'��ͅ����x\�e� ��/��>ʚLa�ӷ�C8���@2�e��,�8�*3l�X�cB�%�˓ʗx/�S@�r�6:/������JS�}؏��Ru��B�>��WCu�熼�|p���]�)��_2<�w"u�c�p�i�yz]�?~���W���v�g/������ ���cz=:1�dZ�py�{j��
��J���4c��S!�SmW�1V"&R�f��X�R��kC���{=�g���K�KX�T�p�b�c?R�bؗ���4�������@����~OMC�\���<��Vk�kz}�
N. �,3pL cs�:Nf}����
��Y�I���>)���Votlx7�C+Թ�$5yF��9�ƀ��Z�-N����1&f�?���#&�؆��	�O��)A��4TFL���x)���^�S�L
DN���!V"V��J<Me�R���O��,6 ʜ�o��h������ �MHL�'/;���f����a30)�Ij�������d�7�}bNW��W�>Q�C�fX�TЄ��!�;Ĉ�)~c������^��%���Oa������&k��1g�<�-������� 6���~]b/!]��$��&D廍w�{���O ު}B�b����K�B:k����ϸ׎,t��kS�c��[M�s>8�����8u�=&�b@-և��4��jS꾆���[h^�-`˕zԌ�?/�c(��2���xNիX�s����������J�u��>Ca�@i��a! ��Z=�<=hQ��SJ,�&���&�I�w���t\��ϥ��gJYc��d9����p�R�:����/��3�I��X�0��v�ߓ)�^ŀ�oi��2|�0�@o�!Lbn�a
=��������է�ّSPB��#����N��πqa����CAǽm��6A�~:N"1`rL�1.Z��g����PW� ������ UH����k튬N�<���-��n���,aߦ��z��_��pe�p������c}n��c9b "Uo�����9hR�����~�S����s��]s�>�W�w&�����ҙq�=O�`'-��XA��'񗒿^XB"�M,���_��G�CH���-�V[�%1��$O�=��y0�=_�懧mR��e�n��U��/�?*ol��
���4Auʘ�p<���`�VB8����.�L�V[eǄ��G ��J�'T�@�?�1&�Wu�yS�#<~�v}֖Tݱ����1�\2莍E�R���ߩ�6Ų��0����?x�]�ܱ<W���^U���W��˥Q���;9� 6�2�	ЏJ9|�WF�=9&b)%�^�b�"ݏ�6�՛r����<zRlGJ}䷡"��ߧN�ߚ~��SJ���b
b�"��]C�S�%V��)�뾇jחX��0�@�t��������5�Z��zǆ��� �+(��t'�<=?B/�]̀?�Ћ�V� >h	Wk)���5���*q*H�'���!�'���������9�X �>�M�߯��?c�1֦������-VFا����1a�p<�س������;�,Ǟ�#`;/w�E�2�c�.�M�gJ��s����p���佪v.!]��+O��ۑ8n4�Nt���/]5�J��TZ���&% S��%B|*e�Z��Է��0�������?xU�M,��b��Bn��M�{��b���!�WN�(���,�@oXoȜ���16$�֩c�v����M
\]���t�
N. �L�*ƜH
W���pl�	��)�_a��T��6���uN)P�����$a_��@,�wؿ����j�!��ǔ��	�)��O=�S@Y����KD���ڞ9C������[��)�#�R����k��t'�?��{&�8Q*NI�y���TV%�;6�l\���%P,��A7�&�1�����߱�;�F�ׁ�o.c)N�^�J��ύ]?f� ũ��ػT9~ܛ���_l�ð�1�bX�ާ���?���иLI��f����س?v�{	�
N^yzzq��^�����䏽�C��<WVz����
�1&'u|lB�|��Q²Rm��~ j� j�V���є:~kC�8����6/􏍍��$�c�S��%`��S��T�j��j� �T=�5�E�+8���aL�V�����㗮��F<�/H�&�)y�(�)�$�M]}��O���X<R�ı�S��X�*#Rm����'�7Vo�ekV��)P2%�kÔ����cS�5e�8�6��v��~�S��@���@<���W[����W�䕧+8y����_N�c���>ڟϝNJ)�dH �&��
/�7��p���U��O�XǮ��KXf,��ߗ������ɿ>nޫ5z�i~��c��
�X;�z���z�&%���-�����/nC� ��g6�����_(Ln���C)u_���?�.G���ד���'R��T��;x���'A����ucǸ6u�;OM���'� r��cSV�����(�yi�N���4��1֦� </����,���	͡�l�}SA㷤ic3�Ƙ�X���Ş��ک�Y�X���ϖ��s,��wWOj�򒶅������S{�p9�������D�	��!v�e�ٓp2r'[}���/ć���Oƾď.�ʊ�q��`��E�ϡ��
2��B`5u<b��/�������S��H^9/mH����ȇ�8�M���5�6��6�7VS��뇀Zl���!�b*(�������������S�D���R������&�)PzU��RL������6DǀAj� �phM%a�C�Oa��cB�̐{Ưs��]=�1;��c��D�i�MSAܔ�a<�|KC�(����/ʇ�chB`���ީqq��f�&�sV|!Ee��t�5�oIWp���-��z�Ձ�=���dv:���uC��|���5VNxM��T6�Ō�b"�kR�OBb���>E�Ǯ�:V^�o�LY���9$N뛲�N�'��LM�ߺ��=gC�w�)	�7��X�-��bj������}���!�n蹉-fR�F���m�T��2~Ә�kz��
N^2���a'�ɽ�N=��1�b
'���!��~+C��b���cn�M�-�Q��"�c���b����r��~;S�B�S 3�mߒbs���0MC a(��J�}b�Rl���g;���0F��~���3v�b����;���OWp����0�B=� {��y����+#Vg�N�����X~�'����Qj���I�ql<�R��9v��v���O*f�@���T�~Kz)`cSR}�ˍ�),M�}S��R�'ņ���c -�g�5J���8�ꚲ�	���.��x�r��\B����@�L6Cl�i�qF dfb+Ⱍ�<��R���5!�����7�|1$�B�1�	��X����C*����9�����T�~k:t��\^?p��_��?���á�S�W�!�H)�<v�[�E����ݧ0\�@I���B�KHWpr	_�3o�#�P�?��'B��i@��*;!��bR��!�����\Y�'R��a��/bC�#dR���) .
R$��� pFA�l~[��?�Kʅ&ug�A�h�l}=��y���z,�(��qm|,�[<I�V	�8�Ւ�ͧ"��#��a�c4V5���쾧�lb`'��Ąk��Ǟ�cw� |��Lh~�����QXw��X_�����ɘ�A�e�+8y�	�b�3��PT,x�V��d��Y��'-��� �d"��w�^�_=/;��J.�(�<��������NV��݅�|C!%�cyS)��S� U��2 �U(;ĥ��6�eW��޻N�C��'3Vo!���Aam�����r\C�0��L������&mu�1� 
1u����R�䱠��������_C"���� t>��a��y渭R?���c���G�J���l0.�uӁ�4�ڎ�<�j���C�\*���'B�2a�ήj�-	�i�\�'�wLU5�~�X�X]~}�N�X����gpM�?]��$������+��D	�����&���l"°W����y�영_���SαX�>L���RЩ���W�C��d5Lv=�*	tp�V�20a �&-�@���m����w x0���k��{A��\�+L,X��Ҁc_,V��>Es�Zc���d(������8g�ßt��3��B��p�^��+�X��{?v}�js
,��}؞��!��o��j_���@|�]�������.�����+8��D�Df�jl��:P�:b�[�Bb����w8q�&E����M��U�����G,\ Z�#5�Z�L�KRC�1������/z�[�U�h�^uV�g�@�<8�Ʃ��}�;��eX�
��2X8�F ]H5v��6�N�PFJѠ �dX��^��,�2E}4�*��a�U���1]�NEXdc����i�e�?���س0�،��0_�NǎO}V�@�P?�k�`"=��S�i����ל����'�3_��LY����/+F���c���;�W�K&�Tz�0'�]�h#-�k��bN& ������0VD�Y�B_��:���O��% �9/,��B�, ̑hV�X6B	'B�J�m��ҫ#8B�c9���@�G@�1�hY��{QU	�@�9P?���gUT&�'Ӊ�I�j-sc@�N�^R�dp�`����� ���^;Ģ�T��������R,��J[bc"��{}M�3]��$e��&���,F�&��xl9�,��~N��m��؄�=Ī�jlRL�=��T�T�&Y�S��X�o?Y�қ��ЩP\~����_b	��h�m���X��
4P���-h�Vd}� ��Gw����,���Xے3CUz˜X��U/�`Ǣ����!fp�]! �c�G�f��w��b��L'�7����P��Z��	<��c ��ȓz&RL^���wȕ��o��j�_G8��)�Kk�_v���9~|�YERw��
��\@BX2io�5��ԩ���b8��؅��ܩ:��c `
]?�RL�?ɿd���8P�]�l-������a�hV����cH�OlD��Ϭ:�E����k�S�t��>p@���X��$�kP�7���#*s�P"���D��0�;�1��0��I�}fہ��ڶ�=��>g���V��ic�1|N�=w�����9�����X��5�w"��uǞC���z$��bO��#�c��/f���uO�a��t'�s�ߏ�"�ѭv�mp�c/jB'�0����'�{[��Vo�gx>�R`&l��pׄ������Lp�D;��Um�f�.*e�C/�٘VYf
��k�B�#c[g���ň-�1����،���o�2;\�����#O"vGx�Lc�9O�x!H"u;Y;���;�]l	���SF}ҝ�P�2�:r�3E]�v1�~�?D6u�ТӁ���c���?�:������.�!���!,�� ������[S���;+3���!&3LW���HWp��.��1���6N}�L�U��;��%�?��OV�^�c�E�	��)H�>������rb}��?i�A�˭t:�� ��v�IH�^1$un�=�0�]4��.�kkl*��%�G�eŶ��9�d�"]{��]Z�M���$G6��4z�uQVd4�X��6 =���AS޻碑�X����:�`�p3%}T=�ɱ�9���6˱HbN(�?%f׭�-��v0߉���Ci�t��w�
C�'v<|&�p��x-�E@���-F��C�-�3,7�h	�@�'���Օ���\D�_�i�1�Ҿ��LM@~yc ���������S�{�R�������	���\u�ǜ,�?Y����Cp�Q��)a[�ΰJ�!�;F�S,�7Z�E�^bRH�B@��F����S,�!|FǞ4΃�� lđE�>���c;������M=�Ŷ1���8��D����AK��,el��Y͏ �h?�Bg�;��ݜ��)ihƞu�>	Y� ����c<c�����$�Y=��)�o��}��os�bf�9"P�Z8Į�z�����+8��������V�	���;��U�T�{�::L@�E�]�K~9D{�H��2��`�����������S���c�߷X�) ��pL�@F��LM�Q t`� 7�UX:#( F��L�6M�eER�\��ȗs�6� �}�iؔ�%!�e�Y�~/��p}:�3Qc}-֑c����Z̟g�v��е-0�N�v��`n+�1X(��:�*R�mOB��^���UΠ��K�U�p�M;߇��cm������}��'�`�� Ya����}�E	����3�gŝ���P^߭������Ǟ��mO@}ϼ����EC�/��3�?�cm�G�|����ϙ���ҹ�t'��2~1-@9���+0t�R8�9CV���-��N	ߓ��\�RWH�&���\�H8|��+֎��K�u:泟�FNN�w�r��Dc�$�K�8V��:	�n�eBZr&C�\G�ۥ�[6C-3tt]���p��#=ή�H�}�B�k�+�`C�q4�U�贽*� �P.��?�I����u.���Y3� i�jKn�5	��0Ω�å�*t�A�%R�x�t�f��O%�N�I��4�*�Ҙ������;�~��J��!��۬���zGb�}I�]�mZb�f��WWXr1�
N. ��j��Dh�!����j+��=Fzo��X��J�6�W�\�;��%����s)
9&����5�$�������&�_캳IX���a��V���J�X�+e��P��Lu|o����lAg(*�Fd�$�I�7=�H�l��X�B�*؆B�@��rlC�]CV`r�(9��	Ǩ����Ta��a��e�o�mf��� �:�L�V��W��&�**��F�D�Y����ܐM�W�	����\��Y��%������geH�ʞR���!05��捡�SX'��H����������է+8y����`���UIlR;_Iy�㴂X9��0�1g�I��~ݡ�=��AL���P�c���ت6Pb�'��2�ٕ�&�q��IǑIJ��~˶&��!�Ь�\��3#�B������� �
���C�
+;l_�n�����փF ����1�F��;.�X�\a؀�V
%���>�Zh��[��w1>d������]�^��"#��L;̿�:͌w��h+��ض1pӆ�v[�/c��+e=�"�7&Ƙ��4��f���������}�
���BaYC��e����f]��IWpr�jb�o��UT(�c2�O��PS�Ɣ�7f���8��!�|h�KM�c��A����~�zt�l(jD���l&j7y�l`Y�-�w=��|�U(��-o�U3'y� �X���1�f��L`˾Q��K�4%�)\|� ��r�E��a�q`���<��m;�\�������w޶p�'��}_�^��K�UlB^=��{l��EK�"�؋=
�����4^;�� �&�5�=�l����2��N�)p�*� t
܎��}x�j�[�K�	��Եc�٘'�����/CL�X~�m!�J���V��Z��\@RYnt��>Qe�\�	qw,tM�<b�2R�x	U��v�B)��}x]��H���Jl�Q9�Q*���*,�[f���P�k������73�,�EF �f�L����f�� �D�]�w�����aV�w+e�U(������k���-aGl�� ��E��z�Pb���F�Δl��\u���R�X2^U-��g�~����a��P��d��^�Ī�d}�v�- n��Y ��	���f�u��-�_���]�lu�\(�4��X��˦�MږfDb����gbL]�{��%R��X��L� ��P����\��.#]��$�:�j��݆;�[��&ǡ��V/���Vu��a*ʤS�*�)+�P5��23c�O�e,۝�~�!̎L�b���Y`p�S�P�"0�~�ê@�{��43x��p_b�[��
�:����@`2����V%0[���PTUo��@���O0(�k�ˬ��g�x�����Ĳkʩ��U����+5��#x����b���6+|��ʰ�*�`��T���ia%�
�;�-z��la6�3�4�̰g1f%��%�FF�?29�sc�g!����)�>vM
�O)o�9&a��:�����cmw���l~�Sr�����\B��Y����v
L���\
�&��m�ņj�C9���44a��𯋩��`��u�{��e3�� �(��S+�T_��y�-����iaM�_��!��Pܒf���Y��n�{��mg@2����� ���w6{hLE����
?.JX"H���|����ao<T����U뺃_�5�|&��"V����r2 �q9*PG�n�B����w9�a������n1O�Q]�������o� ���y�����~�B���v�`A��lK���Ӊ������Ub�ۛ�Pwߧ���3�b�r~�~�]*wj��+)P�:c �^o���H#Ԇ�� ?�x$�S��&0��?e7$~����KI��Ю@�|�p��M���L��52~�C�����CUX�b����~3r�r[E�g6ș�a�
&=
s��:�:��3�����#���`�� ��n�������j� ٚ �X��n����^�>�+��`��l�5���0pSdP! i��I߬ڜ�亳�
J�Zgs ���F8�U���f���`�S��אi>-���w�+���A�L���<�g�Z=���a�����s��,�����I�����z��ؾ�E�5 �f�㪾0OL��D%�!{{'^��cF�s/Qg1+1�eL����5�����vi�:�^���HF���D�9p��ϋ0)�`����?G!@��N6��{	}Ϫo�	#NBp>5y�"����Ȑ�7sj��O�ǉ�P�	Xq�h}��K������!�?"�~�3:6(�	�qם�(��tㆍ]��(�[%ߕ�͂����묖��p�}�^�S�}��®+ �K��½����5��TP$X����k�#��5^�X�B�y��T*~N����}�+e����V�)�����m=Z�C�ɝ�l�di��N�j5�_�P??A����f���Яؑۻ𳚑7��I+�������fv�ۿp4؆7Sα��>`C�������O�R��c�X�N�F<6���T���^�b�~�˚�.
��{
x�������Z�w5T���b��c�C�n�ůϕ��$��k���HWpr1��ԭ��� F�nR0'�3
�p"�� ��*�����KT ��!:}�ݩv�ׅ)%h~KZ���!���CK���F\a���,S�
𒣰P�%Ty_6P��k�.�sk`����C����7x�gC�˨�/�A�+'^ǱD�*���O�F���F�K=oh��f/	�V`=���ENDO��5��
ʪ�|�������QH|*��y�ނ�gP�ʜ�F�~�y�����oa;ۼ��	���6i�I���*GOQf꽚�/�������R�¡���O�)֮�!����������-ꘫ*������D��W�8;�	�4�dMM"cz�p��;W���s� ��=59���y�y�ޡ�N�M��v�������r1cҳ���kt��v�Z�p�׮�cd���U����(���]K�?�����z�"���hm�a�IR�������=th>��ȃ&�a�i2S���&�$�)<����7nwam!�S�0�ru�
�l7�ݒ�-�-n���@��� )P�XT�.�s-Qb�{.���W�v��j>�;�i`�u8&4Yƀ�S���z뀴���WmeM`3���=��3�����1�����$տ	�֛b��K����O*���y@܉�^}���HZ����4b��vB�$�J����g����$v>UNxN&�ӽB�5����|r<�36�%c��XN@�`��.)$Ĳ#�>WY	]�q^�j?�����q9���+X�|���u�3��%����Z��uzC6$4$��I�t�۹�>���0��&&�a�310�y���$k!�'�!5Ԣ]��L��Ӯ����9j�
����
���h�/'kkX"�xK6#��SC������_�i��箄���9�3F\��ظ)����1JB�k�?)&�[���,FJ8���#Uw��PM�bx� ������@���}N�7��k^O��W�]��MWprI���C����l��ac+���^>Ӫ��LJ�=4�W��^EX�6��p8�f5c|�㦅a{�Pֱ���x�c]a��C�����R��K�Š�1�"����i��6/�ݪ�w�����_��j���j� �P`5���e����iizȻ��XJ@�6�;
�^��D���)qm�"DDv(d'�+1ⅺ��E��ṭ`�n�Ɔ�a��/4|�<�v:_��M�溇�9��OS�]�8C�������vz�{��Xʶ���d�"JY&ȴª	�r'ST/}���X�c�y�:4v,Ŕ��J\��s�Lߖ,����hY���;��ʞ��t'�D�s'>["��~ˇ�!�p����$*�X�?���~��z+O�,s�ђ���������Ҕ���ɇu��m
cB�D���З�fb����0�ĳ�%V�w��y߀�����-�W
�/s����(��f�u_�!	� �7U�㈪$��
����
lTê��X�gd��"�mFhd��c6�6�S}�Pb7�
:)�V�>��aY4x;���<�COƷ%	��i����`��@v9[pY�����6�S��'���A4%�E�q�1��7MsbHL��.t�N�
�P���C <LS���b>�XΐII�d��5���1�c�O��n��%�����'�;(�k�{V>�1�����<�gJ��bT��n>F��b��S�Lj���@���
GA�Ƣ�Lf�2"6T6P�
~E��ض쮻|������MYæ[�������|P�2t%o%�A�Ҭ
�!�rh��_E3�  ЪAy I���[�`�{XuO�}��wx|����r)~���eض��#!V'#�$�=�m����v���J[X���K̷��
1 ��A4L26E�m@���ݻ�C�a�]�=W1��oz&^�z��lF��>P�������+ec*�1ur|T4�c��2��\@��J�m�m�m�,{ �.��D���W~��	?�,J�p)h�v�m�ُM�a��=�j-զ�
05�����\#�V�Hݤ�U�ҽϘ��P��@g��氇�y_w���� �j��w��:�mwx�rע�M��ۡp�?C�J6� kưMH�ZK95\����g����J��	m�������ި�+̹¶�J(��2�P5����,�f7喀���_�|�n`S�x��������� ��È���ƶ0�����cR��x�%�����oM)���R�[���]�L111�PX��X����)`���ė����R�`j�:@!��	�� ��&�G���ء�>4������z��,N��N�:L��I1B�+T�ۯk����#�$�,�d���C�K4V��%4�RX�{�{�Qp��=�x&_�`�_ç��󭆊⤴X~��+��4^%��{!-�3F�!�������+`݋Ie�[�V�@�!D@��rȲ�j�b��ϔ2�Ţ7����;��s�Yi�
v��6Qû����c����챎,�C 5��&?����A-F��d<���$��SY�1uD�Uq�_¬� ��4��IՕb�ʋ��Cm��ͩ�fx���ʜ\J���HYV�(���0��AY=��\t"��cB�I�gE�؈�+��zȟ�&���Y);��4�6:?~��sU�t�a�vvz���hρ�2Q�@kU6XVہn��~���W��������������PP�T�I���y�Lv5
�=���p)�Z�1;	`fZf@2/�l���'�VQl�ҏ����l�j� �
�¶)PA63�u�����WlG��p���]�����y�]������l�@�7@� b���G�/���@�����^6 G!�k�'�Q ��IƱ\������\��g��1)�1�F#|�c�~�����C &|�S�dJ�b�I1�������t�R�\�%�+8��d���gy�����5 $��J'&l�=kb���R��]�!���6���ُ�	6�C,�/�Rm�����{V�XSQ��v�?
����З8V���ֿ@�%��/O�7���n����%�����e�;/�j�Y,m�W7����?�,�l��&k� �Y	������װ��š���g��o��6tD�d��2����"�Z��K��\��^@��u���~9��s�[�7o �7%Bh�˛C����_j�K�*���L����C��Ф�h�4L��h#��z��Oj��]�3���UL�ǘ�10U��Ac���|��iJ���R�I��t���[@8u��6�r�Փ�2��\@�޿aJM�!;1e���e�u��5F�����2���ZF8�5/nu24�A�! ���]~Y��6�)W��}l
lr�}�v�y������;X}y�O���[��_���j�B����>7�J"���5��w9�y��կ�����x����|� ��%��
t�8���fp���=�^?�ҏЗ��B��>!�ٗ����<4%|Vw�5����;�='��#������
�~� �X�A��N�=�FC����{����������eW�Ocަ�I��.��ʼ�f�bR&=�SX��L�c �]?v<,;|����)it�dbc�����&�q���<G�� ]����a��<�I6�t�-�NcP����S�n���3��h���15��?�<��xW��A�/���! ��R�z�FW�
����s-�����Vw�m�Dr���u}��/4��AM����\�/�����ÿ�S�87�k�ty�j��=|�+h�4�dF�Q����#�QEζ�(+Xc=��	�r��~�|���6�[��7�"��e�-|�[X��:(�.Z`Y3��+A!P�8�6\��n��a� ���{N�t�L��<�����	�ѹ���jć����w(���~�Ҕ@���r�4�Le��2c��Qucٓx����������d���bM���I5U�� �t��S��X,��1O��c��Z*&�����X�S�Pb��1�P6"kρ���+�gN�g��Lq���i��`���Kȱ���z��m��f�����v����'��}���*^|����F����1[A]b=����ll��|��)�ZR/5<�dv���&�ws�c���vP�0o`��ܛ��챍_��[�s����p r���p@�M�C��^J�/�c�����l���!vņ�'�
._�H'�Z�)ޘP�s�nB76�ܳ�u��0	�ߢ�q����4�����}��ީ�����.f���x����(����HWpr!�F�u���w;mhꎅ���$�f!��u�8�ѩr����ECL��ﴝ�	�% %d]B�:U��ɛ�	V�C�z�Ȱ���¯���9Ժ�/���⩁��a��w'�fs�UĲ쩣[jK���P��|�kXu[��g�����ht�K6>�e
��bŠ�,�?JZV�pP{�G���²+�a{9�,�{Ԍ��r;�p�[5g��iQ a;���s�5�_�y�֪l:Vm�̾��ho@����l���8m�����k����R�{{c�F�kcSyc�cJ��_?��sEXƷ��;��MK�=<�����ך����k���:� ��'��R�1�oXF(�S{�
,�?
���ih2�㤼��$�e��9S��q�D	 �����l��Y#ٞ�]
�sB���T:E�?
>϶-Y���@��{���&�6�刭��Bp3�xQ���_ɶ��I;(���V! ��*�\��=h�����DF����X�BS;���q;#�g�
A �S\�gU1,Z�����D}DDR`���!�9]O�&���&<�氏��:��S�`���X�!0�'̸�����PJ�`���-���%�f,�Ђ �/Dn�+	�n���H��]��عI����>K��pB}Z�/��� Ą����!K?�#�P�j+��ˌ��EƉz��K����<YK�/�W�x ������z��*�j^��q��X0��1�m�k�����1r܀.�ŴQ_�@Uh���Q`����(2H�C��u�����Tx�@��3	�����3�c[�@�|��BY�G���*��ZD"]��2ـ��E�"�f�wR�ꆮ�(�=g`;O���R~���Mj�xEٌ�*C����A�E@�⭐{0=���(���G�u�p�+��㛡�ss����>?�>�GV�83G"��P��!�����_���rw�Nؽ�\^����|Xp�Z8R?.�qG�TJ�_�4��~	bT}��B��(ls�^Ю���+8������>�;�T�B��ꏺ]:&�TY��+�H�ä�!w�(�#���
jL�&�Š6j�JD�v�$L+p]�m��de�j�@g�0�����9π@I>�oF�Z��Kms%ڂ'L��'�#�ᨰv�",��m���v���QZy^����}�����\�J�X*��]��=5cw[�����P�-"U��~�2'ٸPs���lPy�0�%{���~����1m�Ɔ���¹P�b���qw���}���L���&�eg$2�3�]�P�}dP�5��}��Bc��	���&�籗������K�Q�F�Ʃ�<�D�(�G��:�Pv?�^T���-���[F[��-l����7�[���<1U�Kc���o����1��:^/y��+b��t'�N1镏L�ʾ�8-�v�5N�֜�4g��y}2��N��N��+���>�����ʒ�c8�e%:�%mse��x64�	�W^�,t,��s���#��l�t%������-��^ #+u�;tC�p%K��3b�J���=td���u"�is���_{ ���O�nA��E�����9Bk�O�[�[P�
#�������w?6�~���<�Į���1�V�p�.�*H�N�8J,���m|[����F��})�=����z �!02%b��O*�ke���=
�N�6/��xw�2��P�&X�r��'\-��A\e��c!}U^˺��4*['�5Ȏ���h��,q{Ʋ)���������,���P��t�ٵ+���c�TOC)T� ��#SGˈ/Z虶����^]���H<���	���A@����}w奘58ɝ��y��-t��#�]q%���P�)h>�9	��9���,�e���b�������ue�Q�Z�M�l�q�)�]�V���k3�jb8:f8n���t��M�:F9����A6��fJ�h�V}Fk+�r�>t����U����j)ˤq߱`��`��!�Q��C�w"<܆{�}O6"$8h���,�d�+�#;�8��Z�݈ip�H|�!�V�K����6?��BI�}��F�U�(�ƎOd'C�ǚX#�$j�\��#�ުt8���2ym���/R�u�dLh	e0�`V$����m�س-��,SfPgyr[ۆ���#��1d�b"^�>�cc�����0QV/-W�s6rn�����י��������&�r�L&�98@e�Z?�����2Ɍ�)N���Ή1!s vU�	7b�� �	nŬ	UZ�f}N}㢲��,�Eo��:3fU���~Àݛ�6���X�l?a�9�䭪� "z�Ml �2�Sv��e�����n�Y����I-L���ҡqQZ���>3��`�7��6((�=�_y߈{17̀�8!#�Έ��H%D�I����E�7���]E�r���U�)��!�M�����$� ��-�C�kt�d��Q� ����:��P?��Z����`@�i+�%դQ��ʳVD�.f�P;��^��?w��G&�4�V�vԄ��=�T';43���^򦄝 Yz&(�.���h3F�<сJ-{ �jH	�&ne[�[tL ���n���^2'�c�1`���}c��\���t'�?�ڱw,�`���n�ᘓ@���<!e<mb����J,v�l%���{^�*��6}/6!�PV�10�Z����p�No�K�5�dA��Go��+$�H���zh�(� �Ԯ��0Ul#&1vR��V��K�2N=	|l7y��:� J�Y wlbw{dЕ[6L�T �-H���[�ǈ|rc��/�����[��a�,j
�"�̜H9b�����D'��[v�V�LR�ʩ��ș��콣� V���nMy��E<�_�I�b���BZ�J���+mXH��⪐��lkD�/�x�����U@t�Ŗ�$��`%����f��w��->�8�Z��tV��CA�<��s:�����P�sA��(�26�~�`le�'��=���c,�bfl�9b���@+�`w�]�����r*_J��^;���v�+uu�t'���у�e��{� s:u����^���b����)g�T9���MV����Mab�����4�7B�I)��"F���4�z ���Ac��ʖ�ʕ�if}Ͷ+�)rِN[�(������Z���
ޝ��H�d�U���p٬��ּ;/�Q�j%��- #cUIm�&fJ �ty�L	�v̰��!��ӱ���P@����[N�?bhHյ2�
zS ��P�S_kf/�_�ܕAư�kh��x�7TL@�{Xݦ \�<�1 ۙ�UG�+30{A�Y"���̒1�b '�*��`�!#�^�z�� ˒�۵l"�c�Jb3��H�j��s�������P�����M � ��qK(��=��V�(�ozH��sA M�e�`&F˽gC�N�C+����A�_R���I^RWʣ'/���z�X�2��\@��T�������h��^�,IJG���N'�t�%_�ꓱ�r�p:-���ŕ]q6�Ӯ�_��!��B���5��z0�����h�� ��v%"p�Z�Կ��Ƴ�ы�B!�ql�|	 ����0�]lZ:R9u;�O+f�ְ��~1�`A�Y��g�H�j������AأKkA�.����ݳ͉�)�5Vs�Y��v@�Z$��#	[M�TO�X/��3��U�F)�J��ql+�e%��!S\bT�F�W�e(�=�C�`O��aF�+r�c��O!�S�c`�)0����"���n'�Ye��|8�����f�AC��81e�9
-P����C�2��v����}�E��}��'�o���m�g��X3��a.���WavP�;f|�b��k�{�3���A?t�{}dI�>I�Eg�4�^��C�#/�7���9@I�-�i"���M�u翋HWpr������XO	��x��ɧO�Zc����lb�dH���EP����vǂ;g�������`T��AEwodg_���	c��N��F�X�����۲�Kf�w}��`���ٝ���YS�_I���*TÌĎx-N�ܓf����B���ס6�g�iN+�2�%����wx��a�Ӣ����&� k��]�Iu԰-K�oŦFK;�N�����G˷�gpW�5T-��iG`l;f��W�X"H!����x�i���U����a��l��ki�A3�i>Ò����֪L�lL��l X���lce�l���B`��6��(`�LK���;��W�	�8~�gUޓ�\Cgmfp�����0�}�d�\�f���ľ�
�o����ZM-�(V����K�ߗ[�
�gf˪%bl���-��5��l�sx���Z�#��������/_p��{b��ާ�ky.��d� >_��������5�B7�1P����v���1������\@�FO�89$�0��1' e�͘tU�'Fݺ��Fx���v^�S�U�xf� Jc��a5F٭a�o�% ����Y�~ƻ�JV�9
2e�"ߕX��Q�� �kӘ~q0���pN�b�-�C��ݮ�n2\ɳ犸�R�=J�',gK��Q�R�$X�X�Q�l�C�a�P���s�(<�,H(|�`�KV9 �V�����ƶ����-���KN`��uz7Uz^�����$1�ٰ�f�q�_�W �j����_���e�k�5��U^����M��GD+��CPQ�-
e��y���]��~|����w`z~fP�K������rv{��|�*�M�BLI*�s4��;������lH��d|���~�m�r-[�/�=��p��d�,3��)q��{�2�ϦB��1�E v�}3׼a���<Y�ٱ�T�`����� �|W" #����x�����~�g�ü������A޵��(�Q��M?�����_�3aXh�ͬ�	ǂ�r<n�z'��.�.|�b��a~���j(Pd���)k7v�9��̕9��t'��U0ù��)xP�EQ=�=�28-+��{�V�'��Wl'Fl�	o����c翃�+�"��$©a`r��
�U5�/*(q՛�r\I������4��^�h�
���A ���=���LVo��Rd�=��	P@�٨�<]����un���l��e�L\��a��jᏳ�C��Y��]�!���O��u��;\Q�a�C P�]&������˗��ݳ�-�c����wbj���kQq8{�U�Qb��n����
�e�=��n�`#��zͣ7�����7
��f溁���Js�ؾF������B`����>�ҷ��o��=��[��v��X� {�g��MY��2�����m�_7�ך ��)�i�M�})�<���-����=J�5�1/�nlplߔ���Χ��$c������eힾ"�����gx�*��5��y�["�+�2<#~%֩��0��#&����3c_>�ؐ�﵀Lf��|K�WsD���<�J��8��I����f�J�GE���_>�������7w��}�`��?+b�J�Rbއ�آ�U�ή(0�X�!C�����6l�|�6�u��%ʳ7�:=�<d��P�������$�G\���yy]��y����O\�ˆW\�UYN�y��q�t��{'ٔ8�s'��0L�`a3�o��XuL��3}����A�B������2$o�-�i��#
��Ơ@!.���	�D�26(jbGȖӲy�r	�Z\�7O`�9��������7��
�
���U����w4�<�u+l���8o@�5|�6��4^�Z-�Ow(��m�Ɲwطw�Ԣp}ء0��,b;\�?�ξ��?��U9;����|����3l�eO(ܣ�|��!x���z�c�� ��M���
f^b��o��nN6$���]�c�����~��q�>���,��z��"�}#�v>~��
��]�����ݧ}��Mś.�=A���_qLz�Ws������w�%`c`���eP�*�g8������0����wo�p��櫒�-l��$��`Bm��E�6S� "��,h��L������G4G�}z�v�5o��d�*L1O4�F!�j�G�0�v��ם���j3�����5,D���:i|֖���X��q]�݃�m��Vc��x��P���L����3��/�v3p
vܜb����W���������}�� Ϣ_J�:�S�?8�jC��~R��2�&e�	(Om\p}s`P89~[�gP�jt�o���-
w\㉻���?|�r���Z��1�5,�}s{��٣d�K��҈Qmo���5�V$ �(k�){�ob7���B��7���	��mE�P��p��u� է-���?W������Ea��B0������*QHJ4���&UO���blrأ����&C���P#`�B싈�����輻]��̯����nɂ�q��2����B��F�G���}�����{����P`9o�V�v�e�����
�U-�?�����kZ��3ؑZm����,��OF���M���D�Q"fB���,��x�"�X�����#�Ap��d� <#�zFp���Q�#`�~��-�P�Kq^jBc�c���a(��;�ν��h#n�Ěqt^~F�&�`C��$��9��ރ�����{y�v"�����+�q,{����<�6���Ut��{��e�H�( �g�ݭڗ�c�6�sS�ϰ���S���v*�P��Ȯ��L���潦W����Np�ݦp�8Q����c��%���߮����ۺ���P5F�u�'�_J�Γ�#+(�QP�{�[M�X��ZCen�7���K��`[��p�bDۉKko��J���2G��=�Pl�f��_t(�co������ѣ��f.����=��5w��@����y�l'��f�����УP/�
�x�!3��c�$,�����(�tž%$�zR����%Ǡ��d�+
��;7��`��� �æ7��nsV	��#ے��y���`���%F@����޳��j�X�|����AÞ�Ps���+n�{�G��m���}>�mYº��6#ۚf�bY�!��%�8�y�p�8f
$���Vr7~�u�63Xgw@�Hy��#�����ȵ ���:�����#|��Ή�A�ݲ�N��1h�0[a�p[!�7��.�.�AԷ->5����8��hl(�����˸(��m�z�x�'�J�=zɱT�����΍d�s�:�M���oNzM�7]��$�r�Ŧ�QjhD�EȚ�j��*%�/Tu"������͡�氿�vLu+�!��P8�F־�	~�R%��=
�����˲A��UY�_v.F�H{�6�� Y��$	X��߬�E�|�� >o�(��CgI���%]*�$��o!� U���Dn�ļ3oF W�����W����m�L}%����(�(U�.K@����Q:��a�����2�VU��'I��n�&��
%yȰ-��}}Lu��h�6��Жd%y�芢���g�/_!����+�i�a�3Pu�J1$5hz����F�k���"Z �֪?z��Os4؞�Y�̋�� ��#8D@C}�f(	zF ��s�����XjΡ�@Jg�Y##��3��x��ݍ��s1sx#D1�n���wx&f���E;l��" 8l`KqY8��0!`�hi������ղ�����	A�sCqnVd���KZ���dPjȠY6@t�w�[�l^�\��Wb�#�؜ڍ��Y�*��6*�t9�
N. �<kB�o�_���^nY��S�m���?�<��~��N)#dY��t�n��Y ��3(��98���v��'zr�$�Ӿ��ϻ'̓���;
#߲+�A�\����YU���\xɫ'3lXJ���$��|z@a\X��B����V����M:1�-:�Ud/�Y��e�����8�9�U��lؙ�'̻�k��=yX&����AU���ϰ�v�������=Z\���ؠ�_��iA.��e=���ؽf�
��-���O��a���C�bl��<�p@4Q���{��O�ps�>`cȫ�Bi]T3��I7,t�6D����E����ӈ`�<þ�gn'a�7��RGmL��h(7�C�8��ǏmJ8�l`���Ƌ���{�����!Ү�'�jy
�F�P+�i���e��ϢaX[��|<#�����B@���
Ͽ)j(����/�J<��Y��k����->+6��zkU<v��X�,þo����NC%ޫ�;�ᎧX�0_XV\N������z��2��\B�t�%=S�x/��'�1#�!U̹���TAC��Q�p���Y�T.~X��R�t{�7M�{[ Q2Z��*n�Q����P ��Ŏ��l�Ì+W�9���� ���[\���:Ja۟�䑂�}���ΎK�ɪ�~���"�>����ꦄ��|����HRM��H��A�e����
tfE���u�2H 	���.s��h��=�`�f&�F��O2+l;	&G�$�eS��m!_-�5�����M�*��c��ՕL4؃�l�qL]t�^��RtZ"�f�l>>���w%��A8�^C�?3��{y��~�:+�b��A�H岉��3��7��mI
7��3�˦��o���UÉ���Ŷ�b��:����Y/�6(� ok~�2%c�o���n��O�����[2�%��	K/[��w�vlt�#V�%p���nM; ��
ra.��yuw?}�_~�	6�{hz�yz��:�3��7T��qQk���S�_�w�ϟ:{gcv&���V)U}�u��q@�)i��^��+8��Db����7X?L2	[1r<N����V3G ��-)͘ ��s��5��mo)x:$ �CAP�����mѬ�D�1S8�w
��}�Lƫ��@ G@��(�of%��M�A!Y�jԜmG(n�Q��n�����g�N�����'[O��(x�x3�?�h(`J?{yx�}B0Q�	�-��Z��2���������%���0o�fD⮺1�Gb����G���ΰ=	�Ǯ��w���jfJ:�!!#S�<�+hi_�Mv�1��_��78����'��=D���<p�n�U19|nD<)�a�Û[��9�π��K�Αa�)R��
�dց�0���׿�iv����.s�׏{�K=���l�%��g�Qd7�g5�6l�޵��$�ڜ��k/��DQ��ar�E�v�F��!�lɞ���:zV�K�/��6�����g����1��F���ح
6@ֿ>m��O{P�����|~��������e��Ļc���~
ސ�Տ}�I�nGc�s�w���s!p���[��X{�s��և��-Y|b5!�5��t'�?s�����7���#�ƙ����p�n�秘���'�'�І$Vn��� B�P��@ł'P�X�á�	p�_Q`�m�v0�aY��ǎ7�#wam�6[���3��W\���K� ��;�(ɞ$/(j9T�mS���(p��Q>o9rh�߲�����2;%a�W�O�,n��������������ݬ�A	"���;k�@�]�����G���OO��ʺ��%u��_���r#�C�/��?
�N�M6�I_K�`��G�KN.��������!y�P�Y--�!��kN�%;�H���3b���3S?=��B��f���ۑ�1�ob���_R��xߞ��gD�y�Q��Ghjo�3��U[	nRGqtY�PN�)��)%�oƻ<�
�݁X �zLc��,p푃w�B�h%�"m�s��p�ݖ����,g{���C���K�7�c��2f�u�����V����9��5�ݻ?���?��a���c��w۵d K-VY�!�ԡw6�I�����;^cR�k�����reG*�oG�r�/��ʅ�+8�����U�����
�@�a��$bB�	{b���v�H���69��@�|b�q �.g�z����&��%fD��Ǵ�b���c�L D�k\��1�Y^M[��� @��j��JV9d(d��g����ݰ��^��l�x�=>�Bu�B�G��{�P|�J�����Kn�����;�%��>ã�Ia�Vr�-�K������p��5��ǟ�/Hdi�j2�dW`�.���TG�KP���))��(����i�|۾¿��sѴ���hE@F�X���W��f���V���9�����g��zR�˃6B���5���1���x�����Ւm!#���A��;x3����<\J�"�N�	`�1����mǆ��x�<��;�5��S�A]��n4��,�m�O��|��P��� C�f�^fUq�Ȇ|�� ?;����r��l�g����6=�8���5���#(��oA��k��=wȳG�Q3�����-���1\�J	�V�g�b�ٞ/���
�U?|�6���=��}��lg6-G�%Cd6�>&�E
����5d8
�k���]�6�����o�4S����^��LWpr��:�����N����d�ϱB�ڬg�I���;�8_P���i�k��}7��%8x�p\^a�#o�֑�HΑZ�6�m%�
���r����������;K��0�~�p�L��oC¥��kF�!-M�dK���M�S��M�B�Ig�=���v���`�(_�����/�6[\IW��������3۷�0R�ږ����p-3quͲ�����E}�-@ӡ���v�Z2V�a��e��|Z���T!���W(p����rw���B�iĞ��+B<+K����ۋ}6+��^?��f�Y��!C�A��ï&V�%ޏ�؝��FbK��9�x.cW%���1-��l���
�dֻS�ݬ��7|jk��ܦ�uKJ78�Ю����	�i	�GVI֞�E���Y]3����p&�oBlÎ��@r;6�n1��H��15�v3�a��Gz���.��Q�ጢ�!x���)�=��_�;#
~}�
x��wo����l��d֋�z��B��q�?��$(�%�3T�,�6�2ǘ����E�y�6'X}�Y�����+8������z��F"�j�H9�z������ǹn�P�@����C���u��?�T;r�XPƓ"�1Ӵ�����~�B��#X�W|�� �ǎ3�d�����P�.�ɠ�bi�;Z/���5�����I.;��w���|�t����rd+;��w(��[�������߾�!!5�Ve���*��8�Q��-�uU�V�9P蓡%'Z�Wf�5��g��z���J6j%��KAݶx�l�
�{��)���(Xɾ��zxh$�z��n�ۮܮho���_ٻ��O�
ޚ��P"h�q�[���BqN61?�;X�5�%��6B´�1m�`�L�)B+� ��$fj̸C���Q���]@�m���,
x|�84�v_�����e��RE7���f�e�T� ���-������i�ln�q?����ː�,����ےǤ.��q����0���y�;��4o��^=y�,}� l[�_8�Ya��U��|�����h>��{j��l/�?4>M,��Z,�*'|�R���g��ص�yB�Fx�ap�������o�3����(��^���;����+��ᆒI���A8��$(�m�iL�LB�?�{ء�]���Ŝ@���
xQ6���m�Z`B&�
�^�.,�@+�=myJ\�s�����|���P-�ǲʶ��[�{nxտ�?��\��}d+�u���7(0ؘ��r=��}����Ȑ�!c��y	O�����{�f9��L�#"3�o� �H��@���2S�IV��l�f6����h��P��rVm�ј�Lm#�n-$�BQӪ�iu�T��X�*������̌���?'<�#�H�!/23�������}[ϑe�8s�TO��X��K���:��|���c۾��[�4�$@�pok��}s{l��OQ�HV�����=80�% ,��2��L�y�8/[�����5���Þ�!u�e����S$llhz2=0w�1,�^	�fw��V���$g	N��IYBR�;6'�<�L� 1i ��{fp81�ʀ�㰦@h%N���7���>�i�
��Ϩ��d�C
s�Gڵsp ���oh��j6��O2v�ޱ�~B�FQb��T'�I��/TD����[ 9����`�̰
�g�8��cc��\�Y�	�;s{kbFS�d�b��r>����3�%[�e!����^<k�.�lJ��i���M|��͗�t��rP'K@�[ǳ3a�Ӗ������4 �SfDt���[�B��*g6_�&�q}��Ԣ�b9�4CT�U�Z5��&�����ƊYMh�5�g[G��ҡ{0�ݳ<�����$	@�)+����e��#H�sbw�+�g�Q52�+��
ϓ�Y����Ԝ�ܴLol��-���®�{U���;�O��g-��LjR�>l�2�s���d`:)G���9<��p�޽
'Ȭ�-��;��'�nٻ��ŭ��K0�ȸ@fy��infn>.͹5�>�,������L�xe�I�f���2�[�OG��9S��2" �g�s���j��N[��a�>4������b���L,��{T���`vN���� .�ۓ�, ��A�l{�͆)��X�w@a�k��9ڷLߖu�Ӏ�#�`���m;B�,@E�W���.<���dl�YHt�nH�YsĊ�}-�d����y��: �޺C���	ٷ�W ��me>z�k��kF��"����![�,�z��oK2��,�[�``�0ӕ3��<�&�|�1�q�^�l���N�Z�7��B�� ����g��G���+AJ���8Y��꜑�I���<S1>O�8�فԦI�ekr�#
������4�͛�$Ǟ���p�2ቹu�cA
��������X&<��`p�!�V=�eL�l,9洣'	�ew��"�G��y`���2��CR� �h20w�Ͷe ;�I��:*� �!o#��X�6��f��"���:��S��ۓ}���Y��	v���<��j��e֖qZlaƖ��j&�����A�V����7ZP	�a�	c�ъfGfb����  8��g�!��2��" ����7�z���)h��2����I�>A����އc�):��G<ev���?� �|股�b��r�X`&��lDҘ��ɰ�Ȕ���#c�����	���-�k�=�� yhgɇ������p>"�>��f�h�ԠG�V ޚ�e2��X@�W� F�EF��c2�]#	O�@{��C�� ��a�����[��Ay.LI@J����2��ׇ�g�H�m�3r��=�p�	�?�[��1ϸX^?M�^�8�81����ʏ���� �9�N��`sL�؂^/�3�.�YL�b��8�x7��Ve�la"1N$PV�v�2��j�^~�2ܜ\4�#��0+����e$�ʦ�ʂ��#��!�I�����5v��5-�5�α���"iy�d|��pe��n��|`
)�-C�p��e�P�<)33Z]3�-{��@T��XP�?�1�����<kg-Ӛ�4���@��C� 9��8Ud'���Q"�)�������43+�� �m��:�8�;�=xUP�G�LK�3���kv�A $ł1��9�N�ZF��y�08�uV8J+�T;�+�|�I��0�C2����J:���K�2�8];G�[�he��5"��h,c���d�\�!Q��i�FcTR,��q>����\A�aQ�-����&n>���-��`$=�s��<�Q,h~���(�.<�H���4{��a�ϩ��K�y�<T27*�Vy[b�$�.���֏�}آƵ���UR�f���	�,%p��S��uj-܍���N��2�3_�\t�Q�qD���V�`�v�N](��O����ya�q�0{�h�]'B�e���tC{m5�eRS���1���B���h���[k�&ԬN*25���|���hl��p�N�5^�,�r�ٵ�au�A��oC���&tZ.܄{���;��buՂ�#j���R����H�TtM�ns��
HK
>�.� ��B�'[�EB��w�SH	��� 1O�1��L1I����-3�����1#_�,�L�^��=y� ��$�8Q�)��ә= O�b���$5{����4PP@v�E^땤S�$#0���\�W�h���>�%�8�J��ħ�X0%�{��4"CcK���Ըӛ�>D^�d�����*`���\ē��[�� �5��"ʇ�1dMPU.��J�Cs>3��ݛAO�$!i�O1�ż|Z�J�#����K�����=����RP�d1r;7|Q�̂�9S�����Z{]�.����y��2*"�;��-�f���L,`��F���&q?�v�?��A��Tc0d��`##�
�u/r������,c�C�����`�attD҇1�A�b�y�� _��@4ҩ�`h+�fg\qP7
J ���|*��2�#ʇ(�8h/�;�餤�<-�00�!�t*b�w�nAqS`�
v9�حeL-�]YQ�����@��X&�1����3d��s���{������E�H���&IUq�-��.���������E.�r�;�l�/w-�8V�q����O�&s籅k�?\�c�X�p/8�H�DU�It4=�m/�\�,R��< G�)ǉ�2~�Hܜ�C�Ol��AH�"#��G �,��?:z0��3S�P�c?G�5z���G�,���]��?��/1A�K�c$���zO���X�X�>����J@��m�LZR�ދ���y�N���|�V��� �&����q]7��W:��YC׸k��%��b�c@���qtL&�~
@�A��Cn�+���2�iF��<p��L�TP�#w����G�)��	�����e�qT��xg�F��U����+h�SPpKr���yd��D+:�;j0A �U3� �)hVư+��D��΁��)D���r�!UA'�BUR�����9�v+d�{�f�!�kF=b=����:�Ap��|.�P2>V
�̜�?�4���Qd׌O{��,���:s�����2>�IM���*����$�YIcK CdW�V��ȶD`�	E�e�Kg�L�c,����d9Pd)��i���ر"�\M���P9��B�F�9 u҄��T'd+���)?'x�j���nQx37����\�XH�C�� Y��@|����;����{��KH��	��mJ�=��kܧ�>�:��)�Y�8ݎ����)�E��3�7H�d	(��%!ߕ8�Z@Rɯjh��g���u�/��O�w�xG	��d���љ)59�6���;S�+jX:|�ߦ����-TY�k� wN���s�-�S��<�>!��� ��ׂG弨2�$�Rs8w>�P�~�yI2Ts<5�FZ�Ǆ<���L
��~	�U;���� d%/ݧv90��` �,s�{<n4W�۽f���Y��S9���I����8�=�V�qw*:�_4�\�S�ȉ��Ɲғj�Un�+���8�ow^5K�x|�бـ��P= xt�X�d�Q��#(�7��iX�E�K��Q��g�T{9����p�`�KK8o�}q� �n��xξ+���S��I:bt�0 �>2��O5s/��qy�?�蹧N��jZ	�0�O� k�OIܹ����y��/Bs�UX�,L J����lPT̒��f��k'!��L�lH����������Q+��!	�f��r:& �ʁ�ҩE*:�6wͬj�>��,�+	¤eh����l�=L�tbf���2Ru�ٔ�� S�J��j	 5:'��J<vB�;w]���x:�iGQ�Ġ+�?j�����	b�P�:s�0 0��sg�q ��G�4G��q���ٲ���X���8��	<��u�v3Y˼��b$��)Gt�lc�n�f�A�敀^��Ʒ$P3h<�Ƹ���I�Xz�#k��{��]��17d��L��;�+��A���[�>���A!�34�!���EW�Z˘g��&�-�����D���}�E^��e�N��f_��EΚ��0�m���ͳ�﻿��3��rC*]Ь�Y�M0DRQ���clP�z|�);ɉ��3C�zI%����M���&#r�@�qݙ�E�Nj��J���\�����m)HC���̎%.e#��JJ�6'w A�!"gc�Ԩ����4���������X���	(���,�iH��S;�W�r�ݘg�(��)�1�)X4��#���e-�N�f� ����so�8��*,��A�$[΋TWp����4-�+ء8c�s--䁆�������rjz� �O#n��,s�s�87X�i����6;��[��P�4h�y�-*)�5��Y�n��v� Jo���~��ɒP'K@�qi���B����1�~N�t�EwR�-c! U@1�y���|6�,��.�:W�p����&n�.�cX�a<��n��{BR*�T��M��T¸3��d2QGN50����+�+�3`Г;�ޒ���gr�#��\"�5��L��5����*`�6;�Ք��b�`�Ӝ��hs[FV��Χ�:\�qHG�'F܀�,w*�ڵэDfH�臘� ��l;pp"�q��X���,�j�jM�*c��m>�3�x�p���>[�Bc��N��1�6bI��P-��te�g�yV侨����������8���+>xh��ɚ1"��<CJδ�A�����OK��lO�Z�o�_�oī��ɴ�*�Q������O�`0��Rf���rA�*a�.�T���~���齟���ѿ�ѱξ0lΊ����1QtT��Kj��T�����4˾쎻�����L*j*R�4��@%���ԍ-	ٵg,~'�,ol
avX����00!�L#�*��ߕ��M�#3R
�R�9��ReH�dΟ�F���~b�E3P��Cy�v1�L��4�mB P5KOD�&R/��K��LC��8��WdkR�znJ E�L���ɜ
�6��q*V�1�`Q��ܴj�uMqH���\�sRS�mKeDZG 4�U倄j��1��/�/�rsX4����JO�+M�����Y\ל��i61o���}�#d��f�6֍��AU��L��F���P���BN��S7;�����'�ں(0Y,�6Pd�}���̀���Ե���R�s�!1u+��pNLP�zk6�m����i��.�ݒ�FX�N�t�����G&�Y�鶬�nw�5G���e��H��@[�M��CE6)$9!5�2PC&L�UU"a�k6:Ցq̖$J�J�-�mb�
��(�,�0R�~ve+g�LV"5K)���+�I3zQ�4���{J���r�� �Д�N����C*>��ZilH�/����1<&ʛd�����l��@�:��i��Y�`k�iN薋��RM]����T��\��ٔG-�K9敭��m�%'���He��@
�Q&p�����OuQQ
/�}���E�۔j]��v���*�q������eA�T
^�D�iG�Ūnv�b�و�����؉ԙXx����:q���"J�F<k
q�5���T�>[84�p�)65�@��$�WGV�ZD��ک����8�@&�	-�b�fU��[US��r�{�f>p��oT�+w����60�і2��AE)=r��3'�ZyA3����/�i3#��r�Ά���8Ԭ�����k��W��&�μ���vH΍Y��2��A����!�"��Y����)NM�2�����eN��2��4�R1��3�q��ʉ�E>e��@��4-�Q��{�^�Nq=�Rۘ�I�HN�r;�$�( ֿ</J�:��D�3%p�4�q1(h=�කe-��٥K�I�>e��5���xQп��T��_ ��ӗ�n��.�9{.��N�!^."G5{�Z�)�9)`�5��[o��q��I,�0s�273�+���"���~�rv+�K�M��f�����.6F�H��5%a���I��H�ݵ�x���R������;A�r�@�����d_��겁.��������9d	�1
���Q�����w�6�"���!��i$n<�aG�5�N��Λ�)��j�z�k���~3�5�ӗI��v.\����u��o��~�/"_ղ(�3������d���d	�HJ

v`�M�����ёI�乧N��s\��h4�N��`:�f��0+ˊ#{✖��c'�2E 1���)3
���j�w�Eؾ����uc��NѬ1�z7�S�1��0C-�Żl��07v���d����q�q�W�;u�cb�l�E1��.��p��"��[73iES�c�n�,���-�X��)�9wv-�ȼ�f6�ZeFX�i>3��;�^�B�K�1Gc�,�f$wƈ�"���
~0L�0�k'++*�Q��UC���b���	ȣ��yN�Gc3D���f�`��Q�XzFأJ�##Y3Wy��ё�j�Q\r'5ˌ��0�b#ٖ���8���p��l�$2�ʛy'��s)��al�Nt�r~G��E,2�S����Q$,�۵̧�!o�U�}�j�B��/��="I'�Ҵ+qh��1�u"ɳjX�r2���M��Ѩ �Y���G��+����N�{J�d	hmmm�.J�ڗ��%'����]֊���F�����b�뾫��j�ZCn��{���Pڤ��s5���L-��c��\+ö5��S@�q;e�b������c:u�ͿM��ٻz�t��֦E]������CZ�Kn��R�H̠sb�Eƾ-\���g�TǮ�S7�Zg��t�''1�]Ш��(�a#�G������֩����a�E�� we���{b�-M���~v������z��Ce�y$Bk�X�e}
��N|{�Py���m�Ж�� R�t��/����o������Ο?��'Nl\��ܼ>��e�G�蹥N�s�u�/���o��������sx�ɓG�ܽs�Z[�ܬ���C)J��$@���hi�[ ��%ޞ6}6�`��S������ '�N>��+���zDc��^���ko�b�[4-��JuE���w�'@�v�X�<�ʊ1?��_��vC��Ufh�� V�M�A$��W_�����=ڱG�n��_�c��7��;���"m�7�������ї��o��Բ(�U��G��'O��S�N�W�^ݲ�����'������������?�ah���9�N�����p�ڵk����x�N޽{�ч7>�>����x��F��j��ݝ�\0�ѹ'�љ,r���O��|���8|���+�'c���2�����b�$����/�&$��Wϕ R���3u�� Μ9�Ş�?x��loo�Ϳ��Y�S};�gϚ�'O`���2�?n�|���"V�ԥ��o���0_M}�i����ߧ����&4�}yci��b ��+ib�)-�C<5<�,���5��H��s
��#��d�(��% �S '���?Ϸnm��Mwvv�%�I�����slw����f BZ�b����$��H�g����g���f�K���N���E󆀄\��Hc '1�#�48@�����}�^H~�m?���P�$Ɨ��� %�Ν��;;;$���.Kԏ�M~]�A�3�8���J9�݉������?�q@�/��?Q����u��X9��J����D�Q)��8�I��HH�P&K�&��Q'KFv��a~�X���	��`�`�ۖA���ZE(�ػ�(��4qb�'�����)�X��cbi�~�o��3�. )�I�$�t~������?5֗:H���>�����Xh�*��������n�����E� ZTL�j���{�nOhW��/:'�H Bc=�Jh)#��P�j>鼡��!��k����g�`��:�غL򒥤N��p��f.t��Q��C�q�a8��;�v�=+Q��f&/(�L�f�'9	��ۯ��]XÇ�-"��b��Ӽ:Bs!�ڠ9�0B���<�<,����yv|`�N| *u��U��I����\��������S��Y(M(�.���>Z��y EoHB��@�_F췾��~�T���Q�4���S�Zܦ��p5EǾ{�$Z2J�d�/)^V�_�0�Ʃ�Y��DH�yu>8�Y4-�?�Vl"�0���]����Jb�ps]8�@�N?��Wl�u~�w_^���ݳ<��a���Ԥ�����>�=1��� ��j)_KN�!�gS�_-����k���0��q��� ���iʖ��<�����0��ȋ��y���ї��w_�C�ݶ�z������SD�e�N��.\���Uh҈��9�e�,z�Ћ�ލ��}+ʯ��k����Y��2X�WSlc�!�۾����u��1���NB�b�$$���1c�;��> q=��Ql�tX���D
��㚀�CX':�����
QHrb�� ̎T���硴�gKω�{LB�G���}��D${�ր4X�r$_�|���4`�}�GAH�D'�F	�,�E�yL�\��LxG�y���A(�X�$~Xi�9��ȥ�a*}����҂��eH��'QA��P�������4���)���AI�)�ۍ�ڍ{ '� R���u�xLp��9xM����LG_�G�}���&���y�c��\�IIb���м͓��~�л��\D��&殺h��
IPc���[��6%�<}_\_�"1y�s"���ɿ�$.����u	i@�:q<�,r',���4���І�Y��e��=��ە�����OJ1��:!0&��@�N�{���O>��E_�ܧx 5�=������3SB�´��/��w�!Ư�ǀRH��S�.?$�WƢ�Rc��$f���>�ρ6������s利��������D�I[���R@Q->��$Z>J�d���h����2��uh��X�Hb�L/�|��nٳ�S��Iʏ�L��r�=aF�6��T���(\���&1��<I���<N[bs�Kn|���H�Q�)[?��g�+�I��1�Bc�Ӽt�
�6����>�[8�����\듨�F������'����ݘ:>�s�O^Uu~��E�h�(��%�,++�W!�E�r�gB�|&�$)1�
vŻbK*W�ɟ�����wr�H�ܯ����R=�}`b�*��	-�1f�7$Y
էۭ����O��貴$�wG�wӱ�����g8Y\���:b��>���1�����f�~:D���A�b䚶Q��>����+�����f�k�,�k�˪��D�%%p�d4�^��ӟ�\��}����-�}��%�[�<I��]��}�׷�����%?�/��c2���x��w/&���.xB;V��P��cL����*Ĉ�6j0"�>O�PYRO��j���+߿>o�ce��\��ǘ�<pk_�M84oR��'����_�o��U=O!�L�y	��8gI�e�ȥ���=w��ɒSw����>A1F���;p�-�3��JZP�i�b�P{C:���`0�8�E|���I���\���GL������=#�N�,��;�5��cL��M}�b҉Ey�"�M��8�����z,���N�du��s��$i����z\�H��~��$W�e�N���ۗ���	�DݝN�8N�(�0	�>M8��E	�D��}�F�����w�V_Y~޶-�o�~((�q��q�����@�y���ɗ�|�"�
�Z����8n��OE�󁪾��#NB��:�/3���MCL�~�e�Ƶ�M����󬆀�$Z:J�d���ի��~���v����_awb	H/��H�g$��Ԍ'��b^
zA��jU �Gj ���%�ے��И�C�uJ�v���s|�cr��e�!�4��Ů��W��k�˼q�=3��XB�cm��5�-}�}Q��yl\��~���� S���~=��G�mm�>�l���}����;��&�1U��JH�T������뺕4��~���.Ɣ�v�@3������4��p IM����D�.��~�˯>��_�xG6D�k�c��o'����QJ%���k���AȤi����`6=�Y֎�_��d�Y�����dtDX}Ju['ǜ(,�(��F��N�F��O���?�G�r�_�9��C�O�\B2�-�I%�#BiH�����c��I%��V�B C(�\�$~�!O���.�=�ey�@</=����߷o�6���8YB*
��D�"U�U�nrfh:ZI��`\��iLF��E���-�[P2O�#�������4`�-��,����P�9q�9<<�t��Ő�yq8#�ԅ�7��ۦ�͵��k߅k&����j�!��3±`���#�6�H�j�vaTr����U�1g��S������g�"�������)��/¦���QD�ؙL�ލ������rH�+O��I,��X�Ce��ɢyC���7� Ơf��?��e9����rR'KHu=��L/�^hC���Ss��v�L�� 4�2����~~/���h�-�_��_��UI�k��Ov�`���2�S�;w�vt`n`r �_#�q�����o:-;��}�u�T�V��e!��H���I��|�	�������d +cш��������!A�������� dh^���Y)�|�#�j�/�a���ɓ���-�C\�����z����]���ׇ��ؽE�����F? �K�k�޼�x�q嘠������P��8Y2z�},� '�D�^-pbf������>��+�P�`XZ����S�x;L��1}��/�G�L�ԩStL�D*"���V�@L�Cȇ�wǣ�?����I�p!!��<��k��@fmuݔS�spp�i+��5��������3ϗ���)��3|�1����I$E2/R7ڬ�+��9ß6R��]g$�����������7.}��Elz�M�^W�E=F�%%,��1��RCܰe�!b/��r'KF	�,���x���]@�Z�'U����BKlG�/	ٞāD{Ϳ�_�Ȯ4Ъ�$H�)�766�y�����1#Î��Ç�5,�b� R�R�7ߝ;w��G�mW�+ƴB�[�F9:c�e]ɏ���|}�� /�� ���@שU^Z�??��K�:���?O���n_Ϗ�*H�$LTR���ӧ������P9�T�,�}�Z���p�,�ʍ���v���<�҂���V�57O�����?6���8Y2�v�Z��_\�IQ��
i��F)����f�}4��گ�����[PC�Z�Ђ�v���ռX�?�|������-��!�����Pz�'�����Looo��C����M*0?�?��e�a櫩U�KZ������b��ɓ�Hҁ�jР��mSx��+ ��Z�/��E�9�= 1G���W$ !�u�5�q�6�ڳ]�R+�_�C��?@�/��O��;TF�w�\����/%�O���&m�NUJ
,sf��['�ߏ'fK��S'KH�)�W�T�y��B��� �~�Hl�-t����������_в��p��v�zWc4¤@�.�:R$A"cU�/�@��!����ġ����K&� S����[;ݾ��%LV@�x�H0  !��h��� �΃:�1ɸ�};��D� �?�휴�kr��08~K��T�&�޽{4Oh ������4��1D~I�O�]D��P_��.Σ����JLJ�'A��$�i���UO�x�����8S�$Z*J�d	idrС�\����E�'}s�5h�|����<����W3�ϥ
��-�1�L�O��,����C �0�v�[[��N[[[6����}[]]#�$�VCJ#F��';y��f  �l���$Ĉ�t��^aհ��d2�m H��f��Nu�Qk_#�#�i+�@Z���SK*< ��ˮ�ϑr�/]��?o\^ٴ�����q��èu�~�;3�0%��yC�A��>}�ܽ{��>C� R�h�Zm�S�\T���\/J����V��k�"`%.)rRK��K�dI)��%�j�/�,������MpW�@@��]��&����������Κ�
�ow�_��/���C�%�����J�'�&��`�
�P� =�vw����dF��R=f�	�>	�B�kZ��*�VB��TE2R̔�w��t�{�n-=I�ԩ�����a�I�K�t�b�9�v����%�{E�Ţ �!i��u?p�Oǹ-�w'�ޅ6}����s!��ߞ�<��H�岁j�	~X@� �R'KK���5� s6z�l>��"%��"<�r���=?�\�͘�7��"��4���I�`�
E��v��������\��ڰ��E<B$^�0d-��m{|F��8�1�� 0�T �]�پE�,���|��D��[��ԥU?�n�� ����.�0�.? ~�] ��0�"���k��Ү� ��+�.M�㯟� ��#�^=�]?�~]B1������_�F!IG�n{��yu�4Hi��SCf�3���8YR�;b�uťn�q��̂i�N[B�jX�Z�u��v�~Y�rј �j&�&^�&��O�r_T�/L�g�>��Ӑ�@��Gk�J);�����������gOTVr=T����6)z���I���Eף���[m�Һx� ��X���ǰ���]�?�:�_Oh�4�e������Qh���Ͷ3^���׬��b���.IN��8YBT��ȋJ�v1����#���k���_`Bb���y�'��3�����\#���Cy�$H�:R���Y��2����ej�)ۖ5���6��LNd{��^��c��]�E
Є�u���X��tȸ�}.�1�)ʹ��<+f^��}�?�d�9��h;��,�$~*[�� ڏ�g͗�}U��Ec�D���v��_w��k���/���&�q:>��UG*/���u��8Y2��O~B6'ŀ"'��!�.�ڙe�D�S�9��E(�;\d��-t�h�BL+T^�P��Z�?�?�L#V���߼��H�W��Ÿo��0tqǼq���-�i��.ơ��C����6�e���1�L�?�؟���1J=|D@ݴ_ש}u�����ϣ���Hf�m�=,��O�*����>廼?�<�!�M8�"�җ��K�͔��J���$5YRJ�d	�Y�W>��w3������~f�c1��.d��j VH�х��`� 0j���)� A���}�d鳨:|�Ҿ�v��2�Y��7�Zk��6�*'>/��-3�ֶC�*� f\͂-e	�:�,����*:_B&����}�T�'�n_��5B���(��u����5�����韊�1����e� �D��Y]2z�w�?��1Y3�uv1	���f��i�9�E LH��߽�5 #,�n�00�C��e����@l���6���Ԥ�R{���T�l} �r�}n�4H�}�R�B=/�1�����D��� Z`.����	��v�'�y�{N5PHۖH:�S=�O)ח�u�E��@D��噭������踛��4s�Al��k���DKG	�,����Kd���>�ĪΗ�1F_�[�5Oz��?oIY8iS����F���D6+�j� �\�~Hx�<�*���UGZ=�ξ��>j���_kў$�|l}��o���sV��S�mo�����<������ce���t?O0��t`���n�ф��%I��̾��ˊ��_���oo+�k���D�I	�,)��k�i�mB;H�/b�6|tL�Z���ڬ]A���]̻���Q��%$~��YȘ @�_�f� &����ǁ�.F�u3�~��#xZ�2,��&��K{���]�)<�sU��K�	־�F*��mx���	�L���$#�{G�cEj���Ձ�|I�4%�NȧPo�a�f�I�b����������/�^_��ny�o�˻��_��YRJ�d���wM���ݴ�E�EO��,�������5���n�˙E���꺅b;\���6�{ӟ��9�Vc�F���)j��n� 
 ���L*^�_1e>�-����.���1ͮ{-�."eh��}M��!��ҍ�E^?���C���\�_Vq�>�GGS�1I*e<�>':��~�X9ļ�,+��3}k���̵`\�P-��1/��߃����L<�43���s(W�F���ws�G�=�r/D������E��Z:�;��y��'_�(�-@�1��[�ʕ+	�,%p����d?�7z:�4��:$C���^�*h1�//�j��v�ಘ�N:���ZHʡw�!��P��w>���ϽYq5=�*0DrE�49SE�q!���榋m2����=VK��	��c��ܫHˁ�@���.�>�S����lӉƨ"E;y��� �ܵ�Uj���#g�hwq�?0@���3v�lK� ᝳ��C�l��i91�IIҗ'6�� +�R>�2x�:i�ԕ9 p4�q���J�m�6���ϭ'[����fl�(h��ⓁJ�N��1Fu�Y�j��ЌLe��`o�ܺu�����(��Ị̈G��0��/���3s�z4�;��M�,�l%�$��m����g�2�37o޲u<�#0�N�6�Ν7'6O��gN��Q=
7�4��ZP��$���籕p�S�Ĥ�:���VJ%��R�>)��J�S��΋������d:�x^��ȲQ�9YBJ�d	)�'�]��7��	�v(�k��Ĕ��Z���p&z=�0�;����_De���ym�a�?�����57o}b>���k����ˆ��������t�R�G������e^;H*�gP˟  �7���}�3��>���$����@(����ͫW�)����uUw�W�B�q���5>㧴uݶ��&�}饗�p40�?��|z�S &��/�_�h��	��_`�ϴn��_�.�AYр&�9A_Ї���nJ yύ�.��g��z/�󖉷A�*&TO. ��+q{���4�\���-�����Ν�4���ߧ�q���Ӝ�����nw.�L�Y�X840w�	�L��R=8�7ׯ_77n�h��s� n�<~ln}��c����>_ ��������>�<ו��1�6�)��/*��IK��m���̶��7�u�?�+�t��2R'KHv�Yg��7� ����+�. YSnh��a����Yda���s�/�x�Z�ɀa�Ȼw?7�ܧ�����K�.~ee�b���A�q��9��6�	C�!;{f�Jr���(3��m��� �Ï�S}����t�)IVP&�mo���Ǐ�w��]s��	GHId,��7��_$5 Q��>��=��76�0��=A�?yD����}"�����/����]:���_�����r�`�>��c���M�x���?nTP}<� Ҿ]���- |���s�E ;YD�Ç4�y����{{�$� ��`�y�Y�'������8�aA
�[���.�o����Ғ��F<pҒ'M���
�o2�X 8�4��o{��zqЪ�Db"���QP8�Y��<�Q�7�!���n����8YBB��,+j-��]�\���w�:k� �u��t|��#[$�"�N#v �ݾe~}������6-Pm�ɂٱ�mI�0XH5���	��t�m	�;8fJ��v&�����G7��	����FJ��Q?�;H��o}�l�o*�	&"�`�C:��!PƯ�kb�'N��6@}u�nN\�H�q����-���W_�vV��.�-y�$64���/~n>��C��I݂2@�'*R�\���(̫��FF��c����ƶ*c{�_��4GP��9s���1�12p�ѣ�����Y[]7/��rsvP�Z���Hm�?����BR������
��bۜ��/$fP۽��[M����~w��Vͪ����л�o�����k�r�%��,��U�֪�%�ɒR'�GuQ@�S�xqe�'ԧ6�� M��l�Vn:��EL$,f�1��i�*}R���x0l�:���a��î �����
�.�³�dss�2�!1^QS4m2��2����`�`�`fb&�ﰅ ��FTl��h��7�iV�_�)�}lU]; /�qk�	�=N�>eA�Rm�����
�,��ѯ�+s����5��cp��AZ ��>��T8����aQ��Z'ol�P��Ǐ�N�왳��gpjf5.���1~|�+s��w�g��IĘ�5^/$�Tz�9s�lS��'q��Uz�z��`7�F�ܹ�v�^$i ,���iT�	0aN>��~+���<��FRO|�0��߃�(��ى���ǡ�<�$��@��J�d	�.�36'ݝ��Rf�bsI�.p�gFsW-PL���ٜ��Yt1-tR/�ݻw	� d��!����$��`�&� c�/�����pL�B�Ju�M^��4A�Cr��͏�y��T:�&�1k��f� ���<�n�"fP�=L��ŶDK&�,�:a���]P7�+���Zpy l��)��a>��S��o������@�!�h�*��7?1�v��ANF�(kgg�T ,ʜ��zJ�)ȇ��w﮹��g��qj,[p�����ˤ�z�؜={�I��P}�7���J������;w>��=}�tJd���
���p =���p�q�o̗��p���ƴ�א�敗_k���{ϼQ}�TC�>X�l&�Kn|Z5ڝ@_���K@B��9J�d		�K�PײP� D!�	�^��W_��۠�_g�[4cb鶯��0v=s�|޹s����z�u0q�q����*-���H
�G��$�0\���
3R��>T�.�0r�����/�H^��a���u���=�jR3@�q��=2��}1F#��5��ئC<s i���?��|�k_3�´t]������v`����\�w@����%���~ԅ>A�E�0p������!�R`G���wH� �!u��9�yd{Hm&�lT l^���Y�`*��R�6�:�&#;� rh�Hm P�v���?�xjOw�	��|����:��i��q����ޡ-�6꫻O+�h�  )(IDAT�#ҷػ�T�D��J�\�����ɶ�x1�_��T;���]�$ֆV!�HΗ�`����X=����6۝5<l�i}?﨡r9:ʈi��X��n�Pu���Μ>Ӊ���͌>#)@v� ěL��P��1� >��9���0R�9Ϲ�p�����ɝMl"��^H~ n�>��R ,��8��	�L�b��T.����6�����!f��f=&���ƛ�Y�m�� ��Cy��꥓'N;�3�Aڈ��vxpHRH�^x�<�Z`�qx8n�mF=�S'V�w4>$���  #�8�/8�����4
s����c{�.fd(+���n�N�mpu*�'���X��>�����q�/��!`��1ֿ����>ɉ]K��J�:�H	�,!��/�;�,3�d�K��/�i�0��u72f�8�����e�����Z c��<Ғ�A� )���%6������mH #BL�����6Kz���fݨ��~�T5�M�0������wݨ�W^!5����'LP��T�	P��!��<�jbJR	�Dww�Ʃ�Z  ِ_�5�x�[� ���c�@� �p����suu�������3NU6�j�V;Է�wd>����oP|�#F؋���	0!�ט%^�Ŏ�c��n B�ߐ߸`��D~�B߼�)Im ��g��Y�>�m,�[N��3N�=�!@�K'Z`4��w�!UQ�>��.#\Q�pW]�txZ�Eu���P��8YB*�ͪ���b���/�>�N�k�*$n������i�1�/���� i�7�`�;��/K��#������;L��gi�!���6���7�e*pŽp*�G�Zŭ��H]��b�) @l@p `�p�E,�|��S��	�QQIdҶ�\����1�P�`�b �2��8��;w��ctHdV�,m�#�R�T9y���/�c�ͻ��y5��W~�~Xm�O�C�O�RVN2ѶĠ-3b|�|�+k�I�D:�ϑi"ڲ��?���l�w�<sl/c:�7$�R.���ϰԥUu"}P�u9��v�	��z�
���zB�����>�Z,;��C�3&EQV���I�\����}�ʬ�p�֏�����MH�`@����	�ןF���4ieA퓾�VdP�!�MD��4��5@L�Ǝ��{��_&0 )����bwf��SX�f�A�Mg�� �P��'14��A����H�s	�2��@} f�u�"̞�\{;�zN�:c�ܹ��KH^�c ��M��c�''�wu2�C]x��Y1ƅ�g����p�H�$Ҭ\P:@۠`�:�H ���F��#y�i�*�2�R��/I>�[8ڄ<H@���I�'sҪ�j'9i=���� wg<��z���/�
�]�m"�������M�ڮ�V������׮]K��%�N��,әZf�L"�!�m�>ۥ��*%mD��Sfu�-$�5ݝ\_9ݶ͖Mx��`*���wE�`)�l�̓'ۍ'�����nSG�@�>�ݖ����7ȃ�|�9W^-I2$���)�3DM$�A"�p��)Wu�TT%fbG����N�ԇ>��>܎�F �pZ[�0�^|��nWW���
�ѹs��	��p�~�+# 6hÐ ȤpH��"�;7�쳗Q��C i_|�{�F����ws~�L	0iɴ�?w����:�)�)?4�ـ�mA$������aɛ �v c���6��7�2UY7 �U����wtQ����uճ�����9.�����&؝\Ӡ��U�ٿg?��{�N��8Y2�/j������.���O���H���ٲ�8�g�n�e�]}��b���_ן!�KؾaˡVh%���2�Ȧl�	��p��	��#���0&���A�r��MJ7����ڐ��W�#�|�2��sp���8��f
��6lbn��jlk8M�H�Bz~Vǰ�
܈Y�4u�ª��!al��ҋ�).�Çes.�V���� ��{�(\�t�"�N&���؏C#s���믿n�߸��t����m�-�pᢹp�z. ��H�4�e$=�9D/^�x% ��:�:���y�P�/\4W�^���.��V]�7b_��6#z�C����uv���l�1	��U 5n۱��u�C;G���n���D�%%p��d�iQ��]G����� C�jwv���x���0��]�H*���ґEh�]_�� �&�ַ�M��>��S:T�(*@����T
bv/^"|`A�!�Z�_��3���)���xl�\�BA�n}z�A��&�/�0SX���R�z늹��vH9@\�H|�l��RVO ���̍��m;-����;x9h���FFu����q�[��h5����4�׮}��y��qߪF� ��l*��ɕ�^'���v&7�#c$��&j�)y������n�6L�Y�R'9��l2Sw���ʚ��7�A^X�[�Ո�JƂ������¯ٶ"��?��?8�t���U�*�s�{���3�eo"9�����XyzUOL�{�����P߻ڑ�*I�\�'�e&'Nl|����)�I�T������Wkk�G��;:,�3B1������.^�3����VE�	�u�`P���<C���Z����XJ;_x��8xe�P#cM L�^d�������ǔ�������J7 ��>
�	��h�jU���8���l@N�<e���o��A������ ��o��F#��R��*x�9���/�d���kd��:��EN3���9�*�!x�\�s��Å��Y�	H9lm�6����m��'4F�L;"�S��6�i��N��:_}��ƭ�=�56��F�(�};��y��'��7�S�ڳI�v������}�^�X	0m��n~��1OC�H0��i���o��Mb�# ���-�ܷ�������$Z:J�d	�k_�Zi�������8�̔����8�E��v!��DSXo]7B�E�����xbB��x��W���
�|���[;. ���ߣ|X8񧽟Dr"̍vĎYaG5ҥ/�������~A�Ƶ����W��Y'��ŋ/���9�j�cؐ�8��A��U9��r��5*�lwLـ
a��xWF��j�����R��k���gZUڃ%���_���!#�!���� �l�1$5�k�^!@�3g��[#c�\tm1dN1�G� ��o����O���O }�m�8?�ƶ8��=Hy��C~ygD��v'���d�N���&c\�8��(�ǎ�?����x�u���7�:�:�Uf_�+�HC�|)edm�E��m�5=u���E�r�&OG�-!%p��t�ʕ�]?����`��V
,�}����Duؚ$�!a�rL`L���4�Y�5��ۨmI�`��C��#�L��28���l�X.X`IT3�^�X�KG#eӟ�T)��`wWCA�`ǁ�i��m��x�H���K��N�6�� ���Hfd��[-�'`� �?܈qV�9ሥCۇym�D��+'���Il7����I� �����7b� ��NDV���`\Q'l7�\y����~�c�$*�f|�|���s������t����2W "�w��Cz�[}���Dis��� �[ۆ#�#0)��`{e p�>u�>C�͋�.�k6�b��ɿ4P#=V���A��ާBj���5y��� ����љ3�ߺu�����ui-%p��Tmm�������^�/u{,�`8,��	;.;�v�oL#�����c�uI��Oh�.z���SX"s�41Qul���=�q<��+��J���d� A��рb_����30Y��{�nSa�b�
u \O!) 3�Y2h��"p�p�+`t/�x���}9U�9(CU�W��D�#*���`nx&П��>u�>��
1m|�����4J�u���X�c�JP�=`4�\0����y;��f �z���V7��b33�Qԝ{�B_�N	2w��Is��#�(W�t�l�M�H�!�}�[?�������]v/����	�(H�Ж��
N�6h��O�^xd\F��y>h�/ĮF�ե���ǁW��63��Ne'u�B��K%g��U��u>���#Ċ�x�$�G�ұ�o߅_��֛c3oqI�\R'KH0��������77n\������3��H�"�ɹ��u�3[#W��w�_)��-u'�K }�cQ�]�" �chG�H�FÐ����y��!K٫gH�^q�S�8����}.�.U�D8�e3�`�����'���	R� T��TH���ƨ(���N��QtS�gm�sq�����r���UV�?��V�NVRQ[e���"}���[�N���ŋ���S�<�Yљ����4v:Z2�w��awW=����x�h�"����"��=�26\�i�vH��4�>&��z5Б?̙��S����h��aTV�=�Qu�-�}��;>����8�l�9�P��t%�8"b�� ����Ӎ���׮}㧷o�N�dI)��%�w�y�<��?����ߵ;��vG:�sDƴc�ŔE�rYe2� ����S n���Q��S���ڏ�.�!W�����t�s�bWȢ	&�'ߥara
���s[o�植�`�@ej4L�a3Z�I�ĎC�ӑ^58�KCj]�ψ��E�J;VNե���\��~�X_��3��z��uH�>G�'�K2�ڀZ�w����y��ƤO����<=���P ��,�F�4��%09,�6*��`�e�>s���ٳg?�t��/�~+y�,)%p��T���K?��Wj_���y/9� @�����_Xu;���/>���v�! ����&��e�t¨��Abs��fQ]�fξ�_3�ڝA���S����r�������/6�r}	����+��'�ğ{�-��gml��F�z�T���{���^��@�CH��%PS�G��ӷ����Cs���'m�B�kAS�qѐ�J�+y��jLA��j1�W�O���<y��[o���������N�\P'KJxi-=��x�>��ɿ���>m_�vPI�y#�K���~��4������3V��o��e�^A���w�2F����f�O��[~W�i�:�fn�~v�yxL�o�ܒ�D)vO��K���]��!����u_Z�T̤�}��?���Q=����@�{ru,�E����D�7_�J6}���}Z
=7���a\E�Ԑ�X�Rٵ�'�o}���D{&��R'KL�e/�����.�m9�^���=�	^t���&�@�Xp1��;EY�����o�w^|&9�LDT��z��O�C:�\��5���°$��!�މ�Έ����5He��g���X����1�!|������K��N>$M�I��Z;&~���A�E��Sv��(���
����/�-'o�Y7m��ϣ��(	�|��TH2���uZ��1�i�?��RZ>�5������Վ�ʌ3��R ����{��z�?�w��mP��d�)��%�w�yc�֭������w�<yrb<�a	�Dxȹ":���	u��V���`c�!�:��H��|�fV򠙜nx�!t��e
��� ��9�^1N-�_�b`��C�9�U�?��e����N�yǀ���%�.ïo��w�6��U_�����R3���S��nڰ#F�6�%p�h��P��EA�?���c_�&��'O� O�Ǐ�}Rm7Tw�\��_�]����W���&KN	�,9ٗ�~���t��_���9g_��� �F
>5�q�8�n6~CSF�I����H���늻�o3�y�>�k��7f�h�_�N;/�	15@���Y�o[�3�>����$:�$8}����HsB�=Ծ��7�9 l��/�k���$�g�o�C}�{����$4��*�חX�"2Qm4�=�� Ξ��g��ؗ��Dd^[_%����c����H=���o�G��zl-=%p��o~�7?���x��������q<_8<<� P�*�����N�Bx���.�&J�A��A�-��bh���-�����rbV>cR��e
,���V�����$'�]>S����1VB�Q����bt�ϓϰ�ZDK��I'ҽ,[$�s��5��~��P> ���Х��d����8��n��>�� P�Z�u���`�?Z���'�4���Ν;��������?��w����(��� ٗ�Ⱦ��p���?�;ؿ|tt�;��{��{��={�,��r��^���.�r�o��e��E˯k�h���E4�HT�ڏĀϼ~�[���$,A�Ru�z��J����{L}&�4}�> ��m����K*f�O�$�b@u�$e��PM*�vc��Y�}_�L�}^���<�o$�o���Z@�M���HL`to�ɑ]����W^����;���}�;�IF�_J��+Bv�8|������������3��������p���|�̸a�Y��nm|Տ^�"����/�>@�M�0�yx�y�m�t!ؘ$%F�6x-wi�i�:�e��͝�:��LZ����CJ~_b҃X�! ��oW�����5�����<4F�{�ZG�X��=R�׸$�N����]Z�(������[��f�}�Y�9����;�m	�ː�m�lQ������s�̙�}��W�Ϸ�z�?����OL��%p��o~�w>���<�7�������[{{{ûw���0ވB
jOa�*�!p�8��j���Qbw��������$!�9O�����.䵙SL/#�"c�O#�Y���N��(̤�$Z�Jbj�p�/\1#)F>8�퓪4c��������i�؂�����'�=��=߼O��4�|�.�k�}�w_t�p�u>��'�2L J��!�%0��iꍍ��3gN��W�^�?������~��{Y�i�N�B�q�O�|�'kk�������粚�Y��۷?���fuuD���l��Q�A1 �k�H<^�.f9U$M��������dB"�]��֯�{��^�6C�����X���B?�捫��j灡E��S��A�i@z�滫i�R�T�[֬TJ��}�UR�Ʊۿ�'��ʫ;�6��S=���_��}|)�<O��%�>�O��"�3�P��x�Im7G�����.����L��7�x��}��G	�|�(���ٗ������ߞ8������O���cmmum2�d�~z���ɬb��wA�'��X�݅�]t��������B�����^���1�.�]�u�o����E�җ%b�����}
�1�'�I�ZD�� !
��fˬ@�=f!��Y�C��`�C�=Qi�]���j��p�������zm�~��E�i�VXi`"����V%�=#I :*�)�[0��=�����^z�?�����?:w��?��o�ƾI���N���$(�O�8�Ǘ/_������_]�WeY�ڥ%���ş��<A��nl���?�{�1�.X���_lCyC��dt�pY5���m��i�#`�z���l?��4�},�O�kd<i���wc�j�ETI��/�3K0>فk	�/}�S??>PkUùm��Dۊ��.�\��$�]�|a��~D�@�+�>�μ>i
=�z��s�p��7�P�DӅmb,�С��AQ�F���}�}���~������ǿ�������0����N��� ʓ���?��~��/\�7?�����ѓW삳�8:Xd�({>�b8,���T�{��?�[?��X��UE��E<V��;����k^���N?�̻�HD�EU.��tǰ�[@�Q�*$�<k��7؍�]�� ��ԇ �ʓCC�0V���m1��}�Qj��=�_N�`��:#��� ���[��;#c���}�1�5b0ZP2*WWG[kk�������;��6���\�rh�IR�|�)���09=�]@~��_���v��G����������&��(D���
��}��n�o�)�C��1�Юq@��m�����y�o�qhP	�?!y�B�՟+N@1���Vb��@Ř�E��֕����пfQ�'�30�k��.�`�R5�Lِ�}�^-,I���7�}�o?�_��)9w
k60P��Ff�T[ԯ�~���͍���6�~z�ԩ���+?>y��7�|���˗L�D&��Dv���Į���G?�?g��t饿�����/ww�^��+vO��.v(�A�F�e��ԧ��1�E���]���ג]i���t��� ��Y7Lc�n?�7W�Y$k�Y���	2,��ǈ�_}��ʦ�ĸ�\�
gY&�5���
�-���Y59�a������~�2g�m�<���w��iC��n���onS��9�7k��v���sw��uۖL�6F���-�]Znw;M�3���i2��	��݉ ��Hۥ|�o�z�M�θ&ٹ+(M�ֵ��I��qI�ݳ`�.�SS������A=�]�k�kΜ>sk}c��WWW�KY�����������_~�ȶ3�q5��I""�0@.�c������͛�����3���;������흭W�#����0��r
�IV���������B(�ȠV�,��u�7Ԓ�4]@ e8*ݢ�2M�IW��q�6C~�<v��[����ծ}`�I�Zh�u���y�_�RQw�Ty�/Y&�)�9x�kK��u�uʲ��S2a<�����J���gY�ڂ��j'+��=�\V����S�iЌ��i��&k�	�f� i�� ��X��hۆ:��Tn��͜�#̈��^�R��,�l?*|�/��W��Vd����1B����rJk�>F����t���7�k�dj?W�+5�\�-�:��E��ȖE��.l]��I���p۱�T����~dTTy%���r�W�A^Z b� e�;��p�7���Q����p��6�>q���'On��99+++ۿ������I�Nu(co�����_���������p����/���5�ejW&��Y��oڕ|e<��p��o��ͫ��UK\��?a��o]eӲ"j��ղ�nw�M�ڪ��n�-1i��j����dЇ �03��1��������iK��ql}|'F�K�S��+�������g���P����QVeM�~���K}��Zc*����\���+�2��VĘ0���r��v���G	�Y�$����J�5s�#5Wg?��UI^�����V����GE��Ӛwi�~5���v�%�%`[���ǯ�ۼh`QK=�/���i35���;�ep���1��R�0�%PBiل���>{�W�Ƣ(�sW�gsd�|�ퟎ���22����/���c���T�'ˆ5��oi�;��~�VPŌFr?'Ռ|���W����ǹkGe�Ԯ�S�.�:u�~��`Obo���$�<J�$�9�����}����ӧOo��q�ƙ���+[ۻ���ɩ����`Z�����(�bX�����v�U�`}�^^Z@b��Ns�����)>��"Y؋��t��]��w�N,��8PUM��auR,���ӂZ�]���eLB$Ms��0âE��%�r��]y�E��y�8��Cp�Օr!�iqo�8�����m4�=lY�4���Y[��=۩����.���J������<�<H��c��~n�N��'F�ƥIƥ�A�C޵���6MB���Tl�����&}nmmQ��#0�y����H���im���}н{�p���p�B}��m�~���y�w��U�9Sߵk�(�O~���;�����y��w}�ZG����?������D���8I�9�+�G?q�?ܽk�GG7-�z�2���|�2�</��|?�77i1$���3Vذ{��Vf?���.Æ�!��d��:3d080.x�SY��,S����Ւ�ϟ?_߿�� 3B�\�_�tI�Ƚ0���E~^�2J�'Q��s��y�N��B7v� �D�%J��R'�%J�(Q�g�8I�(Q�D�=S��I�D�%J�虢N%J�(Q�D�%p�(Q�D�%z�(��D�%J�(�3E	�$J�(Q�D��)J�$Q�D�%J�LQ'�%J�(Q�g�8I�(Q�D�=S��I�D�%J�虢N%J�(Q�D�%p�(Q�D�%z�(��D�%J�(�3E	�$J�(Q�D��)J�$Q�D�%J�LQ'�%J�(Q�g�8I�(Q�D�=S��I�D�%J�虢N%J�(Q�D�%p�(Q�D�%z�(��D�%J�(�3E	�$J�(Q�D��)J�$Q�D�%J�LQ'�%J�(Q�g�8I�(Q�D�=S��I�D�%J�虢N%J�(Q�D�%p�(Q�D�%z�(��D�%J�(�3E	�$J�(Q�D��)J�$Q�D�%J�LQ'�%J�(Q�g�8I�(Q�D�=S��I�D�%J�虢��������    IEND�B`�PK
     uK\QQΒ�!  �!  /   images/5441ee9b-7343-4a92-92bb-e3ea11bfaf7c.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  !�IDATx��}k�e�Y�Wuν��ow�L��<�xƎ'	�^-!���GdЂI�+�f�(Y�?P��E�R	"-Z���*+�!�'1���`ǌ�cϣ{�}���T�����ι����H��|vϽ��:u�|�GU�n�\�m���&Ȝ�m���&Ȝ�-!��?���YXY]���8p z�.�1`�X0Y��<����xl���7#��y�@�zn�=�9lo
��~m�}{�{��节�a�7�ۚx>��O��(�_��ѥ����Uv������}�k� �����z��/>��?���������z�Oۢ@�%[�x�)��Gv��7^1Et�$ Q��$�D��%����-�1���F�ق�a��c�I��_|Cl� ���y�8���r��������/��/_|���'�x��?��/���V	�;��Yx����忆����>��_���}��>}�=��c	�Dcg����/��=3������삹�@g-�� ����^�#t��W8�%4�����c[�C�lnnn=�ȇ�4�ǥK������<���������RU����ϾG���s��=�| y^~�"%�*�"�H aw�qP	A�xR=�9U/A�Ļ2�qD�h{����5چo�֘�(u�(IhL���g��v666~����q�������o����'�&�F�O}�7����cp���#_��7~owot`��L�	�?�����h%���ɐ����N�IJ��D�����*HNt�|O�MP�C�Q�+c3,�E�H~js�����'���?����UhZ#ț��V�ۿ�[2x?3���O�<��K��}3<4q�p��_�ܗ�0�qo���4�H:
�=�pVGqb�#mK` ��T��׎7�Y[[����ھ�����μ����V��A^�x:������]8z�z�2݂��R�H�涠��$�u&Q(�F+�����s�17�_�D z�C(�;��e��g��A��A��}�v�:qв�����PCP��[�$N׈K|,����X�3v�]���FT]�P_bH�y?%��+� U>�0SUUx&�����'u�Z#y.���c������S�k�t��&��Qv��+���U��D"�����WWDHR���M`bJ$����y�I�|�/SW��HR�v���ԑ��L��V�U�4�`�s������LF=���	 G�5 �뚐m�{����H��;��4$!t��}���D����/`�xga���I��LT{*!A���i��ͬ�|-Т�[�lW�.w�區�j��e��2ן,�@���`�~9�%;��7<��k�]�������=D�U8�����A�k� �&n�Uب�:�܃)2��jsR�RWs��6ѐ]lZ#���-� �)��~��vdD�H~�&c�t�?�:
֙��"��X$j�2zZWPu���i�r>����%���7`�D�ЇAU����0�}�m�(�{]{��$�"g���"����=������!9�X=t��vp�"�^��~�P��'��[�Q
��-#��,/TG�C顎;���_�Q-����8��;��k��R#��\��$rՖ�@��b�$�F��A�/ؘ7��=��;�����E�K���]k\4Ҏ��e�V���H���v�|�R�U���� R�4�&�9��ev�)59Q1�����&���/�i�W+�8�:��v`�-#x�au��0Br�Fό�����N���%E���$�v�ze�M��;�ɵ����� r�ͨ���m@�F}�H������\M�y�p�]�	m�^�Ȓc0��-���y?�blh�_H��q@�� H@�fu� Je����ώ�j���-A2	p�W��c�u[r�s���xxqa6Ο���X[_�}H�'�X}��!�@��6�Ƥ�"��:�/�yN�3pt����!�_�<dڵ��nr�qa{����.����q|=/�y�3tF��a��8(+����N	��dH��qBS6�~��gCꝋ`�m�'�r�>{��U�_'@��к��Bk���Z����$!�1� ����bt9��Z!�&��� �<��S�{��^��(�!�� �cug�@`s#Ѹ7��jVnKk�s+!l�eൄ�rp,�������K�ِ��:EM�)g:N��L�P��@?6���ג�Pg��SbB�/1�*�9��J|ytA�PwsPIMU	#��}T���`�2��HL�ת���<H	��q\�!yFܔ������
�d4E��
�m��1=��u�\�`ψ��	I� ��@�����[Gn��yb�\(!LMI�P
�Y*��-z|b3���������V
�yZ�2�U�W�lC^σjCg�Hщ�RS]Ff��\���Z�&�(U���yi�F>>W���_	�b{1�|ك8�f^���l���N #`-#�qę�����1R0 9!��S ��$�EZpkZ#�x4f G��5�֓s�A�\c9�g�f*�2.M�S�#���;���>(!�����R�!�����(��в�j� �Թ������E?�������n�#�)B6�u���L΋���\d�:�Ϫ��ī�q<̯��34Y�T7p�߳�Hp�O�p��7������ψ�.��R%8>ڥ|L9��>]�;�}f��TeEU6S�������t��#���R`a�U՘��:WK����+�:_̅�P���Ej(sO���K�q�r����S/�,ʐ��t̖���sjD�$O�u����=-��%� N�S$�8��5�Q�O��,DC���=Wi��������:*u[���\��s\>���H9����U"�h@⇔�*X�*����E$��E��
Qr�ܰg���L�t�s*!�^�?�+�q��3$A��8�
mD�D�׼��$L�թE J,h-<���n2R*�ܮ�:Ir_'��G(]
�>2�U���M�I�XK�l�	ړ[D��M����@��3r��C�Nv�����V)�7b�)�r�L�x	�jl�L��~=\�B�:��_^�10��|"�@S�&}pNb>�@{���e?�����i�spa\5����#��S�m�!j.;t�l+X4��$�߃���
��%�#o#29��u��+7�$�u�45��h� ]��dv �#'J
Ĳ>�K�	�G�r�%���&@�/��+ꪤ놰�z�d�pe�R�H*Io�m��c�f����4I#w�o�h�mԹZ]#��8�ުQ��̃Te�Ȗ3	)���
7��>�A\BRs�Pq9>3�l]4^���3g�\9��3�к��xY1}zlFo2)Rې�7A����7�*�5GP�ta�w�%��2:C��wH���������3K-AB�����>ڄ	B^�z�?�%�L�Z�3�'ȍ(yh;�ߚ���.&���o�䭪����PA����M�zU3���C�`ww��;p�С@��1�����I�z [(��A�m�.��;�lJ΁:�9\OG|"r!����0�2b��X�/�qE�m�1�� Yx#�L�����+{�-�ի/�}��._��n	�F��X"�,ڝ]9T�@� �6����v}��[�i��#�b�ѥ�GrRL��9ŕ�4�Pv���>/�9}�4��̸�Mho��uuC�lg�h��ϑ]�M�Qp���}<����.������Zx��~��'Q*��u��j��S;t|ow�k�:��B�A��,ez�D�el�� �^+}&du�>��q@X	j8X,�n��^���	ڌ��^�G��{��"i��٣�riM�K�z����x���J��{R���<G��V����y���lJ��Y��y����{pje�y�(���]�����<�1���щ�M��s�5a���D;u��Y�A-$�h�+P��lC���.R媨���3�¹�M2Υ�n2�/]��oy�F �7��+���@>�\"k��?F�7�rj�p��L&���A(ub�J 袘<��&�s%U>��i�ee&�����Q��a{g&�4Io�N	����z甁S�H�pŐ�g&�{�%��S����[ԙ: �c��-F�e��f�n��{�<f�4�������������KK�Q�>H/[�TS���X^���~΀�6�c��i�V^��ؔg�L����f���;=C�f�!�o.+�'��S�>ا��W���X9�r#�0'dchZ����^Ҵ|,q�r�e5&dH��� �X��y���5�\��ؾ�¬s��q�[���G�~I��<������s&�5����SNM�0�z�/�iV%s��j�����]=�$�Mh/R�Y�1�#�/�Ƶ�~]zT���2��������bS���
F鲃@\?C���"4	��m��4�����Y'E�)d{�R�4���:H��.��XV#��:1�A=���� N�GW�n���*�=:AnJ���ǯu���#�no߀���0^^Y��Ḓ�%�tmAd�)�R�K�ߴS���l���	�Z����ͽ��x�0��=��=��s���Ƣ�2ij��K6�Y�i��r��ܼY�}����?>�Iex�K�k�VUV��)�5��WY��3jE9;$%a�\T��0���ʎaP�a�Z���7�0�������<ߣ��@�۝�?q#���-�r���Ҝ(���������aM�|����{�N�O�q(��vlz��Ц��}��$��Q_q?Y	���Ḅ94c����s�t:]{#zE��
O��ǉg��D�I���0�Eꍼ�k[;Pv:A��8RwU�9Iۆ���H�m�O�_&�Q��rc�#�Z_:������C���2�e����!\�2�<�;2�#ʧŭ��=WWW��t{ٹ�Y3뮫��p��9�
ظv^��"\�r�u0��D���~�_-��e	���Z&W�Dl;�����u>����]�hzC�6-u��3al={�$}��+������l�a�6έ)�����eL:���7�liV)�^'�,�L�o���>ƨ禥X -������n�(z�@L���}*�(� �)e/w�s�����^�Nj�e����jC4X*�����{}��"y�8�v��,��߃Ԙˊ6dN	�E���5����8_6�L�I�x��&��M�5wj¿���g�Y��Y�`�ye��%�b���.��<�IDj�(40�q��)4�N~�Hܒ����`V�`V�1�G���upq}��s?b N���mU����I�ՐۍY�=�ڕ~�����#̷�t����!�Tg��&̒�iN�XD7Hi�!�>k��AMo�c:�PUY�+!Ԩ;V^p�ѦL����H9��yS�bݩ��,�eǸ��砒��6K�5�_�CmJ]�ږ�VS'B��mrW# �|P=��x��=>4�Д��a�Q��^�z��e�������{͒����YS�ͭ�"�� ����	t!��
F�+��6�i;���A'�4�i��r}8f��.�>��˴,J�2�ª݃�!�>FEӻV�����q���Rդ�c��&!c�l��8�`ڃ�!�E��AO��m^��p�݄�U�](&c�;H�����^s/��t`u�E�8�d=HC�����z�Ϧ:�^7�oZ'�mEK��8��L���ke�N��j�CA6�t��%\�,3�W(���wT�sv�k�&PZ`m�z9��T�L�_��t�#��4�M���p�<�F@�T�Ӄ͞+�5a��>p�F����Y���X�ظ�UKpg�l�8X���p٭��-��^v��ՄW]����W�lu��ݷͫ�[@��e,6LR.���6&M���ɖ�����(S�
��K8�3qHM-N����u0t��k)-�)yr^��k�i�f�v/ef��Ju6 �ˡ�����;�Z�U��ܑ�C��|��^��`�A��Z���W������X�S.V��B[,����x���&Diǰ膼0���Ү״�jl{��3[3;hk�е��5.$E�A�����ҿsZ�"0��8��������%�=�%�q]q]IRl#W�	s�`Q5����ó�(,�5kv�X�cޔH��j����X�أ7' 1I�^�a���tq�]�2�p��s�8�Na9�~�Aw+���Z���҆u��2�d-���3;��a��+���`�ǈH��s�Б�+� �{�O�=$��d	���}+fG�ux�Z�M��U��>�p��d�/�����D�����F0�Ncؔ\�v�A�2���jZ�!��t�>^(Ivd14�Kz`�W�a��lu',�!�$Bҥ	*$D��Z� 9
�J���MF�:��(/�Ax����)����% 틼����vo�_�j�Dr��������RI�>�}r4�� s�e�l�l��X�O�'	]���y�`ԑ�����Wvf�^�}�����X/c X�T,��.��*��2It{����"L�S���Wv�ybF!Uù.��&f���N^	B�"��,�6P&�� ��8{Ad���MH�Xު���>xr�a��������g�,4-����q���M��`�j���u�}[�m;�*A\���}�嗯<=�޷7܃�h���&1�k5R�5l��k�����<�eg{;�I��_��/ý]֟3�\ud�}N�4�N ҟJ��ZY�����_����/�=��;��%ȯ�گ��y�?~���r�;<Ð��g�����ً�s���t�]���Ӏ677y�/#�CB��N�$dN'!H�JI���ҷ����H�������>��O<�m���Y'����=�W҈��~��v��'���Ɔ	�)Zo�+��T��Zˉ'j�P�H�������TC�r�,�$�X��Gt��؄�|��w��-4��eqS�J��ҁ��Lw�!дCsL��5��xm�Z<4��)�ץ��u����ݝJ�����˗w�J������\߶�]�n=��B�	�����ʔ����B_iw:��B$a�v(K���B�>٬��� ��*�#�ړ�R�$MIҝ�c4�;"�~��Zh� ��7�A)�@C'�(��fZ��y1*�ZU�B���`��gMӧ�6�D��}�c��d�P���J��m����4��+r[%H��==���'>NZ�C��^�������8~�fQQ�/_��h���dn�kn޼ׯo���ð�_a)�)��?�]X__��x����O��'cZ���籏-~I��b�*��a�(ӕLˇ��Daہ�H�����q$[@�<����J�������
����~�Cb\�x��Y��-o����m<�����C7���⽻�_�s�͜���>���g�=����!���7��{���kx�g���~������5e��sH��$Q.���hYe��-�b(�M�����h���ë́|r-I�ɲ�]~-�' �����؅�H��9�!d�<�S&^��hpX��n1_���q�1:i;���+++l�ڄV	r����0���gu�~���As�I��3��Ie;z#|}m9��P=]�7��{i;,��������}��{&�	���o�k��ZZZ��p�oK,�>}oNC/���1�a��y�O�����f��ṅ��SǏ���w�Da��r�
>�i����o|��"��=/��w��4|�P�����YI�	U��w��m��'��~���h�Ջz%��������8!^���c'�uw�rXFritO[sD�?��?��o�,��O�,��}��5�J�w���p�����?��U��G������>��6͍gdն��k��e_�&c�j���W�TݞC�H3LԅMAe=���@��L4aJ�T���^i��yuu��_��_h���ď����T_��?������?���ϩ�'|kk���q�@������^7��(%�d�i��'���KrYY8wb�9�|��G"��d���	]�_nC��A���ʉYH�3^V���]����Ͳc�<q��g/\�x�g��G}چ�TD�O�3����|�����?�?������T-�
T/���,>+��Uƚ
3�b�7�*�#�0���n:�I��]��r};��T�H�,�e���G�*j\c��a`�{�.,.-�~��X��e��G?���C�VV�p��ux�G��n}��bȟ�N��^�'?�)�x��y4��E�W!�E��*�#.���\��z����;8-,k��s���ä��Q�S��H���=6���#�.�B[7�O�6��~6�]��|�#�,��Z'�������m���-#�mxup� s�	2gp� s�%��bi�,    IEND�B`�PK
     uK\J�-E�I �I /   images/10aa979f-dd42-43c7-9c2f-b8fbfcd42f21.png�PNG

   IHDR  �  j   ):n�   	pHYs  �  ��+  ��IDATx��Y�%�u�7��̬���"���E�H���$��1`@h-2`k�@� �~P�x`x���q�z0@c�a�0F{<�/�ղ,�2%єHQ܋Ud�U�b�Y�{޹'�N*����8q���QW�y+n|q��;�s�o.1������������֒���dff&�E��h�����Hz�N�}�C�>�
y&��|b�r���=�3!�����3U����T����U��}���.T~,$�y �ȳ3`�M��y��^h��P�O}?�y��-�m�	�������L��Ѻ?@�1�L�z�恷�й$���Wa=��3�|B�ڟ{�Q���n��� ���ź\��yk[�8�ģM��8�����$My6�}aa!y�ᇿ��/|��d��K��������g���\�t)9z�h�R��p�� =�:�A���,A�J^]�!��~�11*!F&��C%֓�i^@!��,Ԉ��ɀ��̶�b9Π�mW��<���g�K��vra�m�gF�2k��s��"Ș��'V�c���p4��=^[���^��`�c��]�밃�dXN��D��������D|N�:�|��_��N�<��'�|��dJ��)���'._���o�����{ɱcǒ���t W*r����:�X?7�x�|n�X�W�5d��*\x�id�� �~���ь�\�z`��a�'ru�\��u���h�\��X�XQ}��UL�Qv���B	S�a9�tad�i-�0#x-F车o�p��G'Kq�z�d�3k<�;�X;?h�b�w�}T0���Hn޼�����'>�G���]�Y�.�.]����JZE(�L�5�Q޷�\������0�������Z��s1#�X]k!52�� ,�R�E�؞ږ4BУ1�w�-�<��1���ւ�0l�x���a�P��$Qg�g��<:n��K�t�و�N��>ل`�1���՟#�p�����̭���F?����f�/��D��O��g��~r���o��o����)!3G|�;���T�w�}��~���D�I%\^^N�ʫjn��}�*uQ&�\��W���	r��
f��=s!�'��-m��*���fԔe��8���:�U1�gIY�u�f�>5�K_�f���)���s�hT0���E62�s��`��q]����cz��i�S޷X�na-��uM�U,���5�ֲ���H'?%�G��^{M��?X]]���>���\\\|��_�b��4��	������_��_��ϟO.^���[&��R	%�L~nmm��6��v�}�Tz��x4�yR��]����h�^`�i�`f�C��F�5�!װ�4u*���΄����.�~��i3A5̾���#�iA��*�#}���i��/�<��1�y>+s^���G�J���n���~}�k�0�s&��1�)o��6���������Iu4dF{W�K�'"��D�*�o�N�_��'��/~塇��G>�dee���������̜p���/?��sɫ��z��/��ȑ#�K��R!u���-D�j��m´?�@��,�C���a4C�y���ԧ��Et��� mA�����7���df[��Y��YXo!c	���<�� ,����yK�8+΂U N֑Eȼ���|����}>��i�,A��멓o_�$�AE��:@L;})�~�:�&Ə��;���e�'E����L�L���d�~�֭�̙3�k^�}(y��~tYf�d�*����Ǔ�~8�da�[0�"A�Hz���D��C'
,�Y�^�X�3��&�z��<S��*�3��ګ�ʰܒ���쬍�,X���E��f��^7�����8]���d�ǂ��A�^*(U݋ц��s�X���A����}��Zb��L�`�W���,wΙ��V�k��ޱ�kl�`��%�v!d�3��%�l}}]~_NzLfN8y���������/�tb��J-�NW����׎�i����9ad�QX[����Jɺ{��G3V��4M�}�{����d���%h]�8b���z������@u�K�}���'o�� g��i\�vA�8s,F�(�NC�-�s�9btA�|�u�i����0T��e��;�}��S�8f{��<@�G����3����o�56���"ǽ�)�%LGu����ւ=zl��>�괟�MG���=�B�cB0s�������2u�v�!��^��,�y4�0�Րk�,��{{�}�!"@"�^:�E���g��`���"˲�1b��x��&�gE��`�F�V��b�,�i���Vڀ����!�����z�r�`k�t�)��E��{u��,=�����c�����4��1�Vݏm�q��t�h"�K˛8������9`�g�`-�X����}�y�u���R0�vz�׻�y� �5޺u��_|�ӿ����j�CB0�3g�,���<���y���ן|������7�L�ь���1Z��"��X����Kc&s,z����<`�1K,bzo��U0C��qad���ѥ�w+̈́���45x�x��O��c�XG���Ɖ(�@�kl4�aO�1s�P�P�ΤBٸ�=f(�ΈL�����)�yt��S�4�m�[;f����Vtof�bbi��H=���=:xT��ߡ��׾�5?/�򟓨�7�x#y��lss��-..^�w�S��ԍ�'�`�/���'~���ϯ���?^YYIVWW����'��N��3�5�3�y0��el�Z���!s�Ș�t����+Q�6ILϯ*�N�'͈��֕�G��#M����Ƭ�~��a�=
�y��ra
 ������`�r�aF7��!�+�<'������x�E17̊�����J�	s�F� 6��!���{�`m��s}����L,�ڏ5?ʮc����1���Ж}>z/���L�]��?��w	z���7���o�8q"y����r�ʿ�җ����Y�;w��7���'7n�H'PY&?��A��	��;�ႍ���s��UWPo-t�����':����E�;�}"��S@���A�FSg��Qa���a��m7�.���A��ֳ�k��x����IkuǈI�]]���x#��̶�D�K}��Sr1�U�2����u>����4��L����U����P��L�Fd�.σ<S(���0@leu�]c�r��L�QL�#����˸t%�666��g�&�/_N�9��T�>��gF���!���ye7o�L�_�������W�������b���Y9���tK���I<b�e�ׅBf���vW�0�I�s�-�%�7wU� �3���m�c������`�QL�Do��D�7�)#�u���>C�r��L��i4Wf�Z��N���ZW��f$�WXy5�n�O��h^"�1��-)�
/���3��ˬ� ];z��U�]�m!{��پ���>��#,{K�3�&��xci�C��>���ؼ��W�����t����ߏ;��W�^Mߓ9���v���?������>���%�	��VWW?q�Ν��� %U�Ի���2]'�u�A���u��~��	(*,2ϥ`M����sd���8(x�/��]&H�[e%�<�"��L����v�o�nz���|l�f��-`����F����G���z�x���e}v����C�zWg��zX�0�0̎�@ҫzv��H����ӂ5�H&ޢ�����eNk�e,�~D0c=2^���X;�y�>Ba�%��؍�:�j��#`1@#��z�5�s���=z𾌽yv���&= ��y��'��ɓ'�
&I�n�(Qf�������a�ް�>�X�'�v�轘^3^ˆk�`=�ޖ�c��,BX^Q}���y���3�Њn#d9Ob.l�����ѷX��6<f��S������XG�e]h�CQ�7�KMa�шΜO�,T�E`ΩY�s����u^!�^o�Ҵ�O�=��PV�Z���o�B�b:�W�:�"�+b�9�1m;L�?{��SR�^����|jg�v�����5>���:`aaa��8�.�UB��hdyf"xT���,X�X��7��tk#Ƞ���5�E�&�â��({��s���� ��~}���	fY��-�B0�	{�=�i_汿��t-[���xf��+0�`6��(�|��5 �K�)�������j�<�vgak�?s~g�vDi�]�=��-�;��	�k<�(б�DU Q�끇�l�\[�$�3
"��^ǒ�Y�s�=��CJ�Uy�h����g^N���Ho�i�ݬ�}Yu��P�\cm��Z/
,PX���=�M�#�AO�Po�7�&�]�~�{��Sf�$-�u�տzl/Lc+=��Z����F�4����g��ֆ�|z����~E��aX'=����^��,�4`G�1�Y}u��X�s"`��e� 2��<CȫɃ�V�e�'m��e���P�?SH��vH`���[�8ǥ��d�|��#[��el��C��p�^�=IK�����4�L����w�l>�!�u���KeY__?hࢲ�{R����������^ō�z�1=O��K_�d�.hg.~Yx�OtB���`9U2�Z��%x��[,�Ii�d�-��+��6�o!�vc�u=`��z��LG�F�&b|���g�2�X,k���ڲ�ڑ˫�X�`6��QU�Sf�u�R�`9'�0}�<k���0.�Iہ~����3�兮���U�H�q�1��~E׌�����p���+Rƪs�`)"��>Jg!�!�u��[�y뭷��gϦK��6���C��݋�0��Q��o�:�v+�.zH�%mx�L���US�#�X�D	������X?Ҏ�gB�}x���4�ҳ�w̳@�30�aE�y�nL����xTw�ǖ������q�5�!0a�~�(:�l��2�Q(��G���ޯ�.ě�Ӣ{U��Ν�t�p�4~��Mƴ6E3D�c�G��EM����*BF�`��A��~m�y��=֘�l��������dn߾����~�x&g��-����`����-��7o�L��"���[2JE�l���,á�53`��ͬ�¤cay�!޷l��
�S	������	��`��R4C�շX�73�5��Bp�����:\jx��o0�S�nbM<3'���1����!�y �Lu��ha�7�T]�L��̠n�u~D�&s�g�^Ym��F�[;n�`{}3�c�b���:���Y�u�5�x܆(:�8n�ֻX�Z?ӡ�����	e�-��޲�����;�7R.�ԕ6�x�SZ��ڱ����g>�6@ۺn�x7�L��J_XX����:`TI�x衇����t� ���F&���VXO(�6a���xF;Y�ֽ������g�GA�YX�9�ݬ{f{azk������lkVz�t!��u��U�1�<�9�����@���|�sdo�Y�>Ð��nh��չF�`Ea�-�y3f2���u��tˬ�{Y�$*�����B��x��ud����7�"a4���7�����{�T��˧��m-c�<Om�Ϧ�g8:bo�3�$?D����HN�8�|��O>�����`�+RQN�>�F�---���+k���4Y{��&�}S,�]xky���]Y�g��2��:\���7�l�����g{{��gV=`m��^��M4�|�"���핉kVX;������~?k��U쭎�A�"Ȥ�b\c��G�c�)L�u�u�(}�	��`݆ Qt�q�c:�`f+��	E��XG(0�X�'C��?sY>h�ϳ��MĢ�4۬�m	EzKPB���!���""��!�w	����Q�Y\__OVVV�
���v�I���l��ě��.�$t1ٵ���6�	f�k�X��,�ňQK�aN�<�?(�>�%,2#=��i��-����Wq���b����KYdM�/�"$x4B2�:,A�����쵇^7.��r�W��ff��ǵs,fm�׵hQe �s�2�D�m�m�l3��3�	g̾,�P�Ae�[~.Z�Wu�ת>�-'�63�y&��Y���8���z�=�D�I�����r�B0�Q%9}����i��U39��ɚz����h�f��5�`�Z�#x�ض�6@����3t{@d��M��3n0�	�מ��Ƚ<�,3k��u�-|[]��r,��sT0kk�D�}�2쮱���f,��e=g]��5.����0Xu�ٟ�`�y�kP�=�Q���8C��؏�g]�H�4�Ǻ�g�)���u�
Xe�g�_�~�q�bP%Nz�<�.5L;[0�J�e��3�f�~D0���y�=:����sB0�QE�W��nܸ�
fR�T$�C�* ��@��F ©�<b@�3��b��UTc�gQ�
������kD�ǅ&�GC�08�T^�0o��L��z��<�^�}��6<F�����!�s��`k��mfa�Y�y�k��e���8��3�p�t~�v�kncY~^��]��h'�X��y~MA��:y���E7Io\:L�R�<
��w(�"lR_���>�e����O�.�/�s�ۊ��%�(G�=xIë�``�̳c,�f{fZ{=v���e�!
��<�uz�O��s��F7T]��c�
f��C�5�>�hz���M�w*:6�"�<z��dk��)��F�^U0�I��y��"�A�}�e��x,�R�і�m��h�I�3Rd0��:mR��T���XN�L��u1�Ε�ǥWt=:?G��,�q�,�q�4�}P�:���̋|��ڱ�=d�W���M?Ì�*�tb�Ek���3��u�6Dê1��Ҷ4�L�c�C�[2�����y�ǒ�Ǐ��E��h,�I�b�P�/s�:��1 W�:I�)�x��`�ub��i�+?��jfO����-0aX����2gA빷��Nϛ�3����r��e���j�Hߒ�~eFV斌�󡙰�|\tG�:�j{h�,Gf[G�i먓]�:<�0�W]�gY�;�9gz]eu*��l�jWbJ>�!d�}�*�g��٩��Lj�T�b9�E@�y��n�qi��o�sLϸ�@a��h�Hz�3Bv�q	趢u��.R�^��ɳ�K����c}}���`�ǎ�p��T�0"�I#�s�΁�6�W4��gN�V�aN�-��+�I���I�Nά�����5L����b.~��t]��޷,X�3�IY��ύL�%=F�A�6,#�`-�X��(j��ǳul-rY߫i}*Z|�md�6�I�2k#�Ú�L,�y0K�)�W+�|Ѷ�6�2�C�Ek��H�G0�����ѹ9�$��V_��qQ���������k]߶X��e	fhzE�LM�	�sf���,��qQٿe�C�3U9�T=���R��ʊg$t�Ν�&= �XXXXYZZJ+���H//�.�4p�!L��ϰ��z��>�m�,X/��
�P�\Zz�Y�"3�{
��%L#����\^^��#й���b�5�� �K�s``-��8�X��Z��ǈ6k���L�Ne3������*�EXs����͉�w�3i/bW`x�3e-:�:��(���Q�45���Ω-3tMϊ�g�/�㬥�;����6iZ�w������q9�A���$�"�k�m��	�ot�E#̪�W�w}��s����{4�YKz@f0�\�]�d�<Z�E�d��Q�	�x�N=�u��5�?�^�|bM���3@۞u=@�n{L��fx��e.�Y�4ϑ:�>�s!�������iţx�1�<>���_��������4�|R���3u�7S0cE����:U��^E�q��o�Ї��z�컡m�����)�<,a��I�/d��o�u��}����O�-���(EϞOK�)?f�M��l+���U��!�u����i	C\]]��`&�eu&9�<�z^Uy�:Ok��əe[`z�Z��(��i�e��L��9a� lT,=ڙ�}tqϊ"dF���m�Y~������0ϸ�8�{:�nb8gE�C@����w�ԑ<`�����s4����]@���"UiMb\�v�?�&�p�W���tRV�����g�v@��9�c=�.&�����6��θ.0�"�0�Y�˱��1�(�ѵk���{e�$Z����gk{�9���cI���^��k/^Lnݺ���������<<�5)C,�L�������k�}��>úo�ƣ0l-0�0F�u��W̳UX0�$��|�2�"}5s�[gA^��,&�F3�!��P�0��q.��VJE�c�)kOt��c���H�ͤ�����9�`���V�(�fl�n��rm�٠�P�l��`�X��@�.�}�k'q����b;�q}�by��
3UX�k�e!/R9H N�1�(�:"�����<�Ȋ�̘7�x�ĕ+W>���&ׯ_?�Dy��ˬ�5B�bh�q���nH�L���4��`N�2�+�2A��:�a�5���Y{�`.��2F����gB�5�z�pE@� ��N��H[@��E`��6SS,��xc-D��C��D3���vZH>"i�XU Q(,�=ܣ�F[[��<��<Fհ�Z�I����R�d�@U�X�)�Z۷�<@�W4/=��{�y�tL+�c�~�Izm��Ƚ��l��&���s�4Z�9���?�FmU�T@������� /�vcc#�[�"_XX���̌Y__��֭[��z�jr�ڵtQ"w{{�@}e�LXޛ!��:���hoL_t�*P�"k��ퟁGc�YS�}�gB�(C`>��u��(���A��֋{��#���]x	z�;Y�DJ&ˮ�B	�|�K�{S��5�fҦ���y���iе^1�o��C�U�\Ɖ)���`�traa���u�-�"��t�^d���PXN��Qo��_�����!|U�7N�`ϑ��Aٳ�sE�3	ޢe댳u�|\]@��qf�k�����HP�
f�
f�����Jz@f�\�x�z�w�K�.%7n�H�a��2�$f�����!�4Tz��Yci�dz�y�i�^ [{JZ�Ok�=s�θ���o2'p̲�h��+}�w=XQ���l{L�lK�u�e|C�п�-ʫ��ÚA[�]fP�c8���A^��>��z_'¬���͑B�8>Z������K-���>%<�Wy�N�Q�Lu�*���Ҧ�B0�__W0��>��M��<λY玡4��ڬw���Ձ�S���3akk+}_��Ο?����`6!?��?�ҥ0�K��{��ǎ{W~>������Μ9�x���'������{.�D(�JtWaMW�l�E��/+=�>,/:�+�c]����>s������6�^�A'׃����N}�\d�?Ƚ��܋�������鄵7���_�bQ0�#=�x��׹+=�0�a��y�z����f8<�v��X<��8ĪS^�a�su�|d	3�X�Y;�h���R^mu����M���fb�V�y��h"�����o��ϟ={vakk�����lnn�:~���_��_11$�	��?��3*�?��1� ��{o2*D���=����������yنqmm��7o>��� �r�JZq���"��o��Z��g,'�}�o���>/����Kn���A�dL<���m�}�\W���␙+ϻ�*�[�}뭩B0ð�_��ź�Y���Sn��<�{jG@��`�a�K����(f&}u��Xϭ�
��H@��e�N��%X��W_M�~��o���[��{�������Q�[����D$[__`cc�A�J�}�v���~��;w������#B0k�s�=�k�>��|���M�"�I�l������#G�L
V
Y^I&g��u"�I��U#Ͳ)��=`�����0�x�kY.w����Հ�«��^��en]W<z2��ek-�2�b#^��G�Qf�����Xc�y���� �Yb��4N�8���f��:�<�r0�s �2F�gU��	�>��W�M��rA�DَQt�7�;�h#��|���O~���-/,,|A�i��,��D~��T3y��G<y���`����O����i��^'�͛7
�@ډiGv�ȑdyy9�8���K���ye8C�S�Ҙ�\D"��(���`ճw�����|8��E$
�\��W��ު��⸷��u�.~�g�xgYtїOs�0��S����:�b��i̬�!������[2N������b��b�t���|4�q}
�ã`&��M��<:I����=�]�!u���-L�d����z2�\�|9�x�bzmV?QDD�ψ`&ל;w�+gΜY~���o'�`�9�L�Q�(�����_�J����nè�	R��|V~G=�<by {�%����=�<����e8��E$3y4k���uA5�������n�ɤ��4�(��q`�/��[�����<��i޺I8�ҴÜ�D=��Y�n��tf�0����A�']ҖZE3�EDCQ��^�9�wyIБ�ME?�ȴ˗/������!�5��7�\|��W��lŨ
l6�P�pBA�H�%�,iZYT)�kE�C�����z�[�N֞�X���X�>H���W���:�x�b��Gz4��k_6��Y{�y�-��QX�	���,��c�uL;���]�z���<�r��\�����$}�ld���E��.�KGnk"j���K@�d�]�q4jʣ���[�F��Q�C^�ҳ�t+��=�3��L���������җ���G�x��W�������o�����b�!L�W������3yɿ��*���WUR��� &
̽�{y���K#:�h�\��e����x���$���Y�W���<`�<
��E$ϭ����JP"��*�i��F����9β�I�5,������I����pȺ��Q��Q���.
��V0�!�C#:����lǬy�\�F���RU0��z��k�����%�����}�O��������Lf5������������'Μ9#�����X��h��O�^�1��*���&��z����x& {�"�MQ��u0�e	f�h�J���}��b�a,9k�z��^dYA�E<f����4R�c��P�����
t�`�i�h~�x�c]n�OD󠯻` xt&�7����֎),��>�6�hu��4�L��C�ϊ ����E��流ܼy3��������+W~��_����O���Df ?����ۿ�����O�ܹs��u�ر�Ф%�,���v :Q����*���fUV��U]���������Ӯl�.��-�<`ۭ=��E��� �}zl֞�L���+��z[<����F,o�a����9L�����p����F���el�W��B����U�w��k}�F��`��X0�s�S��^���k�#W�~�O�Z��[�2�5�U&�r/�;4PHй��%��J�)/��d��ҭO�8��~����g����/�����=��Gyd+i��@^z�o>��s�8�|ZأBI_R���bv[E�Z�"��K�V��DZ�]��[*�m��u�<.
X��.��f�G�l{h{a
%H��CD	梎�G��8����s����(��Å]_�6]�����Y�ʮN>��5tچ���aa��x�o1��s@d�̘}��s��b]7�4�����]��F��)�K�`�UH���=X4�q}/�Lʞ�Izȳ�sNMO�zשּׂ[�D[��ʲ;pݹs'��O�7��wٚ��ի�k����:u�+������#����B0�����_�я~���_�p�}�%Ǐ?�"�I�L,�\�H29�L~f+�V�����!޲�C#��:�Di#��{j~[N>�1����N�X�L�U�č6�.h��^�2�1zF ��y���i�-����2�b<����-�йb[·<>�(j-tY ��x.fd��zǤ�s���w���t�1~@iy�=���(ª�{=���z�EiR��ҷ�����3�]������1��ux�@�F?��	Ev=��`���|���'��f���ӧ��~8���Jߓ�ݺu+y�W�_��_��}�k!�u�ٳg�.q�ڵ� ����������۷o�?E��V�ߥ��(��v+ډ�V6Mֽ���*�"�h��n/Ȥ����W��ݐ�n4��Ү��iz���z��q�p�y���-"D��h�Ϟ�Yt4I�5��sW=z>����rn�����ݴ]�ǲ��6XO�\ʺ[ߋ����:wC�C�c9������τ`�� e�̷u��J�ˀ��:�D`���uR���Pg�9J�H���ra�e���z�Ov)���g�(J�_-A�ݢ�n\&�0�>K�yP���z�d�VT?������Ec��h)��;���"��s�=ɣ�>�|�S�J��L��������=��>��<��	��ʕ+��R�K�-;u�T�}(�Td;F�x��������TݏS���k��"�^�uҬJ]�1@'B(�`mx����(�"D��梎�O� ?.�:��c��u�h)\X���޴Nɿ�=��@Ģ�qv�s��)~W�,����q0�<���UVyΌ�AYL<�y���G1�9�8���X.(���yՅp�:����MkQ���1#=�v���Xu
}nd�
�3�̃Y"��c�G����%����U�
<M����xt0k�Le�{�*!���c����E#�d�>yi ��&�c�=�|���M��nܸ�n�x�������_^�9�Hf]���yB
qii)-,y�{�iAJH��f��^Z�"���Z��S�ʫ�g�s��	=Z�Y��3=�X0���+����Y���3kd���9a��Oo^�B�L�^�>�t!�ģ�3�X��Zu$ϛf���b;����]���S��K�y/La�R0��@�Fd���~�sKPOP�^���g�Chz�k����b��(���sKgKf�Ì�b�:YF1�9�nB�	xX"%��3��z ����~뵸����KA�L�����3�&�g f�é5M�����M����9��N|���O�nQ�A�/G[��"�=��Cɇ?��4��7�H�n޼�F����=��@f �n����D���)a�R`�S�M��	�nèF�w�t?�>.8�X@!0b�}X�/;�L*�1A̼b\���q�k���u�KSc_�2�k�?Ө�\�4쳄h��Lo���E5p0�<� ��i!s�A��_dm�k}�|&�>
��ipAEQK��o�z�u����,�2�[���2�������=0=��1�[T�uzh�渂����b���c5����֑�}�V~2�)KG����ӱ�+EN�M�����)����t,�K�+�]��w�X�{�O��UW� $�b�%���\����Y�����y��âljETTX=tND��u:���"�I��˺A[T��޴.�߭���� P�G��y�9���J�j�{������C?Nhf��MT���zn��]G�kbn*��]��<'�,�c�C����iY;(���1���X0��22��L��l�:��3�Vx�XX��s��;�T�Q��*����{!�����;�X�6�ڱ����Z��R�]�y��9K�.��jS8���U_�;Kg	f���X�1��r%jL�O��tސ}^�>qL4��|N~�gF�?��@f�
�)<)A*����o��:'��n�(V��QC
�2���x�6�[f���M�mmxB�bM�[���P�n��5����3̊��N[`ԗ>��i����g��G��.�3����q��⭾0��hz�k����y����%]̗�ͷ��b�4j{Ų��N��p�4X[��̈Z�h5�(t���[e��HDA��*�9<�f=G�`f�lP�~�oV�S�X�@m�����[�Z�o��U���l��OD�<��#��hRVp���h1ׯ_O�y�T�g=F��k���5�����Q�=����
b���.{ej��j�Q&/�7Y_���X{[p{{��2�EY-T�ޟ��c��K����),Z
*LOI$}k#��f��M��u��Ԉ�T�ey�
E^iM�i�C`
fֆCkA���L��x��}d96v��~�af-�������f���|�Hf��h�����˵��Q[Ӝ4=�n�"��X�he׵�3	���y��3*�1�u�!���uYƓ�KʰJd�+F��G�L�K5�oe�>݂Qґ ��g�&ǎK�b�?.^��0��:��%-�Y�j؟aR8Rp:A�I�P'��Au��R	�@�.��a-�0�%X��̼Nά���,��ӆWɤ顃��'�`��?`�<k���Y��c�T���D�-*����Y�XX?�˜i�A�&n�	����/�9[�,?�h&���7�L�6�[ΩC{���*P�=��տ������3� �\LѰ�^h�={�v�1rk��.D�*��qM"�M�F�v)�:��^E�an�ۅhVtm�o��U�]�|.�o�c��'�R��t�EMgmm-�p�B�$��O��}��ݝ������Q�/��%�������ɇ?��dyy9�t�R����.�i�PÂ�/)�G��]O<�1X��:�5���~�^`=P�0��*<ͼ����ī����z�e��`;oaF�0�C���I_]V�ۚE�)��h�L/(�/��1�$h^��EX�$�}�mƲ-0�i��Dh��sZ�(�M�a�ڢκ�2b8��e��߭�b�tE�E^��l�(Ϫ����W�$�j��%�=$��W^y��'�x��|!�U0�ċRX"vI�<�|��O_RhR�N�<�Z�=k������fڷDc\s�|H�'�]�y>�(�_ �̱����6�u�hY�h{��?��I�9�1�#y��&�y>��iO3m�NR$:��aՃ��i���>Nw_��i)�(�"�����<B���TT$��Q�{��r�=���K�o�&��d�FPj뻄`V����D�IA�~���G�'�|2��'?�n�(��K/l�A��<O˒.�C�%��h�.��z����=ɽB8k�{�
�m�<�iM������B"�l����F]1�:��]�3�6t��4�i�0CF?՘Ȼv��"��Þ�ʧy��B˿/..��K�ňp&ȵW�\9�&��e��fR "���&�<�H��B|����ȳ:�-A<�-RE�xJ�n�aI��E�}d0Eue0q��(ʊ�a�S^�'E�aVt&B�s��."jѿ�F��l�aL5�	f������@�J>�u������%�}��L�����c���"�閐���h&��}�ݗ<��C��۷�>Y�d������:Bϲ���-�?��:u*=�L�i���Sc���ma����G�%��`�b�z�u\�#|�-���Z��g�u�`��:ϔo_����~e�F��<�2�R����NZ�(��{uY���9���>�ᬑ�lN2�>�u��w�a�-U0טMw�(z��A���9dF�D����$�I������5�
Fo[�1)yIE�F���uƛf\�!�Ba��빻���h{A�t�m��3��.
�-a�;;T��5
m��-��0�:���V�}�k�<,T���1�6E������=ìnz㮩۷�sְꧼ�e^�'o��z�
����e+� ��sd�d��e��ϖ�@���̲�0�ْQ3)�;w�$׮]K�;r�H����lmm�v���!A��/�"���f�ͷ���aG�U���X�N���e�ZE-j#�y�����v�Sކ1ڞ6�s�P�g��B�����a��gUT�$� �/�6�q�2�$�\7u尐O_�Uq,��}%[1޺u+Y[[K?#ooo׎J�Kf\�x�˺O��er��ٳgS�ĉ��+++���f� �_0�I,�0c.�j��d��z�之��iz�i�����O����3!�m3��R'D��K�I�6{F���ݛ�ݢ�֍�{�����m���)���i�<�{\�HZ�k���'�i��-�e���OA~J��^��1�Ν������[����ϟ?�
d�fJ!�ߧO�N._��8'�f��fѩ�>�|�ܑ�[�g����hKkk����}�!��2n;����h����z~p�>ߺ�s�r��mQ�;t�m�%��F=gaݿ�0ǘ�kۊ�G�	�.[���G;n�kU̨b���|�R4'Aw�ĘV����'�j�`��H[o���5����`�Ϡ}�<�l�(AL��\�~=�N#̲ߡB0�q����g�}�O���3g�,^�x1¤��Ν;��s�=�{�5��￟����jȠ��������4/lY[x�ʛ��wk�#�X�7�&��G���|y�s�XG�y�������-�҅�� ȤI����m�0�<���}`K_�m؋�&̩37�_�V�f޷�NY}�:x|��{`w�dg��0�4e�Mua�+�=��Ma��LgvKT'�h1�J����A�,QL�1yI�?~<^��%�a��믿.�?x�'�%��B0�����?��Ͽ��/��e7n�HIE.-0��oA
L^�=x����z����|�j����T�!�;�>O� ��Ę�D��D��DЬ��4�6���CvkE�_tKF�y�ȑ�ԩSɇ?����D{�-����6	d�����ǣ��կ~�_��+�d��_|�/����9s�r&���(�R�F�=z4U6��$<P�2��� ���3�!��'��AAAA�g�[����客���R��C%�?�x�ň&#�����kɝ;w�@&�������?[[[{�����<��c�'}�C/��X��s�����G�F��$��رc�K
H�K-�����%[2>����H&���/פ��{�����AAAAA�5��d�1�m���<�|�cK�䚷�z+�]�3	p���LE3	~���nll<0z��?���N�|�^0���?���?�9�l����u��Ƀ�35PLޗp@Q8���u���������	�d�H�^��AAAAA0d�b�W�[4�D������'�N#�f�O�>�c��}�Y�	�mmm�?����SO=u���j��?���<�̟\�t)�t��2A�MME3�]D�ӧO�QhR�"����mq����}�d"VA�/�>�<� � ���'��t�j/R_�g"��nZO�:َQw}F�@����g���9�>��S�����`�ꫯ��ַ���?>�[2W
B�I	��?-)	���\#/Ҳ�PV4�*����?}H��'=�3�K��џ�<� � � ��τ�"h�nŘݦQ�2�P-F����vvv��������_�� �~�ԩ?��׾���<ӡ�~���=���U�1L^�ɒ�"���dZ8�nݺ����{r�Y*��z)a��J�fA�!�AAAAA]�bY�8,�iD��`&�Nt�VWWS�L;�h�&�;w�$���z��3����ӧ��/~���u(����/���?�r�J���M&/�T@�̖�2-�˗/���ɹer�
fA�W���AAAAA���#�T,�SMfee%�D�GwM����'�ڙ3g��^{�B0y���������YdB��9)�dA��$�L
E�L�2�|9pN
��w�M��C椐T�B�F�� �a}��\<��6���3f���\�U�2.��-���d}?��<��AL�Rm�ճ�kW�ĉ�ud>�l�}>��c?6���J���C�g��Iٜ1ʾ[���9&�MS������zr��E��p���D��Ҡ%�F�5�]4E��~�ٯ���K�>��Sg�<ߡ̞y�/��替'J�l�(�?c,+��X&��\�ҥ����jJę��kR8*�)U[5͈��A�Y���!ڂ_��ŨA���O����~:�b���6���9�0�)AC�.e5���׮]K�#� &	Z�E��D�Ѻ��L�F�-�K4ڛo�����+��SO�wu���	f���̭[����h0E��s���3�䧈iz�����`&�� � � � � � �Ì
]��˲[4^�z5y���(3��O~�L��gD��F���h3yO��w�^x�~��~/�2^}���.\���7o��eM��R�kD��?)�p	�����^>AAAAAAV��K*��w������~;��O�϶��S]F�MFu�l ��k&N�q�F����>�����羇>ߡ�����z���U��L��T%SH#����'O���
����������fAV�Q�f�Ǹe��Y}AAAA^P]FF5=k~~>}���=�Lu�6;z�hj��ʕ+_}4�"���N��p����	_rVYV���2��(�-��(k��0�D]	� � � � �nPM%{�j4"z�+{v�<i䘠���G�S�L3�677e+�4��A���	f��z �
ay#j6�O���-O�>�*�rf�l�(�fRrO-�qQea�� � � � � ��0R�_v�?��h1�]�z�`�H��Ȧ�֣�|fee%�p��o���K�>��Sg��;T�����iߓ!L�
Y��U4�H4�4�L~u����ih`vk�,!�Ap��>О�ү�D�AAAA0ͨ�B�0˞iV�F�����"Ӏ�,��h���=]�xQ�>=����lnnޫ�Z
"~e�˪����
b���|F4�2����lTY�q�AAAAAAp�E����g���v���
e�3+�}^ޓ`��ׯ�Yf�2��i���`&f�%� �gJQ�YV8�=0����3���~��A�)� ���[|�gG��SAA䉹���zD~A��v�>�KV��n���NEQhY�L�j2��iT��d�����c��6�,�0�mEa��u�d�/U,%�LX\\L�?�����SB��AӟR��l��U~�z0��+H|��us0�}'��������(��ɲ��1v�	�ւ2�nLm�g�.u��Ey�5�Y�ԃ��u,��e���#�ζj��������%��n���$HI���Z�Ȳ�{eE3�k������B��P	f���t)����lɨd7� � � � �0TAA��_[�Kf R YS��N�<������;�.� � � � � � �nϘ%���j2�s���mh.!����Ia�P&�2.,,�Qf��ʂ � � � � � 0��,j�q�?�L�4k��j�?�L�2�H����T�B4� � � � �G�g�AAP͸m��-�_V�`V���*��ϼҙ�LAAAAA�a&+�嵓���YB0�B����vww�WQ8ำ̂ � � � � � ;eZJ>�L�F�����`V�t�L����$� � � � � � (&/ti R����]�&3 )Ŵ��o}/i�YAAAA�ʎ	� �6���O����eE��Ư� ����ҟ���������H�]�1���O���\�UH���M�s��T�>h��xX���J3{f^�EQ������Q�N�4E�+��U�u�T$�2F�[�h���*�vUu�n���w�{]h�iٶ<�L�Ht�C���߱�b�z�ma�1A�2d�R4��[���z��m>�̧:�ե��w�z��й��|��k=k=G`�M��Fٵm�R�sx��z��9�e�[��J�����56t=���~���Y�Xm-;V�a�_V=�Z��g���9�?�zJ����:�7�_d�-��5�~��� �u�4ɜ<��d��l�Ԇ��[6J!�DC�sq/���*RU��� X��:k>�s�>ǾG�{u!� �$k�Ѕ��X<���o��@`=S��O��NocL����\.UϮo0ۋ�1�՗� ����х03?ˮͮYx��Yb-�Z��8��OV���~H[8] �]֘m]�-�D���WYC��B� ����z~��G'-�`V�q�� �Q��`�<���&�0&�FY-%/������6Ip��	-Q2�%��W4)p�D�ϓAk4�o�	�u�XG��;���h[�V׻����b"Tu*�x�Ѷgi ���=�E[`���r��PyjK��6X�X�,�{5b���h`��@L�j���=z�{K}&$R��YddmŌ���ɠss�u��h>1�!��=d��o�sE����ta����}�˵?Z7YϤe�?���F��h6�/�0	g�WB0#���H=z4Y^^>�P��L����{kX!��&�m>CS���h��-c����;悦ϑ0��!�`N�Y��X���|�#<�؏����ڠ��еv�h�^�s֞�m���7��i�n�k��h���h�DӲta�{l'_����̲�Q<�=��ڞk4Ma��=�ڹ�r����Wy~<R�D�Ъ��,ebY�g]B0#����:8---%'N�Hj�Y�U�na�a��G!a0E�����b��bY],\k��p�߉�`�f��FH��4�8�Y��9C�q]X��,�9��QУ8��52��Y[�9�s\&}u`3�X�u����P��sL�8�o�b's�6$���<,��{}�� ��Z�D=���:?��N�=�&�:��0jt�lϘ���1+�Ŗ����B'H���'�o��I�n̨`��X��5����:�-��'���`�D���F�^d1�����&��UX�:�X:�x̬�7�B��yK�ooώ��,������s\�9��"�l����1��ū�ݣ(j=Y�[<Qǫ�����c�Թ�Z��s˸�[Zu��,��c:��h�|?�s$�����o߾�ܼy3Y__O�E����(��$}af$��E����F777�����<3A
	9O��-Y���*]���ڸ��?��R���-%P�[���r/F~���4j#{��0�LV~���=��R0c��c$��|B��,c�8��yo<�+t�e�=�i?m� ��f�H�q��ģ#���X[Es������7��j�@�M�9�u�z/�&�%l� ������-w@��è`�J�� ς�L\t�Ν�ҥKɹs�˗/�uHt�T��Ԧ���F�i�ϧ�b��Au�)3�1�K
S& "�I!��e�8��i,b�Y�`9)����ǈ�:ޛ��f�1��Σ�}&����H���xF��~�3=��J�s˨E4<�s���� �����h��Q̕g�z.��k�f�����k��$���z�3�m��t���)VF�ސk�g���:b�
�`�\�
XH�ʚ�X�s�X�a�X�x�"��ra�w�~�c��G��:�I��жg)d
u��$�L�_]]M��:F�ﺎɊeeh^�+/�5)�̈�`�ꧨ�N("�����fb-�0A'�����F�<gz)뽲�7�.�g�&���Ú�g�0��ν#3���>^�}���nǨa�ap@a��G�o��s/��r���71�	ӡ��%c�眚f�h��%�_��Ҡ�ĺ�X��]�Y0�9j�e���=�LLq�z[Jo�#	�u6�z ����hRKq
}nV=g:13�����2o$�*�~"����ի��r�ȑ�=���3�#+�e�5��ˡ��V>�h�X͆�X&/�*��̤Я]�vP�E^�M;hV�6�W��a_�뒶�Ӥ�o��D�Ϡ ��n9i���e�h���:�N�,,=�Q��Es��)tџ{N��,�֋_�Q��(R'-FD�����z�DsY�������.�Ÿƺ�d�9�A����x��`mYȴW0�Q�f��3���.�Y�*��:N�M�������)���5,�r���k��4�Hv瓗��F�	��d�I�uV���I��B5�NӪS?�`�0.�&+�i���L�̶���ߗ��?po�>ߩ�@3��G���`zYz���M�`&�F�,�	?R�� ��2�X���ȃ�
f����[]<zE{;�Wa��VJ]�=��*�f��@oLs=�縖��b-`�a�s�4����̴V[g��֎0#<�9:�:�����ۢ4�m�}����^���|ٺoѱA���?�,--�R`Rv����}/�Y�ڱ�s�`f��V�����$]�2y� �js�uV�T'��4�C'^L���z���)����&X
}��[���%�m4�K�6�ș>����vn)�!}'������Xl��qqς]��τ��ۘ1��D`���d���4�\�}?�z`].ְ��^��+L!�2�ţX�Ezf�`�G��|�F|��|ȹ�,{�[$�$��K��7�kBa�{j��#�tM�=���X;ipRf�/�l$Z�0�Q�kcc��/8��5�B�$f-h�n0bܧ)�af=IG����\`z3��Qv(H~Z3�2���7���#i��%С�� w�qrA@=��- ��Q,��ж��'�֙�.�;�A�v� ��2ӳ�n@@�i{^یe�j}��5�(ʤ���aC�5�Z�O���E�7��R�Z��SFQZy�NTQ��*����y�����%3���^����hE=߬����j�g�ل�;���@=�L�f�_��؛�
�=j4�J5."Xf��v4��0ð�"�Q'�gbM����=
f�A���OǑ�� ��v�m�轪@��e��@�ЪqTk��mݮ�`�Kft9rE�`	�g��q_�^����a�UÀ�k�`m�`����������6�Ff�3�5��ta����-�Y�kGo�6����r������HzM��"�5�p�f:�2�N�9C���A�؟[#[%�ye��׼�]Ǳ�L4o��`֐l���0�ߥ�x�رRQ-��儿Q�
���T���i�]�`�L�5HZf,�.��z8��"��	k��<;3�Ʋ�t!��th��ڱ�(�2J��ⱞ3�|��g�}��SF��dg=�D�Yѝ(,�#��z^�k�u-���݉�uKF�S���XG[�Q���:�<)�ˎ���)J�K1�(�6}N�U~֎0�c,�����O$�H���\��E�e�*z�.!�5�H(�)�{R�r�]ѿ���)����M�����g�8Al�=X��:����\��>��"$�}S�8fT�/,�E�h.f�+��HW-����:^X�@�*R"�9�fUzh�e��=��I�5,�����gb����e�c���ښ�K�f�	�\��g�x�_��^_��ڙ�[~��!���?2w;r�噐�;5����#���	�(-)Y�U���`�)�{!X�O����Z5�D´^ih�?�i.YM�(BM����z�$��(S��*_6�,߸�������,o	�%�ο-��}�F�1�)&��m��!S`F����!�x�[G� 0'�h=����m���2kOW�Q��ߡ����z�i2�A��Ne�=o�
���p���%����c����-�о�����B�ezL'�.�UX;$����9�W�,I]�V��+���`���8�0`�g]��<.���L�[_�S欭++����)Y�mRB0#R�Zf����J�����U%�^H{��	fٿ��	1�2��g�̅��3�P,#��A�:�����a=g�׾�Y.L��Ҡ�~�q�s)����!�Y��"�}03Mf>{:�Z�O&�$�G�1�����L�㭿c����*�p
���NuҴJO#J�R��sUz���q��kGk�y�����z���G��s.�t'����m�O���28;Q�RȢ�.--%�N�:1���Ȣ�*��Q#�%#�d�ژ�q�'�]3�:��:>���7�[�����ZH���ˬwm/Z��7�	��CYe�n/��"�	]�w]8�X�W癪����G�؟{�ژ�b��3=�Qڬ/M�^�`���Ol;���E��M��<���`fَQ�gK��iٽ�ָϔ�<	t`�i�bXW��h>�"̬m�\�DuȎ;����N�� �?�"Z�Bv��qcVf-�,32IA5 ���?~<�0[\\L�S�JX��cTk2�*�@BC�=vj]E<)c��ƾ���5}~&�����J��}^�fc�W�z�[����>�u6���΃��2�h���w[Gw6M��xlݿZ����atZ�et�2{�z��<w���f����������u������2?�ډ&�sk����a�D��\Vض2��:�8��O9�P��FD0���N666Τ�ϫp��T;��j;Wm%��>G��VEf M3�-��U�|z�[�7�e��1�N�e�% ����z_�}i�lG�a�U��f}��.��u���~N* M�0�LpH��A��n٘uBRm&�ֆ^�YM�j��)z��=�k�'_��o��b8�0Z�ʾn]`=S��I�z����@��5,<���2�m�J��N���c����sY1��,Q�'��am�������<l��ؽ�K�� ���3
Y�L���pJf5(�&���lQ�aދ���T�1��~x����yH��Q䙘�2��E�mC<2�z$��Ewv�Ts[V�$�OK�LR�6�qky��O҆��~Q� Z�Y��WвC:ֶ�M�D(c�Ĥ��,kWQ��ҶH�2�À�wz���6l�����"3c�y��)亝q��y��n�ҤX�5�r���_�1���y���h3A ^�Q7#�z0�[�H=�ۘ��뿆ю�yΨwuv�`�3����}��z*�#g�YQ}�xlWLX�x[�M�����b}Ft�bsss�t~��Mf YO��0.2���8?0�a�B��-�C��L��U��u��y��������䕘�KxA��g2����a*��{�yc�/�Nw�~��o�uţ3i8DEX���W�ւ ��U�k�{�5#��P��i��˨7�>��5M�>���:�X�;��>Sp���c��^'��$V[oV"�i��]l+�qB�a����'q"h��������v�,Ĳ>e��V��l���.&��$�J0�7P��iOo\��j�|��W�s�a���.H4����C�{�	߇��/3V����I��c$>�E��Uel����r�h����'N;]�gF�
8x��|�1A�g�ם���g��W�����P
fM.tŢ����{�H�&mQz�A�M�kJ�y��}�	c�EVU]����O(�m��8oѤl���Սl�£�*M�M�죆���R缰q0�Tݶ��<a%6ԝ�[�q�Z癊�MڀeT�g�A`9XZ�3���+c7�I��w�к�sX��Ys�I����LD1�C>_ۨS�5a��,�g�͠��eש^��-d{FA�l�(?ggg�c��T,��d�ft�g�kah��}���C鶷��maa!YZZJ_���C+F����,u��T��G�i�5H�!τ�9:!Ϯ�zRк"�<�^,Gf#t�9)�v���w�iH^!e��9�3���Y�d\a���:�s�;�Y�X��c߂�c��T��3�Ҡ;I=ȿ���e�jsn�܋5���b\Ús2A�D�8���_u�Y���Ԭz.ߍUϙ��X�1����Ǫw�fy��X�s�C���k��f:��C��s������^ej��C���i�<g���Z�OH=��lsm\�s��<R_�g�u2WD��qMљUMa>;�&�A�6Qt]�̃������<]l��=��H[���O����:�>+�e�����g�zy�{���um�N0k��F%�VC�������dmm--�����B�,�SPaƊ.�>K�M�r��>7:��k��W��);H����(�E��P��Q��s�D.�e�C�sL�c<Ð�`�	Z�^U}��xê�cJ�~�Q����]��C�2?g�����.���@�^�Q����B`:�!0�Z�z�U����9��Qt���ȳ���)�%�3Ǘq��:�Y��7U�1�L���ۖT&X]�_Y}*,������HK@��L<
f�S�|�w���l}�ƍ�L�Sm)}�����&$�idp]ke�������9s�Y^,�^3ek÷u�K�몰4��_��S�}��3!��sE��&�MYoA�xF1���z2�:nXzâ�b����k�ٶ�L���l��hz(�>�5^y`�L�[���@F=�-=�Qؑ��2k#:se��Ft������f�}&�\����l������eU�X�9��Yھ�����O�u��8����A��u��A�~�Q�4�I�
飬w��t붅qK8��j_��+rg�;��x��+��~Vu�6���R��Z�ZyD=~��A�l˨[�d+X��,C����؇v]��ƚ�X"]L�o-V�G�o��Tvok�
r����:�f��f	c��'�,�j�b��L�k�6&LC"�Y{�[]�eg�'�X���'k�����̭�=�FФ�1��F�*�F{f�gy�i̦���g	��P�v���F_[�'Yv��U�� �ނΑ�����z ����������]թ*��ښO��e�Y��.z~�$�D���٭��!�,��K�<�l��� R��N�J�����잙e�Y����	8z/K�>���X��<G���]R�1~�2�`�j�u=GΛB�@@�nW\�LM'qM@����q�f9-}m�B�<G�3�3'��"o^�]���q[\�qm�,���9��yY�B����q�����ZLA`�'��9o�q,����k�/����e���>��G�?s\hC�'\X�C�1��	V�Üs2���`�hu�dE�IV0�1D^����F�ɫ�煲| ��& [�j|SO9ݎQ�,;v�X]V%�e��̺��۟��D]��`N-���ܫ
�`��}��h�̰2�x�O��(V3�L��h�c�Ok���Qm�g���b�)�i2�����k#� ���������z�:_���`������Q������ޜN��Y��W�򊙗���
a�N�u/�>�q����H�[,��@���Ǹq��5*����_̱��5�$}h���Hn�`��)�ND���d-�fz��薝�f�a�!�5 ���K���3YZZJŲ�G������UY�r}UcE�t�*�� ��,��X�(R�g׭>����ހy��+H�B�j,�;��Fd�EQ� X	�g�|$�	2�F�W�S���U�IZu��/�,3�zt����wUd�e��q&A����YX���g��҆��>B[� ��Uu�)n����-��s!,@��=:�"�
�v��6e��@_E5yn=JcR���A˅���:���[2�uS#�����7Q���L;
kK_����l�{1m$LQ�)2�Qv����)�5y�����K�����t|�L^2O�z&c�����5���ü�V!��Y(�	�
g��4dPX���/gv�TV`R!��-��c����PPC�e��t�[������됅��	���#2�����|��u=�������X0�aM�m�|`��}.L�KA[�ƽd�b��is�P���Sb�Fś�s��5k���Q�x�lH=`Y�b:|5iE�a�#�OUu�9�fF�Y���v�^�2�!0׳L�5輅���!���P�*�/�Ḽ���㟥�¾ˁ��!kl�,��i�Z�K�K��h�WL��6�(f]�SVW���:e<��TI�_W�f}O3�w9r�`^����cfm�,�!�2�7��s��;�P2[#/�^���B�
f����@w����$�P���+��}�
�*��a��{�:fg�ܪ�!������#��~h�7�&��lX�o
k ,��EQf�g���hz��L�۬���^E��WX֋ft\Mʷ��D��:��Y��d4=V�J~�5	�c:�2 ��0ҫ�Yl9~����|]�41��2�X��u�/�waDg���]�cE�xl̨i������C�����)�i9Y���8�0��� ��A�g��ڋ�����ѹM�g���`#!�c��b����Ub���r���x���K^�Qf���KE2����L��}N.��'c���|����wF��7�,�-$����n߾�l��$sG擙�Q��_��O��/$;" ��I��&�uӬJ��6%e�#�B�ep@�;av���h_F����$߯�h�����&�NH$�u�ۤ�����qQ��܋���am�nB�}��l�{�ϭ�&+:Y`-����j{�8[u*d�}�}C�<.J��L�6��E�yS�B`�������
Ĉ\g��2
" ���t��wZ
y��7z/֢(�k��y�����=s��x���S�G@�k2�h*�N��M5�d~^'����E��R�E����H~W��D��5�k_Q;����z�~V�J�;fWo�s��%�����k��2d����f韣��`6bo�F����(����d�\rdvT�3�AG$���d~TгR؃d�n�K�ٸ�.���W�K�JX?W�F�"<Fi5񨰠��$�{�6��Ԁ�L���~1K�̣Q�EߝXm�#���B�n��^�}�3���g0*���c?U&6y�V�mݮ��a�G�ܫ�Q�9����L���t�ԡ���*{�I�7�~_$��uţ0�J�����MYG|#X��iY� ��;=F_��k+�M���L�ئ����fzEy��I������n�G^=[�wy9���r����p^����?(N������f��-��7VL�ӟ�p��_��F���+W��7;�M�������߹��w��ٹ}nL���d�h@��aܯ����X��]�T��c�s�e-*!���g�u=`������U����Ÿ���M�Ú�׾�#h�d��}�<�o�e�dn��3,�(�����˾�̐5����z4��2�Y�Eϐ�],��<�M�Ϟ�37)��j,�sѴ���.�v$-Fz��Ho��c�sЩ9���܈=T���:�L�},���E��-�ysM��/��9�hrݝ;w������ɹfh]�|R�*����C#���pa^�F��]�R�+կD���KQ�,I�D3v8L�����}�nQ�}ܛ�/�������dm����ntY�`&��>˃��m���¡XNr�rVzLPQ�a4�hX�"=f}B�:ZXX�����X�hĨ�W�̺��~���G�st�(�sY��F��A }&&��ж�&uŕ��W�NCH�d�W��оy&V�:wC��U۝�=�ú.���lu��8�y��9&e�C# ,w���f�=�X�i�<�#)��1�c�sEK��.D��gGQ���V�t����<s=��;Y�qE�AќZ�#r���T��g���^�6�ϧg�	٨�:�� ������d�J�E��L޻����9�l_��[I���YO�VW����dv��j4!�;�:2�b{�V����B(��5���g�1�>��M�'݉��ˡ���u��ǳ���c�U�g��Y���c;f�.��`������X�1�(�n�����O��Q�Ƹ�~]Ѭ��Mo����M��a	fmO'5��M�o>¬�!�7�p��l���G��9Y����nޜ���?kǢ�sΪ�l���{�a��	e0H$-��-�K���P�<�:Ut]�=�����g�e�Y-/��=�~>kw��q�3�?��w�H_�L�fŲ������"��h�l�(�"�5�~�L�b�#���G�9;Jav&Ie���676�;�k���^G�.&��0��4�e�j�8��,��c �o�7�Tt9��
dxk� ��|�����U��h��ޮ��cި@�J��A����0�"�FX�ĒU�Y������p�x[�-��J_%�(Z�f�0ZO+L#s_�e g%�0��:�:�.tY����4�Z�J��K^LabY�P�[��/�_�sMa�0�y�NMʹ��Q0Cj�Q �X;C[t<Fٱa=;��{1m$,��%�%h��w��:S0Cҫ����Q���-4�������.����ב#GҿU�(��ݫ콦���y������۞�&3�'b�p�3�ݗ�T�<8�,�3����DM�cp�a�~�������3���`��>s7����\r�������;�?'E*˰/�^5�F��� �c`	t��O@@�����=T��H'�����a��<���c��h)�3��0��M�̢��ں	�ڠ�Ѡ��z�#0��<�X[��G���G�Fm�m1�3w,���e�ĸ�V߅ѐ�Ɗ@B`��х��O5}��}�X����S�w�-K����sOX�u��\g�����y[�Z��5����h�7�e	�1�x�z�5_FEC�f��0׳}v��r�rn��_�u@Q��/���i&�qh[�ևl�M�B�F0����s�{��(�f�f3����Ɗ��]�k�M�}��V�C��,����x&g�)߶wwF��$�3�ThK�t8�,]J����u����]K�2�� ����"��=A�`Yƞ����1������d=�X.�K�g\#0�"�y\ �{ڿZc9���S52�I�@o�]�3�,!A`g��8o���>�-'�2#"3�1�hS4,�����׍�~u��ʷɶ�e��QE�ci�Aӫs?̶^E��^�iΫ6�&q�ϰ�+�Y��C�/Cǎ.���Z�#��ɶ�;�"͖��Ө2�[���i�O�ܱ":{��y��	}O��&���F0�v��������(��w������d��/2���wO%�B8�L�5�Z�J�`��mve&�e�t+G�v�n��e���br��������Ƒ���!g=�V�-�aN�=����^��ఎZ��ڛ���i �	�̆=��b�G,�mx�O
+=��v�Xz�����`և�_f�([������r:)�skP��b�������=O�E�}�Ώ��jL�s�Ϸ�ߡ��y����X�|&�C���º\X���Z��׹�P56��xe"Y�w� ��n�(�Y�>"�Id��������`�=-�6μ�x��ٯߺ���o�XIvWV���|z��ܨp��3�J�0���]�l_ ��FI�'�1�����`w'��̿[ ����i3����K�*[ؠ���`�ƞ�ދ9	賡�
K/4=M3�`=��������tH��z�=�ʼ����>�ۢ��u^�\��lfxc�"I��1a:Rd˯�3��0θ�v9g�f�����rkN��M�^����)�U�"}��b�f`Ϸ���~����������8�Q @�wM��e�u�>��s��$Y큹�:�򁙟yQ��l-#��:{���#X���.�p&�ͫ�?'�H�Ίe����pY���민���+Wm��Gv67��6?;l�������_����������흭�W�]}��s����'�ΟOVWW��Q�,-/%3ǖ�Y)��K�Kf�1��1z����d_�mE��l���d{}#��3�vqf���])���Z-��3��+�L����Cۨ��^{�w���`m�G�Q`/N!L�3yl������2���U����i~�ᔗ�uԴu�im\d��{ui4+s�C����=v��}��biPab����U�|i;j���y��Fmk�e��d뱸/����b���&u��m<o�|j��G��A�e���ÅuEᴬ2�,E34�:�Y~|W!T������T?�QaE����=�L�f&s��K�/�&�X���믟8��O������>�_�����~��������dnf��_H#�D� ��7d����(��s�=�͛7�k7n$+�+���v2;?��I�Ǐ��f)�ٙ���'�+���/��f��ѵ3��퍍ѽo'��;ɂr2��J�rL�����AAAL���GCJtIQ�Bm� ��#ƀ 8��rkj�T0����Λgw���������/�_x���w�Mn^�����$�s����0�M��*=�V0K��4LAO�K\�%G3�pw/I�דM�3�,�Et�^F5�{�ү�
f����|2��K��l'[ۣϏ�}�葃����wC�]1.� �LL�� ��0�E�����n��ʶ��\����A��.���>�1O��#ڲkY[��P0{�?����;O��?}���'wn�Lfv��	w��M{����dva!��`���dV�1}S�O{v���@�@�M�$��I#�FO��2u{w'���Ir���e����%[,�����`&�jq���ޒٝ$Y���n23�M��f��b�]�WņI�eA4'&�D�c�1!�3��L;�oA�&H�Y��"�?AL'����$&��,�$��9wn�͗_��s/��\;�n2��Jg���lrtn6Y��K�b�X��p/}͎��9��B0۳�F����*�w�G�D��f�4�� "L#����D����������n�8��K�F��ˇG�}~�2���@�d<���Qc�w,�Aax
��.!`��c�E=@�0��d@�s�b���i��"Ʉ���>� ��A0UD�ӏ�c�g��X��x�K�ٵ���g_~�n\����K�]L�ffSqh6�KfG�v��a�/��y_�Ùэ����7ʼ��l�^��U*��%�)7�=�ⳳ略�,�jo�:ywf�/��H�w����`t�a��;L�Et����eIrp��s#D� � '���a�
���U�����k�s�1��ݣ��/o�VD�m%�|�\1`�Ų����������%����¹���[+ɉٹdy�::z_D�����w�-SIH��|0<���J���JW�>�d����K�S�ۏ*�Kw���跙��Ȳ���mw�p�""�B�(oR9l�n�x�5��?	� �ExHA} A��8Ѭ����A����&�A�=�L_Y����_fa������W��������Nrtn!���Mf��i��C鮐���%�������8��,����%�ro_�K3o�/f�ǔS!-�"K�5ܽ�0��X&g��B�g��zI�l�8?*���Q�f�ٙ_�Ø�'��|�����ptEx��y���_bA�OlGȥk�� ���*� ���`��G��h����.?�,�}Xu��w^�^^�"���M��[B4�D�d���L2���Hg�A&�A<
���$@ '���86��E�"MS�%y�y|��wWzUw�>��u�_��ާ~�|��]U]�U�֪0,�xB�ݽy�o��/���|�Ƽ�n̋MnnLfvyV�'45U�_f$Ģ;Ǭ
Yh{���D"2$�̑a��CA:���׊��5	V�g�z����.s��<��sV}.�Y!�
�msS�1��̴ǳ�r�	8�$ަ/�1i�OhG�]�	L��/AZ��]�־�B�<_"xxȒ!LB�D�c��_{�k��g�k�7e���M�e<���!h�]��P�:�I\ ���B�.5߆�Զ&,q���]+�mݬ���������0�Wf�]��v�A+<Ms-
C-6�k�o�۬{F�<!���_�����?�'�W?�Wf<��vW���H2��;O���VX��첌�=y�����K$F	��I,W��=�a��4�+�_Eu�<�%$a���O.4���`�G7�MnN����ά(_�<�M�<��"�亍0���l6����=C�B{��^�����6��aa�l@y6$�5άMO�*����!	��2�L~\�-��<P i1y1
�(��ƇJc�:���킜�B���g�!y����q��8�YeBd�X�%D�3h�2X�ۘt���s��TDx eo�m��B�|�������_�����f����2��v�+?�ǒ��{�e�)�L�C�&��S���Yy��5���� �ghˣmy������9tMEyS�� k��5s���V�2��=������P}v������S�{��Y�PTѼ����˗/Ͽ��?�����K��n���x���[��u��Y~��ˇs,_�	avzx��.��N��L.�U��5h���ރ*�t]�O��v89��8�@�f�l����z}B��k�>��e�']um}��-ο��V6D���[q:�cY�B��Yn���y��Y�m{���4�ج�e hN��DĀ�%������5��a8@�x���@�~��OMrl��DXs�6P�,[�x�9xh<�\�Z?�*f��/:�5�.��б�V+s�2E���c#̖0�b\3�:X��vM�l�6�S�sK������`zrkCS��"w��c]g�4�K�՚$�\d|��"�B\��+�ߐҜIJ � z"LRi�*�1����eX�ԓ�_��<��Am�e��jI���o�t��aC4�+���6�r����kP�@�߽x����ܸ����5����ݻw����<�2���x�ט�4�4$���׏�c�����5OO��`oB�߇���:w��#��$��X��n��Ya���On��a wwWu�+7t�Mq�z21���g(�!hn�M��].�]s��XS����]Y'47�K�Cy�e�޸��m9�Z䵥?�u�I�3f�9���`�I��g�$ʹ�
����ay0�9o.%��ʊK�B��|κN[�2��Q��`�%@��<�����gް���@�S�.O�1��4���P��Ìd�/!+�t�m�L�Sɏ�_�:GX�	�w����7�kv�l���xgA�w�XC��H_y���Ӆ	$_�B�ɽR�ҶM�m��e��8l��8��ۿ����7o��pw�	Ř��]L�ּ�ɻ˅ ����R��u.$cPB�<$��*�F�{�U�V�t��'��DY��5@Vy�̩NҺ~����|:�'9E��V���Kх*��C@'~t�j-���7Ol�XS	�1��ŵ��sl�bK�z�2~�>�J�b?6Ou�'�V^L���q�
�fֹv��x���K(3h+���G6a6Dr�yI��ӗ�%k��kb]c4��)u�v=J�i�O��:Z��k��c�d鮦���/$���E�K^C�}���Xkۘd���c�b�ǜ�XD�Rk��є}Z�{m�Sf?��/\ٽ���[B���)���%{�ufa�\�avw��7�_�I��:{�0����`�9�|�Y�e�13���0�l0H�)NU��e5�W�v���	�����*�L�óV?�/G^{WU�Su�m�B�m�|ܸ�?��ϟ����d	�M�YYPu��|0C!�B-&hc̘Ҷ�E�f�2� ֚�kf-�	�m@���<��tn���V������YdcX�]�lrC[��[�b��������yY�(EcTT"X�1P�1�51?���X"�0u���F8�O)S��Ț5��8ff�{޶rL���:��#c�i��:Ӱ�L]$�\R�hه�fXՕ���M��B�yc,�+x2ߗ;���eNF]΄�ݻۯ���s{kJ���;�+��DYVN�/��)��Z�7>kM�U�|�Ƨd�oh{��b����ȅ+��e�ճ� �;����kI��O?�ԝ��mw��H+ޫ���x���rQs#��7J�Ȭ�
����A�(�Z*�M�iA{��=bR&��t��֔���Rrv�y]l}���7�,�h���ʋ!0�!�s�гY@�J[��g�&Xχ(x���#�>�lj��X���&��b츚�0C˄ 1�E�|��W4�@�{hZ0�s4���$�}_���S��zU��5�:<g�1�'h�-a��b�U&�L1T.c�)G�aܽ�?�D^�lz��/����pav���7�|Qf��v��xu��h2IH�,��a�jrJr>�O��$��˂ЊYnҘ�0����3Z��9'�v"Xټ~n�H�C}ݹAO�ń����W�̋W�������R3�*Jʣ�g	�6���CC	|�`.����V:�) L�m�ej>�X2!6��WX�%����"ȧ3����9��m>X���$����1��TB�Xh~1�Z�k6�@��;���)ʙ�L�4�g&��\ن�a����zA�;MB	���g��u/�M�i���~�1�2˄�M��,ڄs��m�?u>o=�1H`=J��L�.�Y���Ѿ9����ڇ2��?�L��>4�g>�'Ԑ����y�ߋ�o�1$㻻�ܾ}k�3!�6r�猲*��Ͳ'�W�m�2aӲ��w�{���"̬�i�YV�\�4,�{� ��k��{�	a��e��Qs�Y�H����.�����͍y��#�$Ň�;ft��J��Va�� ��%� `*������`Y�&�l��$���*��FJ,A$����s9�"�&̘V�,�cA[y���@f�
�RZ�L�E�f���̚�b�q��xs��m
Htni�;��sNd*������)�yx�\�H۸�)���C�)�0�b�+�L2f�a�CS��R�3�|����Qж'o�gͯ1�¨��"�P�u�A�ަ�eͲN9C��y�~���L�1:rL�����.<��'!�%%_�}�kʗ>�L������s:L^�L��������|�7�vf�1�K�ҷ��� ��
O���,y�:V�?�^b�!X�*�-3�,���Rf�f��}�ȹ٘���<͊���swwWy�9�������mK{W��eb.Z��,e�gʇ�*fbT� `ZkZ)k�Isy�\�)B@[���S�]�c?`n4c}>��C��Ɩ��ϳ6+K+}�^��.�r�s�6�q!�͊XL�oI��k�!�X���i��)�1�-�f�l�\>��3:�b4�d�'T�ga�~}��so�5�{z����@ӈ���jy$ y����+,�>��2��.,"a����{Q³�[����5���	M�StN#�_jpҖWߚ�!�@�C�)$)��������<C���dY�(5E�p��wo�|��ݭ�ee�dR�����&I�����*��x\��m�B`a=ՐЏ�c�6O:}(����ΓJ�Xêl)�盲^���ܘ��d콭ϓ�J���c���T	����gcǃiV��I%JX`2�1�)��
��üs!E�S�t�e���Y��K�̛`*�X}X3���A�AT`Zcо´�D�f�um��д`���ssn�*��"�e��`�5����u*�����a��!@֘���9�k[�3���^י�N,�ᲆ0u�w�]�/YKP+l��[H:,c�!��'��O_�c~C~�`���۞s�GdSf~�30��2����pӷ/c�j��]J}f]2�j4�ҷ,A�k�@�L�tN�r�ؚj(�v2���lHn	<�'{3�@;��
��s�S����zQ����2p��K�|g����Mq2�,w��O�x,3���������a**I\�j#�<Aw)|��`���2�z�|��4�s���QV��N0s�����F�H]	Y&�"�a��з�WB﷧7�Y?�� V0˭�\d]�I��1-AX�}t��X3���}`�S�M������ 
O�P�i�Z_l��X`�-�w������Ơ��!�]{S�\Ӑ��Ĩxb��59�M�e �bJ��6hfh=1����BL�bͳ�c$��s��6%s� Ж֊)$�X�a溇x�Ĩ�fB��Pco4�.BL��X�<����.l�ED���q���w���v��2ɜ/�ѝʫM�'Ƕw��������ڰ��eeZQ��#JL�P�IV�Yu���B�U�`u�d�9��<�q�P�_̳*����|�9,{�%;6uHFQ)��˄,35jk��ڻ�-�y}�[�o[6��n��~_72��ℶR)F%V���NX�)ӳ�&��*�4=��<�b$}�����=f˾!�Lsc�m}�:�^�V���2&��l`��c��2!V�LSnA�R�	�>��c����M��r}�g��]3�X�ę>��i��3��:3/MR�C ̐�4e��eNm#�1cA+?4Ϧ��޴��&�|hF�,/�/�S�D=̎��YY[���3�`�1y�q�eE��+F�[BU_d7Ta�d���=ʼǘ#��̲5���]���
Gnj¬�0�p��c��L4��	�-��Vg�eV���O��a"FO&fZيpCe�+^��OI��PA��0-,��#�b��A��"�&)Y�0��#^k!jô�6sk���&Һ>����t�^�C�
�=f0��Y�V���kX����T����6�ac#sQ4C�׀]�,� ]?�y��Vjk�d1Νڲ�8M���k'���4�;��d1�]�T�d�%_�IQIO�vo޼yc޽{w&�����5f4v�q��ß����QB2.$�n��|�1���B2e5�djɄ�W�0����|�D�|S��ܕ�*[� ��^Z�L���Gv��\ZB�y����2�0s����N����o߾1��o��:�t��t�{-�V�1�>��v}2� ���}� ˃N��S�3tQf�c�:�i*���U��jY�����h�Mv}�y�Ũ�@�2H��̛�@�%�5k�1���"`�e��E��L�L�,���f�F���f�c/F�h_�Q�9d���~=�r�d���cB�H@��^���\ƀ�9ʾ4Q6G����φ'��uv��f�3�a�54~��Y�W������?7www�}���߄Gi��Yƹ�G����ǇßB���ЌGI4���*¬f]n��eO�� �Y�GO��Ć}����(�Ryo���>!̤\�<}�;2-����9V~*��L����Ӭ:3M��p<��oޚ��{s��9Y�`����gi�5fK@SQ�����ԇ&-Q���Im�B�T�j{Ũ��V2ێT���E�y���P�����������β,�hg��t�g��<�#a��>"@������Pk&�b,;�L��Z�Q��9V��^����$I���V�$�@�h!6�f�P۰q,�?�:�Ph�E�������<���C�2V�04>ۮk~f����ݱx��}��f��|��Z]y�}��V>��x8>?<�f�����=���̜���ñ&���j��(�f�����w
Wau��'/y��:��I�yR[�n���Y��-\�	1&5!L�4�����}x0B��yfN�Z� #47�1Zo���C���v�K֘B�f�Y��L��[�g@��.,�X�,b�;���>��,F@��t-f,�5m#m�,FK{f�����@�fH�c|>&�k�Z	�LY�lDk�}����il:]�c5�Z+X묶�
MY�C@����%��[��f*�/)�\i1�:��=�X��A���������sݤ�P������u!������˗/�g���ۀ��&{����$nn����O�VD��<�d�Ќ�N����,��D�0����.88Y����е��uv���Z��r��^���%�7 օ�w4硷}�������3���s��'֒v,��"�ŖU.��A�N�ʅX(\(� φ��e*OY�cP�n(-T@E���h~�:@���3EȹL�� 1���M����>_�8��F7~1���Z���
�p�ڈ�]P�;Fc.��nξ7g���ݚ�(���)�+��s������Q�1:�aC}�F6��:�X�-M,v���:�:���M��s��-YM^���f8���N�6�z��4�{}��ً�x�7&X�a�e��Y���`Q�I}�:���=O��r�CMV>f�OO��*�Z��	�ll!N�S��r&�.7�^�4�|�K���k��0Fœ�W
mk�χ䇦�N�1z�Ř����a��e�4H`�\,"���T�k+3Qa)�
m��5kmc���ڞ��N�ň��b�����ӨO��sb��l]��]�����#����7�S������Xט��݇�?:�ƨ�e�s>�$�|zC�az�1ʄ^�m��֙1&$Y��h�����0����7�x�_���y�ٚ��C�s�ߚC���\��p�>&cVOO3GY�2����zO�%f*������0������x�{��|�IN.,�)�IwS���U�H]ljo39�l�lo^�|n>nx�}���؞�F(Ĳ��1��n`=K��C@��:�E��5C��ɏU.�k�@SI�M��8�kU8��@ ����5W/�.1*m3bTXǨ�0e���(4	�K�l^�J)���|�c�9�mbTD���Z�}4��"��˥�!�>��uI�b� !�:`�)�:�&�領�.5�����+��1H�EO��l)��K���4���k��_���fy���0�}����>��زP���8����ܼxn��\r�ͫ��j��ej*~ȑeH�3��	f��1����*Y�f�*���
~�𧝿���nVj�E�Q�#�B�ɽ�0�q�ϧ�MH�\H3!6e��܅i�����O;��H��y�b���"�Z�|	��´� FǄ�v�BN���®x#�Vĸ�c�i�B��i�2ĸ�]"-��i�g�UylSӰ��ז��:���AbT�.����s�='�	,��5��cɱ~��f#]�Y��8�MŜkQ�u�-G�9?M����	0�1$�B��w�|��5�t�������2��y>��fe�*��Ӫ�����&7!�a���di&YYu}n8BGa� i�,ʙK��C&敗��ka��s�l}͓r�����G�0����G�2�]Y���IHHHHHHHHH��n��������������p�h`]�7��W�䐌Eq�U��u�p��<�|�♕դY�H#�K�ёO�6��@�*"j @ �e�8z�2�3�Nz�3�p~t:{仲�L	=�ò
s&�:+����[�ѣ&!!�:���	K��2:�w		�#�													��SE����wcBicød�瘼,p�P��@���pBrU�X�Ly��=�?�򉗛�_�΍��ڝ2srG�叮�YM�e�9��cgYr0KH�I�/R�ċн>�.�f���h�\�XM}3!!!!���6$Ċ�7z��y��}z�M9����"̪��,7�����0��.+LQ�%tTSf�0��yp�Z������
ʈy����^^gO9O��K�^6�C�"(tYf�Ye�V���Y�ƶ�*�o���Y�ph�V����Y��		�$Y��%$$$$$$$$a�3���}�pº1挶>�l,*���]��:(m��*�̑KEuf�C2��e�|�װ�Wu���� a6��;glcl�B�ռ��ju�>��=���@<�$�0�������{�=�				��%L$�3a�H�ԇ.A�g�w�
	3��
=̦�f�sL}V�ƚ�F��?�ٹ�L�]U�eΣ����'*�ve��Ԇ7ں2��� ���0�g�̅Y}�0����Cۤl�Q�·w�.W�j6#)���}�v��4KH�iVH�GBBBBBBBBBBBº1�����d�Wf�Q=���1G��.�v�q�+��"��ʭ���j�p�ܰʯGh��TX,-.�Wu�����3w���t�5O����=��0�]�S���f�ndٙ,�ʐ\H���7)��Cj�e�H�������������������u��ì����d,$$c�17���n�����{���f.��y��]�Bs�� �$�\&Ւ�m�/��
Yo��a.��ob1��6��ķ�=bM�	�XV����9o����Y�e!�����iռߘkE�eGU��β��I����1���2%o�u����h�<���m�]���斮떜���J3�4���nS�Km�٭YN�<�B{�x�u��3?�;���S��OV�b�������������sB������J�R(�sݧ���~7�w�V�<��/�1d[G����r�n�7�}p	��o�)��!�.lQ�af2���*�h*�a4� �&hT�����?\��� :�/3������(��3!�*����A��Yhe��Gא��P���lʲ�N�#���M^�s��Cf���z	�g������+9���|�U����7F,07���|�	�M;��j�O�y�`�3�YF�bl�ô47c,�0�����M��"z��c��2�٧�����#I�m�I���t��YvC�l?�c�)��`��O��>�����澐��k����ycN"h�,�]���^�k���@�0{o�<1�ާ�b�G�l����m�$���a�����-�G{> |����GOe�c������i����<3��[�8���3fk�̗���&˂�����cH�ʋ�Vtu�U�ŬN��qMݐ777f#�Yyӝ}0����2�\HIs*gS6v>PSS24ɩ.H�ׂ���K����@��D;���À6�`���6�J��<s,Ĉ��4x�����d���9�s�Y�}�����~���E斩���:�r��X7�C�u�g�?������V�2�=d9f��95>B�?�|�&ч��ʊ�X�RT��H������K^F�f�L�=�=�V�tm*P��Uv�k��n���G���G�`�Z�<[J�1U'Ӭ��W���X�5^�>�a�LIs,��~7��&Y�"�s����_�}�{�o)t2�e>c��l�YE��m���oʞ�v&�<��ɲ���]Ϙ�����ę�0��2���יx���ߛ�����p<7v���^g���m�/�zfu�"$.XdsC.�Ж2�,	T @�%�3��Q leZS-T��Y� �R��ؾ(X�.m����f(�Ɛ@��c!�6�����H�B��X\�dnY�ה�Fr	��!�f9p�����:bys1���0�D�K~e�wK���C�ʜ������u=�L@ѧ����/o0�
��/?�{�6��<�7e�+����r���]�shNj¯�mc��Mzi~}y�cߓc���u&�{�V���rBZ��nh�}��G�*���j���'���ztκ��;vl�§y��*Z��Y��p�Y�H���O�I���_Z��Bp	!&��|cv��vfW6�~�7ۛ�w�ОݔU:Al�J�i+oڔ	m��y�aZ	^s=i{@0#��Wb�rц��(v��-@7���Y��u� 1a�-��=k^�����-ߵ�V�<s��T�3�����vB��������hٵ�N[G��=$?��C�j����Ciɳ��Oa=��a@[f>_����|?�H��NX{���昿��|�*���I�F��2[VZ��Ӗ��66o�Ʊ>��'�i�P�����0�u�դWO���6>�E�3�jf����Ҳ͏�m?��O�?��c���;{�We����c�t�3���̱�B�ت�Zy8�۷o��7�=�16/&����T�-�]�|L`y	�|�L�16�}���V�|舑�D��L�vc�?h�����'e�@����U�K�����x�X��%�R9���a�jp���*�/�sk�_c%̴Ӻ����A�f����;]��3��y�ԽU[�s�9����T��H�9�M��yŸ51����Z�Y��M��<��e�2������E�(�&�x���x� ��L��kmECYfك�G�d��?��{�<?�5m���L��\l��e*y��B�����$;OT&X�O��	-J�8��۷�������ݥ��0�Qh�.�y�a�mB�rz�+�I�}y>�>�21���US�0�Z4Ʊ��~��I[��{L�Bx�e�څ��J�g-h�+mknv�	<h*�� Rvm2e��.�H�^�r�<}���l�Ǳ��1��,��!��W�=c�ꓣ���E�VU�1�k�&¬/ݩ����c�}}s�������<Q9`���}���r	Tfm�g��gy��Y����>�t9���gՃ��֗/��W����WfO�ʰ��!�*���?:�L6/EE��rY:B �f��#m�ߙ���L�ߘ�f��9�u�Y�Si��3�R
2�� Ԗ���X�*��Cň=��@	�!̥��cH�k%�дD��X^E����lkr�����C�I� �}(�8�/͹�9gh@Ĩ�KQ����>�a���3�Af�Fv�{1>���YH�yEi�F��XJ�)o��f�yq����0[�3��b��F��EV�	3f$��1�'����Ye1�[�m_>)��	��}r_e��~k@¬A���q�����*z��`�=%51���Q�&�ʗ�]�N�"B򣇙�C<:T����<�yf6�n��~o�}��l������8H��he&`C���0�.�,6 V�C��1��NsÆ^��c]2˭I$h#FO�P�Zڱ�<(X�jD�Xk�:׮m�Y���(ɅfH�Yg�1�˘�T,�9��7�<c4�Q1��]�Õ	tmd�%���#�3�Q$-f�kʜ�~O[ߢI���B��k[�L%f��_����g`�1ceӾ���6m�̹�S�at]�6X�iy��Fp͑V�S#����ߔ��6{YJ�-;y����_�|���^�L���+�j\�6���rҲQ���3������S�x���B)����0)�����*�x}�	U�<I�\��Uq֚'�+Z6���$$�ѹ~���擯~��^<��+� a���V�LH�dS�׆�̝�0ɍ؞m�^�H:1n�4&���I�"�ѫO��훚u0�! Jt3�R� �1	�	3T�9T�l���(ĺ�D�b)3Q��F(��km�F}��x,�L��s���{H~�b,0�C査�;�t~e�dD��{hfHHB�1�#A�i����zQ0�"��j�AS��Z���e�� 6�M��l,a�槭S�1�9�ƥƏ(Ya&��A[��e}�d�۹Wx������c�=�L��������������M)䗿�{�5�5�2���̦�q���{*ߜ��V�\Y����+u����/��<;�$��{e�� ��e֞*O�6�^++�\�˻\���d6�g���p8�{si�g����s���Μ��;�,ߗw��*����W��
�h�%],���A��H�d�k��xL�.�r͘��M9��f�k��P%�f��y��c䅖� #����?L¬-�㔶�w�M��2Ϫ��j_[��T�!
�sMcA�(��q����c�]�%s>X�l�L�9��U�D�IN���z�ʏ�a�bH9wI~c��XrC��4ҒkD�@�>mjk+�/%�² �]�����^_P"L߂��1Cձ�X:�|�"��CO�б>���r�XȺ�Hwn}Z�}HZ�:�U>�^y�,4����o��'ڳg�ܙg�T��xc�����!ay�<��o���JA���2S���e�*	ehM���.i�E�8�d�/wQ�q��sˆр>%g�����O��|�L�T�T�1O���yufY}�{��~�]V׏�?O��f�3�]Q�vf��7�	��M�<c�a�Tx���ֺ1��E}�_�W�L��SSAŲf .�C�Y`�u&9���]��.����|�?5�ͪ�Ij���C7b1zo��%�:`zi�a1�ϵ7�H�ڮo�[L�[lm�]�X�,y�5P�k����I�"u0�o2�Vl�Q�N�٧d���fzWi�A�"��䑶�X�gt�d�A����K��wH}21Gۜ��-�K'3eM뚧��{����{�K��⽪)2��`�]@�������tD`����Mc�3�R�W�1�������>X�6�0+y+�N.W*�e�r2�ݶй��{UfQ�{����*�93`g/���{�)'���Mƶf�:|�|W��(_�|W�t�ӳ˲���E�U���7���)�Y�f��Bf,�h�61
L�� �ac�},�F��9K��$�bS�	4-��P�1	%���x��3C�i{1ڹk��u]L`Z�}�ieP�Ld�e��s*N/��2:�3� m�p�pY��$NY�)o!@����c�'.T�ε�P����wc��S\5�F�ϵ�0�,�,s-��_�H�-�����DH�)C���_�kXy"s>��Ct2�c]���t�χ�L=�3�m� 2BhX�����|�fD�;Lk��W��n�N\�6���
� '�>3��f�O3+�����Z�����-�	�a3�A��WY8OX�\��5wg0���"o�&w�c��k�2Vw�F��x̬1�S�Ǹf�u�h*�,7
m���y@0�����.���f�,F(��
����!$��Rp
��Z��?���JZh�M���t�ۘUOHZ(b%������M����O1*�i�<�P�WC���q���2�|̹��=4�>�Խ�T�l	�TS��48��N[�k��Q	��Ӧ�ems���E����1�Ŧ7e�u�-k�!��H�k@lzc����z<�w%m��iaHF��u�}�i(���ٿ�=�1�ݶ"Ȳ� y�����9��o�B/nl�0��{[�Q�[�1[�Q͇�&���h 4�sl�2vQ������e�Tvij�>����	���ʣ��Y&/�Z{�����5T�eš�v¬mm[�Yi&��kXy���1ʏ)��^���F!�6M0�ڇW7�flƢF�]b�8����hZ��/L#�%����c�wL��Z�D�\��7Y�����+��<��v��!�5^���K��.E�I���k>�q�9o�5���-��Ř���OA��ۉ�f,B��W��6Ly�uuH�5�侩ᑧ�ml�j?!�B����μy�ƅb�N��<�$�m�g��D�<�n�_8�l�3֑KU�M���TT�QEV�G�0���<�*��\��'�Bا�d��QD��!H"���Z�gf#w����(\�ƪ�|C�oT�ڪ~L��f��c��+ál�!�5mK4�W�Vt�A�6�<P�G�3����ږ�h���0��PC@���F!��pY�Y�\H=��}�r��T�Α9A[:C��1i-�A��y���:`z���LC�W��ٟ��5H`�}��ːUb�V�,�y^�V�2�Yd.�K	�$�дXs>��XU�-�w�t�C=3�H�X�I���n*!�M�^3����h*�(Y͒���M�]?��|�`z�k�ˍ1��cY�O����t���g
�.noo��ׯݙe��o�&Y�l�6�_o�z
Vf���g7�� !m�
!�QEYЊĒ�2�1�	�S^���_����n���{��$� AV���X���n��tE��6:�Y�Y����T�3�g�>E�V5^ՐB J���wdY��������,7���%��@�֍{_HF�����1m<�"�L���y4��1�큅*7�
$?�9c#���I� �i���1D�Ũ\D��-��9R���Z������7f�B<��Ĝ���1��sd�azr#ޫmy�m�Xm��(1<��WmY
�w�5S��T�L%:�{��@^�$@֘�Ϩ��NS��6rM� 	+��O�
�X	3m���]�9<�.�k�����sc
!�mp��W�PZ��&�:�,�q�A:4-�(�z��y����0����ٳ�.ѷ]�]�I�PV�eꚋ&f����v�3���Ʌ�r?z���x0�#�*��EL�=̊�.h�U<�ӿ6�����!�U�ά9�szk�����b}E�#ú��G�z�fW�5����/̱lܣ)�Kɝͤ�ò�F���A��pp����MhZ̢@$T��RJ��Y�S�Ih#��"Q�i�϶��T*1�@����:E�XL┩�D��.��Q.�X��$
mRM[��`�\ݵ	F�e�������&b�nXb.`䉮1�!���Zejm���z���6"	�,��j�y�o���`�m���U&k����k�/4��m�3��b*���gLcYM χ��K����A�ھ�(PR��VHf?�Ę�`�ø����,l;���|!����6N2�6�1���x�9�*s&�^>a����U&��e�(��\3S�IO2�#˚��S��l���5��Ξ�/�8K�M�ޗ˚SѰ��(����Gk갎�WT�����a��{�Μ�q��7f�/;��A��n�׼�o��8C~Mh+%H=iZ�-f�0��H@�C����!`��3t�C��
V���kާm��	y.$(�X���P@�c���C�>k�	�:���m��FSӘ�	M�hvZ(���=�5����&�����bY�#�Դ�f���f�D���Oش����u��-{�ĩv���;����%e��!�i���[�J�se�C�}3��ŗψ�PH3�����t��6��R�����|��勿_��~x07�0/^<7'{2�vS���ȡ��ʝa�3�<̌s�쨴:<c��� �Ρ]�,�L�>+��������)D��$^N��'��$��ur5y��s�LM��tˏ�|�ȸ�N�x<���o��Ƽ�����O�d^<�F���g��cU�A�C��`�mɋe骭`E�δD�;��Cܾ�0m���X!,Xg���.�l��2	3V#g�!�B	3M!v�X�3���dZ	�J��l�6LA,E�J�����X��u�nZ�-G i]J�/9O0	kL�\+/��SY��9#=f0�Ѭ9a��3�e���T%(��g�c�ŀ&�3&Om�Z��%�K�﻾�~f���]e��ce�rh�?,=��b��D��F�Gx�Y��	�x����𾦷Yy�Z>G�=���v��_��3�$��pB�	uz8{*La+«"��y^��#��d{��Z���y�*��4���J0��)6S�^Oh�*��̳����]�p%�ui�o�&Ih�Е��|��w��(��~g^�|i>����GS�0cmW�kǵ+=Y�����5�$��K���,%3j�=�E�k� ��7��맶�$���1s� �F_�^�X72a����cF{M[¸A�gW�:wj�7�Ls?�%}snk�K�A��a��5�W朿���簾�(���c)��&2m�e��2�]�:���2�5c�[��钫 s�Oi˸��͉)���y4�l;!�nnn�_IW���U�6W�}�<��<W3�0���\��VZa�'s��y�!�eMn��i�<An��]�lV]C�Y��o���8�\���&*O0��>O���W�;�P�������M�˘�|7��l͋/�� ��&����7V�6+L� ��(�^�Q�7��
��f
��ź�r$&hoBPĨ<E��=��P~H�C�9w�cB��TSi��+��O�$xXޫ���|����5�b���ՎX��7����S��b� f�=a4](���]c�P03��s��`���L]cc�b�חN�^{����ݴ�x��Z.V���$���5_�s5s>�.L~�6�7�,���m����L�1�����#L�˲���OY>����*w<���h����ý9�"+���<��U��O�$P�a�Y� Y�u-�I�>dY[�*k���4�A%o6r����:�W���_�N�~ͅq4�L<yҬ�gҬ
Y��&$���ػ�o���n������-�(T��튎^����{I��$��c	�Ǵ�DBձ��b��Ds��$NY���fLA�u���C��5���c�WϠ��� eB�\hzw��kH\tm�-�[�0C�b�;A���I0�$,�V�
r���K�(��暄9#�%��bW�]����D�ľw�Ҭ����������@��@\5�b&A�@{�"�\?��m���Xzm���sNc*d�ΪV��3]�����6����1��y�[� gt�թ��ʫ%©0>�b�<��օ8t^iO"ky_+�����0+�s�N�ɩ�w�Y��]�+�0���RH�V�N&�eű|ֲ�E٠�(z�ob/w�Yn��$�7e'(�ɸV�M�u���j�C��ڈRT�*UԲ�=k�iA>�f���&�Pa)��Y�}��<4��:E��3�;ڊ5��6��@	_�sZ�Jx����k+d]���IMM+F�L{.;��h�����`쳅�~��FSq��g4��Ch~����@��v}�����B����m�rP��uF������$�P��q)i�U�tPtM�7��e:#�9s�G�-ӡN�|�@�X^�g��1�gl+�P��>2��΄�v��u�#�y�av8��vkv�����!+ʩ"�L�eÎ��m����k'������)N���ɲ��{4�� ��Ueun��=���τٱL��<��������E���qn�!*
�l-�F���S�u���X�����1�q����̏>Ӛ�4��H��H� ! �m|�@뛵�fA�@�٧�NL+޶��ks�ī/��ߵ=S��$�:GaX�M�$��֯�Zx���T�j�1C�$�4#$���H�i*a�uc��WK�,�dJ������Lc�����$��exTa�a�0�D��fJ=�<9D��G� `����j��M�fj�`�uk�"eY�f�WY��v���G��0��T�=u2YQ~���3Ǖ��g�,��a��O��s�M����>��|'�|�̴���:�#��P���s�U�V\�T|�]-L�|���Lޘ� ���$�nQy���mU���Aτ`����Ll�3��5�@�1�Y�ąf�hJ�d�f�Rv��D�ՙ�h?����	�D��#@bo�#��
+�D�k:+� RO,/fH���]R&S<�����Bl2*��8oh{_k�xl����-�Н���i�H���a��ǅV~��US�ǹ�����=�!��í���&���0����$���e$���sʯS�3�0����g��%��҇Y�e	B�u��aע��4&���CF"m�%Sz���ԅt��T�/k�Ń9���5B2����#���
����!/4Sys�"�7��7�c��G�ј�쳐��n�ڊ93�I�3�M��&��7�;�O��2y��\�ZSY��a	�d�5�'���1- Y�ތ"���	:�4�������s�K�Omer��Ś6�=70�b�(A6�>-�z�]��憜��%�k.�QVd�>d��1�wV?�|�k�����M����M�hB[�G��#���4Uy��Kɲ��1c�/�)�k��'�hז�l��:*�0�k{����C���K��m@ۄ)��&#0˄��>�7V���qJ��f�13S��Z� ���ȝs�YiGա���Y��0OI��u�_�@��:G�ﰏWX�8q��w��܂.q,s�[���af��.�ow�g�h��t�dY����?Y��m07+k�O�:@'�����s"�9��~�lL:Q�D�R�9�YB�6����:�i+c���<���v]����`h�㼉���>^4�C<x�������R�E�5����`jZ���'�NԲ�ί֮W�Uv�#sB��9�̓`�\�HGӨI���YĘ�Q&l�~�Ʋ����}C�s��d7�A�5Դ�zچs6�v_�|��L�=�����?���W��ߛ�ۭɥ\Ǔ�h4mǎy'3	Rx�͉(k|�$���K��ZMN��3�l��>�g�Κ��f��"�$k�A���o6/L�1UxJ��2�#s'cw�;+��NZ�-�/�>�zr�(+�)�(/\x��p����Dl`[f"L�`Y�YL���p@-k�𡏕�`���`-�k��Yu��s�5�XJ3I	釞���S��"�kzR2	�HV�D˭i��ק�Z�ɬsd|j���BP0��5g?d��)��ؚ�O��O�<f�h�si~KϹ�Ɓ���̫o<)���Q�T��zM�GS�E������>��#���.�~�����4Di~ߕ֥��O��mMREW��қ����F��|��]���+�{���:��3����w��1�wf�>��������O�������/_�6�n̍�JR9��9f��3�i��+$P�l���*N����������k��>2\6�?;�R��:����s8W�8�'�]�5ٕ�M�ښ�����<LQ֓x�əfB��v����&�ʄ�֚Ӷp���YdD����\��q��:h��c%�B0�����b��Դ�ў�D4r���9�P�3'j���J�9��E�s��!�T�<m���b���Z$�v�1�]DZW���u!�d3�9O���X&f~�(KƢKq�uݥ`��M�Ⱥ���R��$�hH���LBw��]*M�ϧ�..I%��������h��X�"SkCP�T}e�s}_����������lS�~���2��c0�c�(��������9�P�����1�H��<�#�����=q�ʶ��l�5�����`6Y�:YRw������+�-wmo�I�}���ؐ��	>�:�!�VԴX�����=���p\�^V�UWn���U�l���禙�Z����h��˖uYh��t�%z�ʒ!0*S�5�B%l�.�V�����_7��χ�	ˊ����%,F������`���//	���oh!eb�9mt�T�k��C�qk>ߜksna���S1�=���\��ڏ�c�
������m�$�<��iԷVRj ����-�k?⩎������<� �� {G�5��V��%��%�.S�e�լk�Λ]ck� ��9���kC`�X2��0�2M=ј�l���O\��Y�&���iSCښuP�&��f���s��mz�y�{��qom�Lѯ?�p���/nn�;r��ݝɷ��n�	���b5�#d�u�RY�bh��������pJ��$��c�LQ�9��\nϯ9�Ͽ*��tr�5�=YMV.j���G�l��ͳ���owe���~�H�C�B��l�K������Q�_,�D��@�C��p��j�	�q1�
I3?� 3ڊv��l�ͺ��GH	ͱ'y���Ƭ�D��H@7YL�U����l]�͵1@�a��f}�M�P:��VZl��H�:�O�b̈́ B$hw����Z��_�5C�"�LA�!���w����^�����1(��e&��G �M%��t/!���uMc���jLC54̹ƌ�.%m�uC����Ha{j����ɋU�������5O��Y�Lĸ�B�a�}��<ڮ�+L��5��a"��<<�扲��$�*��V�L��l���d�x����^~����I�������l7R(�('؟۪�,���rT���\Șp���5YMzc�|�?Ky��KBIVYM�e�(U����ߊ#��{$ʲڳ<f���P81+B<�N���󑰕�\�:���*��A��s#
�]Bi�d���7YJ{����P�h���������o�$�&U�ڙ��F�<蜁���3�=����D���a	+@�W���E�
�S]ss�Ĝ�4�a�?�5,�F����צP\R���+K(�4��$�X�yK�>�E�6�����
Si����eWlks�G�c*����s>���9沩�<��acS�iK�rz(�>H~C�%�Qñؼe�k��j۫�.}�&6bF0v,�]������ �UOlc�p���kxV�P�a~�j�f�x����~�����3s����G �5i�	*O:�M�s?+�5���T����*w�����L΄���3�<�~~�0�A��C1:�O��yV�dƳw�^��(1\CԋT�Y��,���da��LY+�P27�0Fˏ6h{A�"X���dZ�!`Z���r���>��F��P�SSQ��.�sk�A7u�����B�P��Cӛ�H�˫�E��8ߡ�q< �^g�FCCX���f�(��M��#��м�a���nnn������}М�P%��4Jɏ�)��.���{�䅆�g���Y4��͹:�}e���C�1��1Hh.e��$Y���eL��ӳ���H]^�ި�1	{L����mD�'�d�����5��өO)����O���_��W�͋������YfE�r����&�(5	e����r� Q$��,?�>�=�W�q�Y�K�Xz�,����Ӭ��;ﲚ0�
���\�*A�^�p�r�'�<9&�(����[�b��:���`�f=���T �Y����0Cb��J�!0	3�R����s(��,֦�I�:ԗi�r�v���\��.0=75=��
�X�Ӿ��MA۽S�i+�Դ��F���'���}�kL"̦�Ͷ9H����Ι�T�0�U2kILA�������t~E�b��C�Ec�$/m���w�H�9�$����]����Օ�H ���ty������p����ԕ�)�5ˉD�@�E�<?�qꍾ��_��2a����:|	³��y�o�x�����~�z�ѫ?:�c6�ʛ��"�}�9+S�k�ɦg4C,_V�76D�sV�����5�����Ğ'��w�G�����>����*��ĺgw�X���xt!���t:��myǯ>7ű0o���8ɰ6a��ǂ�}�Ǩ�f[]0�t�
�1��6~�! c%�X`�\��Q4��� j�J,d�z� F�6��a�1KX�i�k~,,A�i*�Phrň9��6咦�3�9����C���f�}h�	c�I��`��L9I�4�'1쵴��X�1ӿd�n�����Cנ�KV�B�|�"%4�1�y��{��u�~Ǫ�i�h��Fz7?�(�1�@柇�����������,� {!��{�������?��~����v#%�'(3)*��f�|���s���LKu�Ӽ~�����Ϗ_;O.k+��*]v&�\�����=�q�(�BSVg�Ud�x�	)v<YV]��p���u��|�ٯ��)
a��J,V:,��<�е(Ū��ZH�$�b��0�L�}�5��ef�!��ph��D}"�i�+��#F#�1�a�a��p���W�m����f�l	h��X�2� �%�`�-�v�4^A���"킜�.ߗ֒�p�Z�<�������6����g��RFO�K�.6��i5uKc�@Pٛ5Wk�u|�{�1�F�Ӯ�ж��h����C�썙eb�O�щ�[����H�=̤�B����3���cB���g�6��O	5�^ ٛ�?���˗�(œ�(_U��,/[�hՅ�]�ln�@DFG�C�@=[X���������nh���~/�(������.��\��?�L�k����|�Mn��2�}y���f'+�e۲�v۲���#d}9FA�IN�b�3�E\��b���1�d��M4h���}LK���T����!����:�f�76y�l
��q��$�b]c�Xc&<{�K�lͶS&V�D�����XyiX��X��k#��x�A$\:�L�g*�r�6ю�5ߡc�򊛡��e��?u?��m���u���"S,a3eOU�^�|S:&Y��I5�qU�ڠY�KB�6��0���֘qØ[�:�{��#�.)��C�N[��z>M�hj�a�{��Yu�-y�H}�@�s�_C����d�\�f4p��Y�O��_����W�i~������!�7��82˖��˓m�g巛���ܟ��f�*��@�He�v7����du���'�PV�x�m���;�����3ΤR뢺h��B���[&f���pmrpY^�A�����s��B2J�>���/}jn>za�&�N=;r\���m-��������X��l+��+Y��|me`�5'X!0���I,��d���3$`��W;��]X^�Eʤ�~�)��cf輡-�i��|>��:�Ƥ�m#4-m��}K������k�B�i(�ܧ!i={�l��uu�֥�Ǫsf��b���̜�Y`�k��TX{�fM����#J�-��y6ֳ-�U3$� �+�|�$̘�0#/F��O��ԕ�C�91�<�r��M777�kţL�/�#޼yc����a��_'�Xǜ�=������4j}����f�>��Ͽ�W~�/��o��n���ٕ!�UyQ�t����xp$�)?�c&_������U>xY6p ZQl�������r!�$d��/q�qd`^YO��#�'_˳�-,+��	��)���<��V��~�7���e���ɹޔ���C!�NB��"bT�3��tabk�5a�b��gL�-�v�
�<��11 	��SH_»a��܄�\}��2DHC��Zǳ�0f�u~��btH~��l	���x�<���@�.������t>�Ҥa����4�S�,a�I��e�3��|4�A���`*��y.C0����2j�h����6��&X@�a�p�m��%)�UC�$�0���6?�g���a�M5T.��r���m���S�O^�zU�(77g�k(M��;U�=O[�M��'���o��7��w���~�[��~�������<��}#P��<�ԯ�p*Šr�9�>�L~Ɂ����8�
�B�mvu��_lrG�IXI�w���t�K���&��ȝ�v���pdY�m�i�)�/��S����n�:q��,�ԓm�-�TD{[1."��P �&�J{�>�֓�R���Z�$b,���$Ǒ2��f�Ot�&�4����1ۅIx��cyS,i%ؗ�v~��=�YЮs��Ch�&w��Kb��d(���9%����Cej�Ŝ_����Bc�2���%�2�;�y1V�!����Ҕt�d��s�� f�O�0C}�z�&�Y�$���<c�f��@ۅ�^�����d٘{4��,�������w�A�_�q�������������{?��}���_��X���Ʌ4�
��*�V��92h����ɦ��pʅյ��\y����˿9&�p*N��`��G�5IW�u�י��&���D�p���$g���|̏�Yf�*���V��9���i<U?ٓ9f#!��NQ`\ڂ<�#�Y�����SK�nB���$]�@��k�h2���M̾�n~Yh�7w�G�c�j�7�%Ɲ���F"Ń�Շ��3.��i{1�5?Ͱ�m�yM9R�%��;FE%C��̟y��2S3,ܐ���3]�:@�ьN���֬K�D��"�Lcdx�y
��e���ǖ�������3��r�Q0e���,I�_����VGmyKB.�q�ѪI/���?����\�ɧ�0�����~�/~��}�����������ڼ��/����y����pW��ɏ�٘�yne�DVv��껦"��7���b9�%l�`ۍ�d��xf07���f�f�5�;�,��A���8��"�	��:�MB.�NGS��o#^qr.��\��N����0���u�����Z�r�IN!��\��6��m�d(?v=eW<��l���Vx6�o�!g�i�^�}��4�{��E��%ĵ�*E�V߬:e�;�ܬMAl����}�����C��m�m%s�Yk�
#F:l�)sƴ�Եj�33����k����ͥd*�C����K��3g}�A��mHїw�kk[��*3���<��穕Zn��{��o��ZsȘ|�ej#��I��Y_<�-����S�0�B��_��~>	�0���c�:ۮ����Ϳ�ѫ������7~�����������ɏ~�����_�/>��<\��2�}�Y����� !P��L��ʔ��޾yc������ �ce���������K��H��_SC<�$?[7@y�-�8��X��<Ϭs33�0s��ٺ���wf��;O<�j32�D�е�m��O[��d���g���0x)�Jri��%���:nB[���ޝ���mV@s͏�Ơ�5�B�����5�s>4�ӳ���/�t��9��J%ڊ������3���_Y"�ƴ����_�Dt��Tl�&!z	�NL�)��DgB��c�SVd�x�!�@S������A�%���XS����s�������ν�=����<��tB��׏����N� �,�6��}�N�����_;���6��/����o��O������{{���-ve�rXn��X4�n���z���ev��=�Y6 �I$ō9�?��7���g�������_��������ݚ��L��OL��τ��+�d!�w,�d]��O�Є$3�_�V�5��v۝��ߘ��]�lŏy"�TTi�=Be�L��Wl%LAh	�n�$�L�
K��1>O��U ��
����-��G-ȘhS����|�ʏፇ�iH_�F~�q�@���6bz� m�x�i�9�����`z��3�µf�P�sb�!J����d2�V3�K3�"/�u!V�,F�A��%�>�(afsa��<G�$�x^۸�Ir�<�X$�o�&A�$a65�.X�@󻄔���h�^U�1�׊W�۷o���{��P'��[!�oz��y���fx��k�����1�3+�����w�|��~�';�_���,Q�zY�n�ؚ�u�<�v�Г�H3��������]�W}�H���lʿ�ǃy���#�vo_��Q'�4SlB�
m�K��C��Q���Ʀ�"\b�m��Y��gT�/2�#�!
k�%`*���Ed�%��Mԡ�Va4<�P~�r6B�\��(�$�H_A�͏�5˓��aH�P���|KZ�wa�m�,�V�sfSӟ�zF䜘��=�P�E"�0,I�]J#���%��K��K@��1fhZ�5L#_�#����钤��GNY�F��@��i!�H@�+��<Y��$����λt�^��^h����1�0�0[3^}�����׿n��+�x{m�N�p8T�t|[��'�LS}�k��ϤZ^{��Sy�SVX�]�	8�gF��>�����r�[���y��y7������h����y�װ�b�i)�T���V�tM������k���U�#�!�"��@,���f����@�[B9�IV��h��@H�k�0K��a�)���}���]!{���ꟗ������o�B�E��u�Re3�6��9�g�����	�>h�qv~��5'�Ό��".��MY�̏=f�H3t�F 4�Znּ��d Yc����Yv��6I�ɐ`���!�޼y㜎�1Z�\;&R�/�7F���{����!�Ͽ���|��?�7���ٹ3��05VAVWh�eV��f��V�؊��*��%ޣ#ׄL��9��e#l���������,�dv77���3��W18MO���-<�w͓?�RiL��� ��pc��$�X`��֛cҊ���J�+/Mr�?�@[��M�j�s�ў���c�a��u�$
�qK��&��fh�Y&f��-��Ph?�� ����G̊Xb[?��n�bL[�^be̋�5F���QX#ii�Ic��.*S#��z5���}�T��K�IPݕ�|����Dќо#��s�9��cg��d��o��\��4��K>�Mx>YWڡ����C�}������/_<d��3Ճ�ybE��P�7I�A��5���4��M���&3�\�1��~�r�+_���6�n����j|���`Y���,+�%,�5�a�1�Օ��XSi�
���\�≙�Z�
;���t��&}57����E$�1n��e
�)/�����p��Zm��i�9�i𵴒��Hl�aie���R[�X+��1��C`zi�i�˂����LK�sXs��a����B�'�X���k�Th�m�+ñ���u>f"K=Q&���	��x��o>g�}���k�������a&(+o�]�b��4�M���d��2�nύ�S��"8m�qh�A����LƸ�A�c��h��<�~��_����`)�!�+1*~��l�=��%��Xk�XH�8f\�G�1��9��q����B��f���%֌kƤ*%B����o�{6�ý�`�x��8Gň�>ۘ}��Z����m����mm1T�LÔX���O+���Y���c�^߼�{��߶��<����%���yBb,�|��6��}��0;W�w�C�Y�a��n����ILN��]	��@��u**k*ѵ�n2	,B0F�xh?@�`����-t��*�]O�:Оϙ!ѐ�S��	������6�m���ƪh�4tb�Q���/���:C�	m+e���(ږיּ�� @�k��M+^�2�3ϣF� ��T�J�|��Uc�-Sk�9�ԏ��/�ux���ڃ����!X�hj�k���J��8S�K����^�i���|�(�τi�ߵ�C�wy�΀��3AXq���������|����%//O����#/�kI���)(0	3�%�k�@���anl5��Ɣ��K,��	�s�E�P�����Zm+lf^L�ZKX�30F��x>me&���q��c�e���%��I���r�F�z2!�h�hS��J�	�����e�V�����+f\0뀕��<�]cX�17hfm�]����w����/M�^X��ᵗb���5��C�w.��z�ˇf�s�7N��W��$�j>Ͽ��V~{xx��Z��0++��{}Hņd[G���6w����Oi,�^�k;��7v����0cY�PA���m�)�ӲF�rU
"�S,�=tS��@IP���7P"!Ð>��ܳ�T��=2'2�t�M��Ycb��1�9e��!x���qt�ŨczR���'`I0���,�?f(b��it�s����{]�{�1"�\��d�I�Ƹ6��|6�#4��ڴIC�}s��C���Z�ԟ�c5~��0c����7S�׶����7�������3�{�w��E�'�L���ީ�S��a��G�����g�Hh����6\��_���F��_O������g1'X�2ڛ5梌�7,0�/F�6��d���ms�Xk0���FS�G�|�7il��-�jC;���Y��8�4C�
�0�>=�Ꙃ�e4%@6�L�(�q#�%<X��L�M��,:oy|i~Kx��%��tϠ]�ޤ1*��c��|l�0dnA���N؆CXb?ԥc�'�u�kl1��5nh����KO�/���蒅W���,����|��Ç�������s�����裏̳g�~�>�E�}���\*H*^*S^��l���MҬy���'����#��M��MGsÊ
�,�.ӂ�<Xi!:Ѳ�E�2�)x1�~��T@2�b�-̱��G�J;�V�K�,0=��ꀹ���LbT���A�!ô��4�D�Yk���zf�P�������D��GL�)+��+��Kmc McYf^��9��/�>�Dy4uN�s2��$�v�\ڰ���ڤD�z��X_$�%��A��L��a ����oȯ��F!W:=�{�3�����&i�x����o����_���>�E��|��g���F��www���b����_��|���oܰћ��5%S@E6��`mF1Z��ʄ�2�!@'F��@{�ch��枅-���/�8D��,A�Yk?g���h�iL�h���v����!V�6F�b���yKU$?Dv�-z[!�̯-t/=��S�kZ&��N��^&I��y&�5c������u��~,m�4�0C�m��s�X����������X�{�+��h±x�;>y�%�s�� r��g仛�G�}���٧�~����1#����{?��O�����ß��g����#�Y89��n�Mi�w�޹��_�~�\����'<��y�C��!�Ұ��EI����I@�c�)���ţ���d��g���o2�T�j*3c�7B���74��
��c*V�Z	3���K�٧��IڤY�2<� kL}��9T��������,ϩ��1������YLFSa9�e�e��>撴YcO�|=ԸMk�k/E��M%̘���D��(b4�����f�%Ǜ�6I3��<!i��_�l�{���|���W�r��i��9��$�_�z����W�j����[��o��o�E���"�������~���'?�����?�ݟ���XV���#��*z����?7?������}�^��c<3*D����YN�k즧�x���ZB��X&Ɔ5�A[���]�T�kC���c\l���K��6b�$@�]�܅�e�1�yj��@���<�jl9.�Z�f�z��,�ޤ4��1FC2BS��u=J��]�L_��E��'ӋP{m[�.+��滾�4o���.ee�d��:�S����˸%����!u�����rZ���-2�������A�^�=�?����_�0��_���w��]��o�_��\�����]y�;�L�++��ޯ�����_��W��������1���f���7����ן�o��?��l��z(+{'�;�߲Q����������Ǉ������?��0+��b�����$�E�"�]���[S_�+&�H� !!!a>dI�]]�K��E�WƖk��t(�5^��L1DiQ���,W�m�V �O��V<�ט��	C��E����4<I�_���������1����|����O�����/������(vc����Af!���o		v���^6���������?�'0�a�J���Иɒ�j�r�AA��	������;V+�)h����D�\3R�&$$$,&1�����#Z4Ca����2!�v+s&bm��׷�?�"	��s��{M=�/K�z�%�g[�.�ž�C��(���Q~���mט��L���%���+�q�g¦u]ly˧���^�+��o~���~���2�������σ�<av	�F�b��;�2�tb�`'ȮEF{�0Up\Ch���z}���蓼݆1
��6m��b�O���c���p�m�ֶKH�Pc8�.a����b\׵����4Y{�6v�R�LK��s�i}���u���71�^�n�����eЊ���=���XEtS��G.	_Vf���@캽1:aVZk�M��"�*�����U�"�ٳg�e������2&av$��x����� �.�x�FW����kA� ���b����ʘ���t-dY�2��				K"ͯb��2餅1��1i^�W���>0�#FR!6����u�]֘�{6r]��F=���)�S������&���}��=Vdi�z ��1cH���0��g��o����QF"�.�4�fr 
����	r��؉�)�պh)���k�,�~p�H$WBBBB���C��7��6[R!�&hGd@�,S�g��j�<5*�DU[~k�Kx�"^GH��X�Nc�}y�E�i��8NH�5��!���6|	�o9½��.w"�.�0��Zb�5��K�%�Z6�Yv](s=ۺ�^�@sM�뚟��x͸�������� HdY?�Dv�Ro,�>[���&��,�"���9��^Ҏh�Xi]����!Ҭ��-r̚ɲ%�|SI�)X��eڋ'�]a�H����j�eg���P6�λ
.�Ͳe����3]����e�Kv��l�eӮ����	�#	�			s!y�^?�M�Km �o��b#�+�Bo���6�)Kx�al������}�M��Y����R}!���[�}��6�BQj��l2�ZH�K~{�a�ڿ��U�d��0�5����&���)�}}��	ihT�de��׆�J�3h!��������Yk����D�\�� ��Z��Hu��T�	s��M0�_#�5%�b$��Jn��3UQ�Wi�׭������BV�]kW�,9�!�B�i�}dٜ�X�zS�D䲑��XI؄�%r2�FWB�=<<�����;���όav�F{R�i�F�lhp��~��B�18�Mϔ�.)��v�wژ}�IX��#)q�J����8K��|�Юsģ�) $ȵ���h�h���χ F����	Av���#�u1�BԮ�b��/�`�c~S��5��`����ϰ{̽sc���e�:/i���{��+{�Z[��[w�>��De@�/�o�٘�n'疹}���������Ka�������������������������p�1��<���4�3�/�`KHHHHHHHHH�G������"͋					k�x���X�~�(~K!fd�+weMHHHHHHHHHHHHH�@R�'$���\�������^�y���D�]!��f1�����������+�r<!!!!!!!!!!!�z��e&�u]W����K�ٌh#�>D$Y8!!!!!!!!!!!��Fȓ4=̚ץ3�V�t�YBBBBBBBBBB@e�b�@�8�oBB�4/&$$$$�͵�-b�d� f
H�YBBBBBBBBBBBBB�80�щ$HHHHHHHHX��{�yRL��&RHƕ#	�																								��`��M�ϒ3��7��{/����!��Z�3�,����LKB9@p����%8�����L���N0C7i�g_���s���a�)�y����K�����F�á����� �m�����C�b�)V���p����D[b�ϙkk��ZK��!k��~�+�C�!u�<���MK��Ǥ����3����tb2w"}3���c�Xk�i�R��ት�@����ʂf��Z�X�:��v�D�bɀ��Q;����N�T~�9�ϓ�u<Ͽ��ޚ����E$������O����zCms"� �X� ;f�)�h�Yv�@��Z�&���7�1*�cT�"X�.c#�����\k#
]�2i�s��3?Y�^9b�Md��!�����*T�I��
�)ʋd�%�Vі��+/�<YĄv?[�~����9x�`���B���1�]�����tވQnў�Y{U����ރ%xXeB����<�1�1�+_~���С�Hȳ2��qM�E�w!��S����Z��d�ֶjss��,1n�ƴ1S!Ϻ.�����B�y�� �	9S��S�b秽!��21! ��Qt��"�c\�P�}	%m2��h^Ri�ڬmٿf�'6�;?�|΀�8gz�@<�XF ׎,[����,�(F�K���c<S`���[Bve�Ӑ<b4(Y��j�h�M��x#��K�0� ec��F�ŭ�J(��0�mV�M�G�� �bA��μf��!�l�m�$�ě�5l�&��B�z���v��]�}n��g����(����
M9��xjK��^���0*���5�MRt	C5�b_���  ��IDATӲX��ŷ�'�uj�uk^�4��ܩ)�gi]�֘4F0׏�s�d�Z��P,��y�1��X@�)�0���QƆd!�d�O�i��!y�������5ds�fm��}f�k�аp����c[�b�O{��5����M�gԛ���&гG��
M#vZC3X$�\�c׺��~�ַ��*S7�1ȡY��0�<F��d�6�c�%2c��G��t��>t�	�ˌ �����i�2X�s+��%�5����.k��a���E1�_	2�^P���,Ry9�r���i¯�M����vO�1Kf+F814�0Ȃ�cq��7��Q������	�5�<]���Z�oμ���飍XǺ6����#���0c�B2�N��^X@�"&i8T��z
�VF�LlYRs�c����kZ��g2 ���h��l�p��t.�6r�nc��b[������M�diO����Q�מ��u�0e7�vY"����i���٭�4��C����F٫��XH��4�s�nnn��K�!!&���pp�sظ��f�{�`yWe+c,w��<F�]�܈q�D�W;6���_{~,a�i	�ʏ�M��5z(/1�XB:ː F�eL�D��DB�}��5���6������5de�7nc�e�)o!���4,b]�$ǵ-\Y���L/�Z�3�A��=:��q�f�5�1����y�,!s�e�Jd����ƖLٍ��Ʈ����gT��I�,1�3�`k�����A=���/�sv"�.@�X���_?��ǄW
�Fo����JJ0�fm��.����D�f�%6Ī؏�]���,a��R���8���E �7۬�PR�9�J�!J��Siix@�>�M�y����C�IB~�Y�k]h��r�v��e�6aƂv�$�^����@1�sH�����,�MbfL���ݵ#F��ΎM��a6��@�ޚy\�D�ċm����}��������lԸ������g� ���d#/��@�>�S:c���3ˮWqѕ��V�)E=X�0�g@ĨdF��F�d�LL��Eho��H�-1�Y�>;&�0����m�����h��x�%�6��r6?)��S��I��u}�Hd"�];a����(b$����IS.[3Y�|>�Wxl`z�#`�a������w����ϴ����9ƀ-s��	o��_8�L��1U�/�"av^�~�-�v����+՗/_�-_=3Ɨ��7uk���7�f�cnEޜu��8tQ�$�
OR{��f��؈}mRM[хX,A�6U ���M�!@�5���!`�I�6F� �l,b$�Qh���<���e��A���֬���LYb��fg5��>F��~����/�����V���4�̱�M1�"d��3#��
������yM�=H�X�2��p�u�t�n��� }��noo���>��w�q/�}�("f��?���{��ܩ|���ٻ�^W��N�[g�s_����BP��1�6��x�iz�@�i�_��� �I� e�`�k�؆#6�,Y�%\]�s���~h=�떊�*��b���r�Ū�U�b����e����_7ј;�s�h�<1q�?���Y7�������}`�>�գ��a�A@�������<TY��>�=P����y9U`�x��Ny1�Z���ֺ������s�3LU�Уz��X�PU�s�q|��F9Ǳ��>��F^�;��M�;���pj��4zz�8��6k<�Ы�>���b�FO��_�|V�.��12�;���`����`�gTU|U��\U���:2�*K���n��1b�EY�£�}��G��#8���7ӊB��:��w��on�������?��?�����w6�	�����1��k̖w�%󳶓XK�����'�Fo��_�8�vB�: Xm�y���\rP)0{��w|k\����m��
�}���=��rq��a=��	GoU�������f��H�vWy�y�����ؠg�G�_{���*�������h.0;���JU�Ī+�{/L�X�K��Y�I�^U�A��4��~�=��7_=����U��{�����*?�˼��i�z���@�g����G��Y5�K�z����u܎gn3�Y���̢�(������y�M�Y�"@��������?��?��������pu�ٟ���7���7��|����G?����_~ڸv�����=�����o��o����}ӮfT���?��[�aV}(z��j�jz�'8F~��l/*~H�#,�:���ֶ�G�e��KL�1�>ŕ̻��K�0}0�;��}g��V�ߩ���	���e���9���<;O=�Ξ���AU@׻�z�>�?����W{���q�S���L�g�m� ��U5���K���'�F�VY��C��-8����i�g���q�1LZbm���@z�E++.�.���^e�@���=F���W��-[�g�~�w�������U��#�W}����m�Z�!e�� �sƶ׶�M/��x-³x=����o�f���{����������0E��t{���������V�������{������O?������ۿ�,���
������_�ɟ������}��}����e�U,O�wc��	�o~�7����o��'Nfǰ�~�-VfnHsW����JePR5�S��mF�<��
��j���ԣ�R��1f�ߧ:���2:0[�ɾK�Z\�?=fz*����S�w��y����һ�+T~^*�?�����_�/�:	���O��ӊ���k���^�U�=z�ѿ	��������G����魵J�G���ܥ���Df��Ue�MUV�2�9�齘md@Wy�����ha�y�}*����T���^�6�3�����q�&T]��k�q�!�ܷ��3�3��DS�Q�����~�u�f�Wu�o}k��<�����ϋ�3`�����s������>���_�<�;��;ݡ�UfO�W�����E�b!���������ܨ���X11��B+8�6��&���j��W%�TJT<���=dzk�z�� �rz�Ot�Y��oT%���r\�z��%O����\x�s`Yu�fo��;��*�g���{�g������>F}º�dm��[YeW1L�j��D^���W�k��9�l��ܡH����R�I�ʋ2z�x��lZ��ｪ��^#O/��U}��.B����w�GVx��<��3�ޖ$.50�jV���г<�.��Uu.�T��1���$c�r\�³���vzٲV��!E��|d7�����0��v�lYl��t��c���_����˿����W��z�������#��=�Ql���i�L,�}��O{?� f}��ȫ��1W�M�ꪋs�7���K�w��?�rz��:���.5�Ua���JK��۵���:��$z����+U����Not�1�U����Gf��{U}�UXUͯ�K�.>����2�>Ĺ�0�s�c�Amմz������B�^����hz�b�se���x���sNadeQ���'��5�*��E��������{���1��\�xFN�24l����K���}T�&���r^㵶�4��x���篇���N�#n��Ͼо����;���o}�+_���������?�����,�y5�.��+1�J��x-¸L<s�r�
������J�jz����}ٍ�!��+�zU]Qy�/��0�W�
0��^����9��.�����̖Nc����'F+�J�|W6��3Le�G�5^Y�'\�x*�w�˼�J����M�TS�w<��qt[y�[�C�+k*Û�c�ʓ�=DUnU�s�Ǔ�?W=*/����r�(�a�����z��G7)ڣ��*�	k�zé��p�f=��W��c��e5��@OHv��_m&��,��;/�k�ڦ��.�&ߟ�j�����=��AfSO�ݸ�ҽX`=��
̫P�q�?R�x.K�>�h�ЬG��'.50�����:cn܇���X2\����Yr��>�M<�<І���[�#�wz�x�*Lz����'�N��e0��U����ޜ�u�*�V�\k�̬10#O�V^�>�[���U*�5�©����՟��UL��}U*��J#?ad��Z�w=F�����ؿUUk��`��%T� �s�U������^�/>Z���%㪺��%�����6縠�r9����M������B�mf�X�",�}E�M���.�����v�Ր��x-��z��gz������.®|~��2 ˲�<(mWJfmy��jt��kmW/�̎)A�u���y:�Iѵf�*���-=�s�_��o_`�3?k<ح�\UUT�\����{䕧K���y김'ǵO��Њ��j<k<�ޫw�:�c��5nw�'FGV���J�g�鴶M�b����1����WE�Xz��t��>;��ӹ�����n�w�.��U�[*â*����y���Ze��;z��P��m�U��ثgTN�r���G~FWn�:�v�s�#/L��8pn\��U6�ގg�8�&c�Ӑ�����K�?E�M0Ff�xO�f/^�X�ϸ��,h.�ލ/p���^5��Z<?�j��g?{��}n��r%�F�@�^����1����r��+.�����Nr��+��x��jz�ۦf|�]Y�_e�2��^����v�p����'��W:e������M�v^��Tu�X�o�����c�v�d{�5Ξc�<��5��+ї|�-ӑ��;�9�?����?:?�f�w��|���Vϟ�J������Ԯ����x���^K����۪c��a�Di�x��={�c�C��}�)��]���}b�w����O�ڎ������z�u��I�-�S��wl:�w�v==7��E�2=ϖ�2�������h��io���Uf�j�6,�<B��,�{��n>��lVbۉ]��4���l_EH������%y}�5f���'/.�ȓ KT���:=���G�)�ӣ������C�U��N�q��p��y꽰a:�m�=d���v�����o��c�鮓j�W�v:3�����Jy�{�	�s���S5��w̮m��£gzK�j?&���m���qm�Un{U����'����^p:���K��7�ڏ�+��%�m�}wW��.ި
Jz?{k	�Fl�ob`V5�ދ�*��oZ��v�V��ܶ�7����oo��:�}�20��#��6㹨0�۶���͡'�0>=�Y���U}�6�v�����Y�<��+kFO��s�S]�}�����S�j�;�w�������y�џ�*�|b�jz�X'�|�N�U���ϛ�}n;�>>&�9d<=�ˡ���c�cvA=��Ls�ɉ���|�~�OϽ甁پ�mS��X{����k�(�5O=aʱ�ٶ����s���Wv��Kυ�y�m���=����{�����4���c�ꠤG�}\e�U9��y���ݶ����c��}���G�k�Ե�f������c��޳dZ���s�f&y\g�Xq��榙��aY�-!0�Ю��)��XYq�}�eS
YuAZ��\��_Z��}[����k���N��,�� ��l�jz�����UO�neU_��;r=�q�����DW�:^r�k�s����Ǜ|�r�u7�}�s�\�F��m��v��%��]�;��Ρ'h��j�:@�~�.���ۖ��*SK��m�>7�xyih�k�Nu��1������*N��b����cǵm�c��"H��#��7�ڲg�*�mj�==�XR�p�r:���g���@��"��Ns:���|�q˾�ɩ[�����K��a�Yd,��d_e�x��/����o24[J`��܂���6���Ϋ�~��?��F}�d��`�*O��~^�}fz�W�*���֥�<�4����q�<��Ϋòʃ�W��5�X�:��q-Y����F~Ϯ�������q���}�߾ionI��}#N�T�|��]N�}�m[�K��m�N�����;�������C�S�u��ڞ�V�ڇY�~�gW�����Uy^��w�ھ�+��z�md�۾���S�y�M�������r�]�W��}F��J>�Wf��U���L��=��u�+���4�������2�+�*�Ӯ����/�7yYVs%�ث������rqda�\棧�c�<�����,�y�xz��'+>�Y�xN5�
#O�/9ٳt:�W�'+=���O��<�Gve�0=�s�����쩞�u���	�ND|n��: [2�S�~_o�����Ss�<�Q5�5sV��=�~�ws�����i�{}mǁK�˾��ږA�1�ҰhW��&w��T6�;�w��c�C��ޜ��s�q��l[N�XV���㘼�M0n���})��:���C{ 1]��61�[�6�8��CKt��q�Wg�>��6�813z9U�����Y�kUӫ���ڛ<���NUaJ�5V6~�B�ϖ���+�G�<�{�j/]�ӓ=sW�U���_���F�Tl;ѿd;?60���`Β+p���>��BO_K�FV����~�����u���k���t����V����P��.Zz�uh�ܪ�>�9��T��}U�{;���KN�W�ЭZwk�z�5�7ͽ�2����L���4V�S���>�����G��h��F����3�S�s��G��8�����Զk�6�i���ss��!�P��e�.���'	�q�w;�(����D����k�{ [=�5M�'�������M3����y���`�'�G���E�����nS=����KOx�p�ｪ����[��e>�����,N�7Xzr������l.�n'��m������2X��\ 4}|�0�gZm�S��5=�w;?���.Ua�9N��f��\������AB�:>d�sL0S��RTgTM��b��zT�˖�vq�w��������w�gf�1�)���P����mӫ\?���U��������l��]OӐ+�O�z��u�}m�߉s��6$;�pI`�a��"�l;��[�	h��1?�v����N��4Up��֚~�U;�$ݡ�T���^��uZ\)�%���K�^�Um1̥N�Ǜ���\왧�~�NŴ����Wd��U�������z����7��s�\�R}B�B�2����pc�4z�����澾xz�9��k��]�<Յ���c��%�{�h϶�m�8��:�2Zbz�`[��Oo_̱�3w�9߿t�W�F��գ�c����������]b<�G̍���.�[r2z��~��/�٧wz#��ܦ�}z>t�<m�����7XO(Z�?8���)�)�k�Ǆާ��J;�߶�9չ�}���Mò���lZa���m���[��Y����� �ʈ�Wܲ��~�M�O�l���RB��_�k�� �R�a��<�
�5�m�7Ti�<��x�A�<U�z����'�F�a=*���C��J�'8F�VMr�|�����{B�b<�Í>1�o��--Y��^]}�r��w�	ϊe޻,{��^KO*;�S�`{ðc�ٶ|��r��>9|��GkL�;��-�|����W�0��:DŅǎ�����c����W���:N����{_����gĸv}�j?_�*�;t<�\pt��������(����&^��|.C��Pk�MVN/������}��Y��p.KsB��Kv��˵ضn�����%��%����N�h�#G��   ������~ZE�V��vv�@�^f      \�6L�V���n�z�      X���l�,��}g�      X�m}�NC��.~f      �]e���saY�[־�3      �.�gϞmnmp��i`��k�q�      g���z�>�      �xs!�4,��a6�4;����
̞��!eys�`N;��&�s+"�P     �k7�����yLV���q�����nnoo_7_V�-qU��1ڶ0���4�l�      ��l%�6����B���g���f      �M���W�e����[����lZ�����m)�      CM�%m`�AY�L�\���2LӇ      �ò�l.LkeH67�
3      .Fx������-*��>*̶g�m��m��     ��hí�28k��Ҿ�C² 0     `�i6����L+��~�X`     ��h�����=<<ln�|�g�Y����s��R�B��c�F	a�      �Y�E�}��}em�2�Lc���>�B��X�ww5     @++�▕e!�2{뭷6�Yh1Lh�p�Z޲J-���      pv�M�Y�ʀ-O�H�3      �.ò�,�ǻ��i!����N	�      8���ۜ6(�V��z�.3      �n�cb=�f�8��:��     �
��i6}<חY����     ���e���[�]����nn\�f      �]�dy�0��2,�&��{�K`     �P�P++��[cs�W�fYe6�f{<-���B[���>�io��c�     \��b,r������Y1���߷���������6n�z���9޼�0������uU�����      �d_�2�o�)	�      8���m�/_����Y>n��V�-%0     ����}.�asڶ���     0L[	6WM�/����c�      8���={������|�:�F`     ������#L�����ǭ}��MC5}�     p2�
�*�x�!Y�f�{_�NE`     �Ye�X�esUbmuٜC��ZW�=-��i[�      ��\�dm�7�^��y����碪�m�1���m��-ޗ������9�vU�      籫���2 �������M�5��u���     �՘�8�<cT��!Z;��{��     pv�����l�q��C² 0     `5��k. �����l:��     �����Ŷ�l[�fK	�      X�}�2�{>�2�      iW��m%Y�ܴ�,�����     �U��,ði�vhXf����ڶ2Y�      �h.[y||����,�o�{�����i����]f�������9      �iï6�zxx؄a���2L��Sd6����m�����     pv��b�_ٶ⥹�iP`     �*̅esAZjC�cZ�     �sUe����>���!f      �]�mkZq��f�T�	�      8�������V�M�5}�     p��f�����}����d     ��M��j�gϞ�V�Z]fŎI/     �MV�M3�����L���m����ö613���vE������o��,r     ��Q�Z,����<<<�|��Ǜ���|-���%���h�q�6ј�Mܞ��w^�7      �����B�dY��AX<�M���)õ%f      �ܴ��i`���"��[�J�6����	˂�     ����M_�7��Bk���>k	�      g�^m_dmS�mȖ�hm�Y{���     ��� +C�V`m��aYܲ��̢y�v��8��{	�      8�ĶZ�&�f��m�`���y�%0     ��5�؆]QQ�����,+���v9$4�     prۚdL�c��Y�G3��e�m�Y�/�Y���C۰l;�ko!M      浡V޷�c�|b����[�f�Z��-^�-oϟ?����[��\U`��`���0�{      ��Xmh"���+��� m�ϴ}���n�6{�wޮ*0     `����7����ʲl�Q��      \�]�c�}ۄ�/���K�      X����em 6�L�44[J`     ��M�^��}J3      V'+ɲ��Т
-�)��&;$h�     pv~�M.�㼵�5�0�E�v{{�y>�u\B`     �*l뫬�,��򬽅x}��
̞����     �"�zxxx~��]XgYq��gK]U`څ�m�M��k����CP     �K��L���e!��m�4�������f      �O6����E��g�m ���-�|�rs��^3      V��2@�0���Y�������#0[�z��     ���6�؆k�e��R3      V!C����da���������~�|��������     pvm@���40Km?g�z�f9L4�(0     ��m�,�7�a2\����{	�      X�6����.k�2���>�Ͷ�m��:-M"�     �?��G�?���V������r���R�mX֖��˵���MW6     ��j��B�O��E�c�\>?�2k�j�|���Oܞ�}�;_3      N�-<j��V��k�f      ��ž�*���|-�l�3��Y/�      '7�0�.�2˿��?�m#0     `�����2΅b�Zۏ��p��i3      �jC�i�f��rع�64�$#      �6��V!�ʹ���     ���U�V��m[�vL%�63      Nn��lI�����"<�u���+!S��T.�?E�     ��"����׹����&o����pw���������������/_�������8�����o�Λ��CuY      �,Xj��",�0,�����*
�f      �]V�e�Yh�|V��kQY���,,m�%0     `ڰ�˦�g��V������L`     �ٵ�e���m(��f�kǄeA`     ��e������uӋm��\>n�b�V�-%0     ���j��)ƶ��6�k��=<<�~���     ����+�f�&�Ҭ���v��f      �]��XT�e�Yf��s���hy�aY۴c/�ٌ�Bl;��R�k�$����     xS�e*m���g�5���|�V�e?gK��Y�iY_g�A     �5�e)���ڰ��2L�p,C�x���.󜗽�!0     ��`iZ����M3      �n.0�>�Ҵ�l��0M`     �*D@��68k��4Ͷ5��C`     ��M�b�7leӌ3      V���ۮ@-�Y�	�      X�i���݆`����     pv��6{||�ڏY{��
̦���V��	     pMڜe��mzq�c[y���f=}�M]U`��ٳW��2�\���޿y����fK:�     �_L����a�>r�9L�Ѵ�Xަ��O��V�\U`     �:e(�AY<� ,nmxv�V f      �]�GYdyˊ�΢�,óJ3      V%B��������M@��fm�Y�f      �]�'Yh���+	�      8��$���������իW�����8�j�j3      ή�����>²�e����U�     pvY9aXgُY�]�%�Y�S�      �kM0��*���?~��[om�|=+�Z��ӿ���S,��X.��,���e�m�smGt�r{��     x��Gm�ϷAX���-�9Kd'��dZ6�2X{��e��e�Id���Pi     �\�eSj�2$k�3����     ���
���Ucق_V�ŭm���     ��k��jðx.+̦�gUf      �BۯY>��w6�خ�f      ��\��6�8�.Ӈ      o�6˾̶=�}�U�     pv�=<<���[>��m�m��     pvQ56�l[u�.�{z]U`�� _M;���u�wwW�Z     �+��3٤bܷUe��2��,����,^���9��l�60     �<��`m�6}�}��z���������     ��ڪ�0�,�`<�      CMC�ie�	�      s�6X�>>$x�     p1��c��f      �����Uaa�߳C�#0     `�6,{xx��/i�q.(��B`     ��e �V�eh�Ϟ=+��
�jS�\��\O;�KSQ     �7UV���If.q��,o�ks�K�|�����l�\q�v�Bo��i2���s��(     ���,%�67������0�����'B��[��-n��ۢ����z�K`     ��e��6����J�m-�mk���     ���f���6���i�>�m�K�      8��n��Ҭ���
�}f      �E��M.Nom_fهY��t�K	�      �����M/��m��0     �b�}��
���]v�      g3�0���b��5�87�^W�m[�=�	     @�]�a�e`vL�K]]`�e�ػ�3������7�>��ի�Oλ��[�      ?#���J,s���,�� mZQ6��0��,!��t��0     ��4��&î���ٖ��B��q�zn�      '��ϱ���ٴ���<k�ȶ��3      Nn��\Ya���ö��5�x�      Cm��>����=y�v�5Ӗ�     pr�B�Uem5�\��g�YEh&0     ���ʰ��x�������ns�gm�m���
3      V/�Ǧ�W�U��#$�a�>n��b�V�	�      X�i�5W1�aYg�is��8�M3�����qۂ��#�՜     p�6�sKT�e�Y��걬0�`,2�6T�곸���i����v��Y�c�K     �7�\X�a��4�֏Y1Mߛ�-%0     ��2������ߴ��j3      Nn[uY��⮰�����5��     ������l.,k��lSm�K	�      X�c�^�     �J� k�	�m�cs�g=��%0     ��}��!X�?{�l�x���4X���&����Z3      N��¬��{
W����.���7���?3�S�<     �K�IV�E��bm��h�ʴ�~:l��
̞��O�7�«
ж%��2     ��J6�"4�L%���g���.�0�"����     �u�VIv3      �i[�kC�C�/�ai�1	�      �²	���lװm@V�5��     ��k��~�Y�i�Y{߾>�Re&0     `����,+��dl���(kóC	�      nW�d����]�a     �Ei�d�����v5�Xя��� ����	     �����XܢIƞ���R;Ξ�L]U`����ڐkI��+��������������?~��tE�uR����as�      xS��Gm���Kh�2k��|>�#����}�e&�y���o���Uf      �S"��W�T�)	�      �m�o�R_eY16��*8�     pVmuYޢi�6P;e���     ���.��R���)�      8�m�X+�;u?f3      ΪĢ)Ƹ�ߧ�,K3      ��6�2 �[�f#�      8�lZ1M�AY[a6}�)\U`��@���S�w	     �?�zM������������x=�����.n�疸��     �u�`-��%2hk�z�!0     ��c�B��5�*3      �n��b�wg��3;��3�      ��Sa֪�4�     �m6�e���k��@�F`     �*<{�lz�}��l�      g�Uc�ŭ�����4�8G`     �ٵa�\���a+��f�������O�^�8      �A�,!r�x�6͘υ|.��������u��t{�;m�Y�,��)     ��"c���߄^|eaR�/���,>����eڠ���     ���B���}-ó�2�&0     �,��[M��a�q{?giWYA`     �Yeh6��.���:,3      ��ʱ˲_���&CeѧY6��O�i����L`     ��dh!Yhò�V��.�a!0     `��l����~��RU��     0�\e)�Ȳ���=m�)��f�z������7      ׬���U�����ׯgX�q��Gܲ���f'�++²cJ     �$m�!X�]�����l.Sɾ�noo7�K�V����ŋ9�z�E`     �Pm�XV�E����oo����Ȧ�i�8%0     ��"$�J���ji`�p�0     `��@k�xxMC�v�|m��!f      5�ES�y��̲���*����l���3      �&C�i`vww���,o�Z��e�>͖�     �*��4m���>Sa     ��M�6����(����T�={���LǑ���cv�      g��Y�e��}�6�����Y�i*yLI     �5���2��
����3{��������=���2�����q��tؗ��&0+"@     ���?2��
�x�6�ؾg��
3      �.����V�e@�6Ÿ�I�C�4�      �AY�Mïi�fU�f3      ήɦaY[a�em��\��K`     �jm�Ҵ�L��      \���={��e%ٶ��~�
�3      �.����׷���Y�]T�     p��ʱ��ء�c=�*0{Z�w?����/�     ��4������y.�ۊ�h�1_��� -�x��Ͽ�;oW��S��      �����V���s���UiK]]`     �xsAֶ�kd     �M�6,�ʲ]�amu�)�      8�6�	��&�/�S�     �jKö�f      �\O�57̩�/3      Nn[�gϞ���e*�      �xs��e`�����l��c�v��s     \�m�d���������M�Y;|�x[e���F`�!C�����������B<     `�iuY(��]"si�x�f�8�q��j)t�     pvs���.C�iaS�h��1%0     �b�g�e`�A�Ұ,�      X�l�1o�w[aֆe3      .֮�+�<�׶�U�3      .ֶ�6(˿�`�٢�lih&0     ���5�8��=mX�?<<,���     �՘6�8ɢ�,n9\�_�}�e����څ:W�wH�q      ���<f����X[]vLXf���������ŋ��g��׾w[u      �����o�S�<%�U�f+��������{34�gip&0     `5��cm�\���}��     pvٚ�4���fa�|�f      �ݶʲ|-ͅfs�-!0     ���,oaZ=���\e��eA`     �����*�60˾��a     ��k+����Pl���P3      V%ð���OT��f�4Řf      �´jlZ]��W�u�V�7}     �ym�c�[����yxx�y����ʲ����n���b�gϞm���xb�|���l���L`     p��	ƶ�)2��BjmN��O���4��     pv�euX�a��      8�ɢJ,C��0�:EK�3      �.�+�[�U�Դi�^3      VaW�X[M�ش
�}m)�      ���b�-�oe�vHH��     �
����[�d�-k�?�YF�      g�V�M��0�\����J��
̞�}�����fk���}��2?     �k0��X�^�'Yfm6����8�p����w��-0��g"OK��L�'ƕ��      vks�i�2����~f�6߉���-�{xxx��RW�     �>��%�+d�gɰI`     �P��[�&�U�U�     pr���,����4$[Z]��     ��k���e��6�j���J;��     �a�fa�MM�Ц��q�0     �"d�����	��>Oóm�emh�>�44�     pr�­i@6Wi6̦�ٱ�3^U`���^U�g95W�׺����     �	s!X��i�I�c]U���}mGrU�Tpn��k/^��y��o      �M]m���ٳ׹M���޾.B�|%�s��,ks�i��Uf      0%0     �	�      �j3      ���     ��&0     �	�      �j3      ���f?��O^?�ԧ>���     8����M63�kB<���p���������7��{r�x|{{��q����w�o���      8�m�Lmȕ��4X��sL���     �����ٳg�걸�Ug�8^?�      ôa����2�{=^;Ew[3      ��k~1e�ٶ����߬��     �!2k�����"�f����q����     �a��Y�"˰��.�9�      C��2�ڪ�68k��m�=��     ���V���0��ﲻ��x�����      8��B�by��&�^y��YۯYh��Ϭ�|r�K\u`     �b��X�\��M1F0�|>+���-C���%f      �\�YӐ,���������m�1�n�3���>�f      ���i��g`����|�48[J`     ��/YaQ]�f�|h�Ŧf��sfmUZ/�      C�U���}�-y�1f      ��0���e6�k�a���l[�6����     �!�
���M)f���m��}��	˂�     ��� +�-mX�}�e�a�t����v�ٖ���li'o      o[Fӆ_�*�vU���	���f�����mss�MM     �k�����qT�E������~���x�b��;�ssww����6kó|��H[B`     �E�ପXI`     �Ej�]M6�#0     �� 0     �jePvHh&0     �bD�e�Ȧ�/!0     �eE١���     �7�>�      � �"Q����xs{{�:������[o�      \�����U�[d*Ϟ=������?<<�~n�޼���,���������     �!�B�]Ä6H��lkjqZ�t�      '7�_�m�/��´zl����      8���>C��V���|��f      1~�U�M�m�"0     `�i_d���k��ؾʶ�     pr����4�V���     ����e�M�+�PL`     �iZa6��b�p�ʦ���*0{Z��mRe}�����~.�Ls+<|���7���     ����?6�X2is�VV�E��������-����߼~ww�Q�]U`�bA�XX��6�VP��     �eh6W�4.�e��{�0*GX���e��$������dam+����p��˗æu�vA�W�̭��ֳ�z���b�Sk���M��5���?ꂽK]�K WL�Gձ��K�xFO�J�z��{�bz�Z�9t<��f�����c�xG;�;��f�gf������,&�e��܅��^�ط�m�\����c�}��6_Kο��;�u~�:�s���+����M ��M�b��c�W�^mnYq���������3��vU�ٶpkߊmW��63�e�'� ��u��7ӹ�����w~k�f�T�m����u��i�C�LX�o�f`�d�\>������bdYm��ϟ�8�+��-0{��m�  �	�~ܻ�o���\��N����J8�s��p����lK~LC����>���h9��E+|1L�co���湨6��"@�
����a6�i��jSȥ��]�ʦE  �o�Ϟ��o�Z�j�x�J�ks��`����VX�r�x���c��C����Yv�*���갨��+�r,ߗ�����ۛa������?��5�8�ٳg���e&�ai��m��N�I% �.�d����xM\���kXO?��Pl߾��6��8�r��{�}(�p٬b[a��s�d?eYY�����~��l�����������U۶eoG��`,ö�,�  �.v��o��s���w�s��xS��B�Kˎ�SY�}�͵���;�����}���|�37��ηz���h�qiX��es7  �s8� ���Y�vÛ�M��M����i�ٜɲ����Ŭ<�������Ǭ�<�я~�	Т���~��n>�������wU�����o|�K_������3���(���#��2ь�?���?�p��bY��}<?�>���ϒ���5��U�c;�m�䃝鼟zۨ�"������H��ݳ�rh��o�]�ۧ>u��+�����~��ƾ�p����y��V��~��mx�|�c�+��J������'�q�2r9U�k��fF/�/�S��[:�c�Vi���|����W_�=z������%�d�>ã��]=w�8��;�G�>��F<ۖ�����m�r?|�|r.��G�x��,�s��Xd,�8r����w����gH��%���F�y�ʲ����W~�W���~����M��
�~�~돞����?����������߼��{�(뛓+-�� ,�����|�[ߺ�����Yɱ�bFj��/6�CnKN��"(�f�B��62l8f9M��'	���\�֦��Tn�=�9�8�|����������z��3��b_�O|���{�>�Y�U�ZOB�#ynP�����>���C�?�F���?��Oϸޤ�ޱ�O����hk�F�l:~��7Q��W������7k\�|�{m����y�?ǽ�+z����<�^1L��y��G����)�*?{�,�}�Y�u��p�x�����`�o���C�l���s�=*Wdȕ�cۏ¦�^����W��)�F��g?��M�K�'^�J���f��~���~�n~��~�ז��Uf!B����_����������������������|�+1<-��O��>����o~�棏>�t(��G�ZȄ37�XyU'}{����r��Y�m�z�w�A�ҝ���<����Y����j�?l+��'�G��V��읧]����sVM�R�r;8e`62��Wl�='�F��m���谺�����T9G���>��'�G�9ί��W������깨��;�j[�]�'OG^�Xuҳ���sBw��]��{_���Ɠ�U�w=�yo��������㍪�q�ga:�\n�����c���5��z��	�ϭ1����g_��m�w>�״�E20�l�K_��͗������_���z����;�����˗�?�<��zگ�|�}�������?��?��?�������,}��_��޾��������k_���}���������|�	�2�Ǉ$�����Ɠ��h�a���i���j�m3_�TW�w��DKT-9�>r���(�*��� �,Gx�-Ϲ��j���UUU��S\�-��+�*�go~�x�NpTmk����{�W��^0��c�5WY�������x�w�>�'����No�ʋ2������lmz���c�<�Oe8>R�q[�E�U���e����Y��p�?.��r]��5�W�F;�w�!�Y��Ez���q���F���h��(!/0ɋ���l��_���o��o�������YҬ�1�60;֯����|���o�����w_�M+5²\�m`�heif�O��'	��N�Ez̉�C�?��Ke�z��!_ʻ���=y�O��J��\Fy �:��c��5�am!�>y5U����7��?=F��Z���t���s�T]�����os���O��M6�R�wyV-�����oڪy��;���R9�������T��}z�?u���z���>3����,�H�l�q[h�d�U���l�.yy��>�]DQ�UM��xղ��,/L���8���h�/^�f���/���² 0;�����l33S�v%�<!��Z��J��F�{eU'��v0�����s�>i�;O�,�r9U��R�ӭ��emF�8��j��PyU����>/yu�(����=�U�:�%'G����z���5����x�����pcmFo+��=��Y��N}�cU��K��F�S��ˠG��Ttk���[}4:0���9�[�oՑ�6�No�wZ�w̡�`.��m��O.t?��}��7���s���?��z����y!W���T��򊿳���0���>�����@�#<�����&��$Vdi��n���@T:�U�U*d��ڜ�¬]�N���p�;εW���~]�V��V����*0���U�lQ��&Z{TU@���{�g+?�������G��p5�}<U��Z�wQ�ʦ����ڎ[��m \�Ev�̲k��+u.��/ǵ�m��"�5���󴫚�꘺*��q������FWUMk�y���r���*��O����������3� ��?������짯t3����r3��`��߾���?����ܘz�w�0U����:e�0�����_>��ʒ�=˾j�*�^�ճn�����9�lF�Je85�oe��ܶ27�#��J����C�ɎQ��X�U]�]�-Q�V���=��i=�Y�*�g�/8y���׸�FW;U��,TO.�V*.4\2�}ӫ<��Ry��s���q{�գ�{��8b�����pɁY�Iߪ�9z�3��J{�ŝ����UVH
���U1L��z�Su�j�Y8t+C��z�P����¶yI�^�xq��o~���?�t}�J$���<�
�LT�e;�����;Ｓy��2�<���ۣO�-�ޮ�f��SU'k׸L��������
��U��[�	��0�GCO��?�n��^︪>W�����p���[��ǡ�l�G���q� zOjW�#��{]�1���U��ȓ������J�wq��z����9>�=Ffk�RZ�Y�'�+�#B�����_���DL���m�^���Y�ʰ�j�����r�wڮm�jZ����{�ő�^]�;L�"G���>�h�}�{߻�я~�y.��<G4�#�Af�|�
�J�x����ʓ�=.��ۚÛ]!Ne�F�Q�B��+�+�����-�\:�k��{Ox��0����'�z��/�ɰ�p��
��m�gz��y�ê��UU��'���=�s,Ի����},z��芙S�.�ʫG�UFǬ�sU���>�WY�_�$Z����o�q�>��>yZ������V�YN��đ�FNsM��?iԾei־qU�����
��ߣϻ�#��2�wS�g���i���94<�٦*�����{�����jy�:²��1�~���o�ۯ��x.��F��iž����9Wrʕ��rVuv�ӭ��De��S=�4�1?�a�7���D����lw�'AF��Ǟ<>�:Y2�C>��c�20k ������3O9�}���~�*��}f�� ��7�:A�oK�?g���b<�����G��}k��z�K�>�����2������yU�dV~>+��;����gz9͞�*T��'�5���^=�/�ا�b��믲e��t=FW��}2~�ˠG�|�o*��ҋw����AU?�=��<�����?k�"<GX�O�z�W��Ծq�g<�mfX�f)���eQi�an����o�f �Y�lr�իW��6c��ǡ]����z��J��q�SUJylX�T{v.��χ�Ku�2j�PuY����,z�`�I�C���'X�>/��:��u��}���m���]y��� |:sӫ0�;�2��	�*؎���1�������c��j�C����8��sgվsdߤ�T��C��k�ɰp���J;��D�)���|��߭�J�j�+�F/Ϫy�=�k���v��`�E#?ǽ�?K��OUP�;���F���W9�K�i�q����������e^��EH����0�����?n�c�hw3��l^�Qu5�9���O5E�ޓ�UӚ��e������w��ْ�zƳ$��V����}�
&�Z���Z����9���=z*�F7��;LO�^����{�����567]9��fEG�S���#97�m�뵝���X�Ơ�����sMg��V����sO����^�{o�5f�kܿ^��^�U�����ٳ��nv�����QUMZyδw0zz��.��f�a`��z�o�,kϟ���V�M�M|�ᇛ��"O�^<�{K`V$��
�D4*˦'+�|�TM�w���̒q͙;a37�)C����7��%����}��w���g23��$3)2)�e��d�J$XJ�
0<�x`
ex���'�F2`�'�<!�U� I,ҥd�3�l���}�����}��/Ϗ���"���w����y�8�>���9�t�0J�Q�,3�=�}��.Z�E��b^�m�}�/�R�t��wu��$���&�8�<&PG$2�+�Ҵ4bY���+-V:��w�v#�:�U����F6a��B`IԶ��:-R ����tYv��z,X�z��k�aO�yϲ?qj�_&���P�#ɺf�9�]ϖ�R&f~(,�'��8��Q&$��)-Vd#�.4�&��oݺ5۵/���wem@4>�!�];��	L��{���c"5���
&�eI���YfU2�ipﳞ���i�k�(�*T�����:G�2�,��/�f}�7k-�K�n�Sԥ�U� yT��,�-Q�ciLHU�b�&��e]0���y��rN2�b���$ Y�Z��eJe��
,u@)��N�!�X&&,I�y�֢k��e��"�0�i�Fj��Z��@c�s��I��:q0�_��ݻ7����0[H
Q&��D�)q��3f�^��J�uͫ�5���l��>I�*M�����S�˽ui���k;�%��$bh )sB����U� ��?��)u㠋r]Շ�	3k������0��4l�S�^ί��3�g�C,���@��s���ss��d��C���'�.X��6���ԩ-��u�0�|ca��Ĝ��?f~�ۮ���dzS��m�JSvZF�yY���g�Y�� �����;�a���w��@e��u�	3"T!�,~)�,�y��a	ck��>�t��{\����۶~,IL��5����J�,��R�aV�[��[��Х^��WU���x�s�'¬	uuXU�ޜN���"���$SX��bE��ry5�f�e*���"T��QK��״,a����KV�B��	VKXA����h~<	�N#2�@ש�~����Ɔ7G�Ȁ��u{�ch�$-k�N�s���n��,[�f�	;�P	3y�=O�d�LЕSa!f= ޱQ�a�M)�:P��TX{֔������h*ˢ�0���!�}*+��E�"y�%{Ј�>�N��R�ߵ݊�����4�����ƒPB���b�;$R�٧�d��V�cox��u>/¬mZC��,0�ަ�R��l�Ҳ���������S,a@����c����ݣLL�FmD���Y_��Y&f4˖c��Z1m�������>�d��rnD˭GY���֧$���7�|�	3"ʝ16��,u�xSbP����u��EێU&�q����W��y��/n�rZ��O��ͼgi��S�1�U�u!�ɯ�y鶩4R�)M�L�=u�6.v�oү�A�+��]��1;�>�\��4c<��,=ȑr3#I�	V~L�,����"���ϛdZ��b�+�D;�N��>U�1�0��~Ŭsб��0�6�#�&�PxtZ��:a�=�:��Y�<����ou^G����(Xk��	,��,���Gg]�Kk$my�]�仒gC f`ڈ���N#߅%-/�Ux"ްC���z�<�LAQS6J2=.��G_B���w�Ӧ�"	I�t%h��ӵ��,rKcü|�2�r�VwMռ�wY��g1��{��V��(�9����溮�w�G��h?�w]�ض.�wwuh�
�����㘱�����b\D�X�
&)��˲L8�5�%�-a�|�Gz��Ŝg���G��"�k���.�yo��"�N.C�Q����������K ܊8G*a�������Cd�lL�8���ʞC2�����+�X��ha�u1Q���{�|�!s�̻��uT�5,I���꺮�k�ƣQ6tyD�.����\L�L���a�W_	M:�e>3?+�Y��.���8��錴��1���~�����k&�9�w&�¬Ok�<�S}�EC8�������Q��H{�Cc�Չ�:�e��%|$$Y�W��B����L�!2a� ���[v�(##������ed�q�q��݈�a�E�A���"����2,##G7r=�!��U��M�3y���Z�)f�驖����7����h�2���@�lX�p�����Lx�E��b�X��;<g�g�)��[)�j��8��}�eb���yds\e�Dn�6,�T��ԁn�o�^��p/�0[fX.
22��1��3)!�m)QX�i�ΡY��E_c�o��k��(�XzD�@����rt��1�A�,w�vߋ�<�->۔%##��Ȳ<�ӭ��ݖ����,�F��̰.;{KF%�dKF%͔D�w��[2&�i�M�F��-*΂2��px4`�E<f�<�+c,C�����,]��Pk,{���|ɢL$��O��#R=���=���5�"���Y��:J=��߬�ZLM�W�i��"�Yu�vH��2@x�+���L	��,�'D��e-C3a� ْ�θ���Q�*Eګr��d���$V���CT���NndtC	������PGF��
���©����=��#�j�y�C���G�m��2��(�&d��z��B�5&��f��Y�=�32ځ��Ά��>��,x�jh�,���m�oRؒ�,)=m��H�eG�t�&�~Ц���j���Ʒd�Ⱦ�tXf�Z�)��rǺ�e?@	,�<��H}�떌��>G�	�f����KQ��{FFu�*����ЇA��6F�%yPd�g�\�i#^�eҌ�\w��~���1�ɲe_�ux�
:GH.��hB�v	,RҬ*�Ev�[�0[ ��\�F��]]]ˈ�U����{�����y>=o��Q����Wײ�s��3.�E]XԹ'����������|��*�,�
Uy�Q�.i.�6�E�_3:���n���2�L��>$Y�w��,
�k�y@��eF E_(��m���*7R�#�ؑ�ˎ��N�/�:�l�,f`oo�~�F3�'�׽ݭ;��p�y�X$m�p�>�+��v̔�6��׹U��X!��,�>Ye�Z�]Ǚ�:����H_c!�c�?k��y�V=g��S�f��c�{�j�뼇�'	�"�>b9���4�X�������|kx3`x��m�����YA�4���E�q�B�m����R�׺,rC�ZOL�\�t�p�b\�D����U��A�<�X�@ֳ¥L&�a&�-���q�$m="f࣏>���>/ktYFFFFFFFFFFFFFFFFFFFFFFF1!�(rB�=z�(ܽ{���_�oU�3K�}��������Ž���q�L?�U]/�/��x<ޕ�?��7������~뭷$�,lll�����������GOɌ�����������eD��D�Mg�	d~pp�}�����~��L&����x<ޑ����֧�����N���5�lll�}���޵|g�0��w��o���?�V������*^�����FS�777g�d�n�
?����Ç��������욌�����������E`��\FFFFFFFFFFFƢ@	O%̄O��>�����G?�Q�q���w����i{{{���5r��5��g��s�΅k׮��{�ϟ}�ٿ��?�����3�)�lZ�/���?�Ͽ�������?k�x+�yę6�����;w�َQ~M~�H���������������������������G��+&��oµȻ-	s����@&��'��^�V�CM~�p�B�z��o^�r�7�i���?���-ߙ"̦����>�菤���dE�PEy�L%��$�T�D�ic2�����������$�'o�������������A^_-?b��������w�^4�Ln�]߅�嵳�3#�~����_����_��_�)ۙ"��ݻ������d2���Ƨa��=&�bMR�2݆Q���������������������������xUg�iВ:�j��|F�Y��'�G�&��$��l�V���<9m�֭[�1M��#�;S�����󇇇����q�#��z��2�&�$��I������������E��0�����������H�:�*8)>6K��b»�������o�uJ�	?�g�)�#�m<x�K!f�Ŵ����6R*K*7�S��r�T�6�6��.�!/�JSv��&{Q�m� �����:X$V�Ym��W}�����r_�=��ɏ9fX�g=����g]O�u񁪩`�9�y�[�9�-oq����K�N�ca��2=�{~��^��)��52222bx����u��C<��m�cZ,��˪��a�.��-c�`��˴m��(Q����=�!�2Z�3E�M+kMXH�BQ*R*��8Ug�	Q&��\��F�)��ě��o������4�4�@nPC{SDۼN�6?���I$4A�.e �+��V�3����(�x 4A�Te��w��?f�B�	�sH~քZ����	����-�uV?G�1�_y���װ�R��
Ly� I�w�m����'+?���D��eB���Qݍ%�2	��]1������.h^ވ����#`��ǃ弇�s�D�3�r�9TZM�}�	�.?� ]?�ꓹ�-����mZL=�%�R���ꀬ6�S�0aI\0�Bt7��,k�\Ƕ	[�~�����k�ʍ�|�缍k�?�|���ȱ��2}�^1nc�Y�<2%�Tw�m�w�Wӈ�$�
:�Lp��2�Jl�=�b
ꔛ�@�|"��xB�a	=�u `t�1g !��	�*b�|:���Q�5Y:J�7��vK���!��Y@��M}
-3Sv"�^�#@��lƂF�}��Xeb.�@뀹�@�\�"ix���"����4~[��x�R�̷{�`�R�ܐak�д��J�9_AnX��"uT�����w(�g9� ��c�i3�&x�8�3�c�e,�7��
q]�9%x$̘�vv� $!Δ<�h�6N2Jvj������Lfe�����c��@<x�q����ƝQ��:f:Lf�rd�����.u^�!�-��POP$���eB�48 �h�eb�hߴ&��}��3?�y�Iɂ��M��4�ѲH^,�`&a�rPBێi�Ȱ�(Q=	"�G<M��<di�Da�G `�ޜs��"��<�ؠ�*
���.N�ְ��פ����#�am�ѱ�����tok�0;�F�W����-�R�w�N�v9S�JP�a#c�$�F�>id}�a�,0�Ցt�^� kз�o�eؒQ`Q��$,$��#af��c���w�ȢT��м�y\Y�l�d��Ӊ%���IR�%A�t��,�=K��:'�8moƵQ�:
k���BZ�K��3-��Ȣ6y�9~ǟ�tQ�9���b��gZֻ�xs^`�h~<�Ӭ�ӡA<�T�em��]c(�L���D�a��K�V]p�Uƙ"�u!���j!*�!�.L�z��x�6*Y}��%�'7k��:���@�C�d���'&� J/l4-��s^��ń5q��1����V(�3�,�Gָ�✳hZ�(4�f�{�ތ<�cc-Y��m����<U��r:��4���2҅7������;V~uz7HS���,0IJ��N	�2I��c��U�NW�9�LPE�5E�U�ߔF|8�NȬ�G��0�K��ױ�a*M�;L2Z�L�_/����\�Y{�z�Z��u�E�e�H����F�����Se�
̼�g��c�Za;�X�z;0�����w��+T�0I<�1��쨓�(a=�#����xʞ�X�g��b9?�Q��:{(��צ�R'�$^��T�q���!�9y��,�����֎���㟮�T�R�K���f���ee�k9S�ٴ�ƥ�O	��Ȳ�=u߫�N���,#:J0=�Y`��3�x�(�˅X�[�t�h�[*�1>�z� `+��ud�$�ncf�|�� �i�5�z<y�h��P�ng�g]Ϊk�R�LOI�k�U&,���x�25a��G��	M�'sZ&�x$�Gr��[���1�z��UM�+f?`�,��H~M�Ѽ<�U˶��g����ie���s�5��ڱ����>f�u�ڇ˄��e�-c�c�b�M_]m?g�0�BL�ſ�I4}�Mں���SFT\~��ۃʅD$ J��	�54]���My!gIYo��
��:`o�e��j��FѦ�b��M@�ZO�k�\Vi�Q�`=�[%�7>�(ʒehy�z���Ѕ�+D!$,ˀ��)k#:�Y;�,Z��Y��s�'�F,�.1�<@��h!ӡī!k�f��:kB���l��j4��ڱ(N�*�e�ur�#	�L��.��`:��Y�����[|#c�A�\�{q�R]9���C���q�b��]�s@��������b<��<�����*�ʤ����ӱ��L/Ao������p���ڸ���D��7+-�r�����W�Q�a���ܚ���L┑���3�+�42�V��6��m�c�]��;�P0�j `E�1�i���q��4�(�`듬�X`�=f̴��'-ת�u��V�����t�iX�[�����;s����Y0m,X��5����#:�X k�SkT9��е��]�c�0R&���n|qݷ�o��qh�]dԙ!���������?��o��v���fB�����Ć���V�0���d�Y�"L�w�]������������g�nnn6��z���&�h G�qA��z���x�N",CPʰ$J�=��*�����^�)�a����VL����SG�4:X�����s�"yuq�aa=�c�x�9��6X#`�cf{4�A�X��}<��� MǛ�`�o�g�#���Q$&k��6��I���Og�>���r׶j[��s2�[4-�#�e����[��X�9_�y�.��'�Y�<PNFw6R�B#'cBǻ��'��tw��6�ք�_��_��|�[;;;/L3?)��L����N˸v�Ν����[����(��g?<��ŋ3�L*S��԰��s�L��w�ZQ�1��O%ʎ�g�_?Kóu��H��f%�2����q�><f,I��.K�'e�?o�W`M,zEa�#�lE����~3R��j	�y�6-���.o�!d�u�ڬ���ѐ�lM��\�x�������*�Ui�g!y+��)�����!��g�j_�I²�]�����
m�b�H,���<F��Ѻ��[�2��ի]_9%��cU��<'�cb.~=�m=��kQrLH�i�k���{��w�������������?��Y ����	+)�s�Nx���i����f�X�0�X�hc����oz���ŋs�C�Ҍ��>�?.{�`f�:@��QX������L������ @a�����3�2?�����2��a�̣����q,X��=O�r��z��,�8f�[eG�E���l\��ֆC�c#�@���*G����t�t(a��㊖�"㥪?1���iuEy\y�G;�G�1_ϻ�;�~n=�)�����'�����T�ɳj	�o����;��Οܼysk?���[�n��>�(ܾ}{���6e�|�~ֳ��]��Ç�[2Vf�Y�:��=7U����w�&���m�.��@`i4�C!��SSZ�O&XJ �d�\�\%�֑��1��Kw��cQ�Hd��b&�h�!��m<��lA�I$�9���Ӻ�=�,��kC^y}��t�����nM�vP�j\�V.f��!̚�.��^��&N��!�����/QR�g]�ZH~}c��h�o��"H%��2P>I�\�#��oauM��0���~�����������-9�K
�Đ<��K�����L//�3�T��j��0?y��0A��(Y�b��|�w�_S{Yv�ʕY��t�{p.
� ���yP+ih���r��2q�2�z4J,;,=��㳏E�<Xz��i��U��e ���t���a���夅��ז��3�x��SvH@ʎ8����~nIp�yˈ�!`�lߦqe-��kx���`�M�e|�E�����h[.� �,a�|MD�֖��(4�&B�Ox N�$W&�0t��]Ɓ�M�:l�����Ѩn_UV5������{Tf7o���[o���/~�Yd��?�m�����%�r�%�V�'��T|L��Ao�%�2�U^�,��W|,��oRrF��f�Ν��.eb����A�d}��%�*�U�}KF�>-��l�u�1��[_�F�}nXF���Mie�7JxE����^� �$�&W�B�i��;����!Xf��L�{Xd�G ��:���pKY浟��i���o��kI��#��6��|2oH��*�6u�*g���!;�9��zZ&�R��1���!�����|£htbj�5��J6��7������,JȞ�������_q᭽���2�¯��+?�[Y���M��S2LYQ=?M�z�F׭,�I�#��VS=x�|��D�(,oQ����&x,;��k�^�^a��؎��6nBa֥^<.2��8Wy$̺�/�M]�U�8�3�W�ݐ��E�c�����OC8�Y���^�Y�{QX�.L��)7�f]"����c�٬��u�p���T�o���-�*�>����N���ܘB]��Od,0m��k�/�#�k�ׁq�S�����f?�я^�������[o�2�q4��D��nO�,l�!e�+&~W�L���2}�u�j������2!�$BO#�؋�Q��6_MeG�������J����D�������e�	jm$@�6�"����h)�ܦ��ǖ��7R���'����ּOv����l��a�M��5V��c>���0U}Kp��<�I`M�	��\�^���t��$�t�ǌ%�hӦ<-�]�tbd�)��5�]*UҬK���Tu\$�Lw
�GbU��U�yU�fy�����������޽{�]�TC�43�ZP� ��dـW^c��_��V�91ɦ��IiH!ˈe�邂�P6��3��ׅ7�V���m?�6�2�`�9�M�b�Cތ�C�N�F�eY�?��j|��ىi4c�o�И�`��[zo�c�/��X������.�^�m�kS�H�ѝLghK�nY���t�k���>�D������Lǫ����{�-��zk]}���-C����b���"�x\-�&���,�)y&<����P�b�3�٭[��u�Νɳ��QE��Wej�\A��Ƹ��[��[9-~�4��i�f�p`��?���|��%K�E�.,�zrC`]&+��XF2���HѨ=��g�.� Uܛʕ�q\��8�3L�����N0r�+Va�������X�m��,���&�eF�����n-���>f���v���:�Ezz�"�����(S�#2�͜fYv�:�Ƽ<��×l]�c#h2��q����y<���q���}�Q���!v�a��^��5�T�i/��V�v����� ��fq�4͘���(?�Ge�����������͛�|���쳲�U�����Pe�ɾy3� q'�ɱ��y/i`m(y��^	����X�]�	�D�P�q�F�B�"�����Ǆ����X_f0=����5-�P̌,b�h^H~){�7�?�}��#�5�=C��-�`A�c�7d,�.ӑ�RF�8sKX��5ȳ�q�:���~�`��hZ���:`�{���t@�ǴY��h]�A��������&[G��ɻO�J�&�\�0��-a-[X�<ZO}:�e�"6�>�Xm���n��#�o�;ƤZU��֍z_���*3�"�~�\��O~���1����xJT) �o];�@B�mnn�^���'li�F,�L1$�6�F���E̠ªO"�+�-B�@�H�����B��x$����j��v������,k�'�v��d�W��\t���6��`�W,uSt\1�T��-��u���>�Ǚu�Ju�B�b���1����<��R|>v�e�Q�u�6e�7/��HYֵ~=ʨ��-��~X�+���*����lQ��\+|���h+�E)�"�d;�>��U9�L	�T'$:�fC��Y#��)�)��j8�����X����ˉ52{5f���f�cnmTE��������L���j@F�Ƣi(X�_��p�@���1ǋ��y��:��б�3M`>�G/l�zB�qBӅc����KWD��x4 {$��u^e����}jY�'aV���`z�[� �n��n4��-;��X�H^L�\�uLgK�a_ӊ#M�4��(�fZ���d�����\��`����tgr���cUi3�d�����:����Ç�pQ�.�睳�]�x��y����R���]�D�u�[@�gL�Ցgʆ
D�H߻w�)�9ġ��h�.DWx�ayâ
?CX�F֘����$n},��r"��fL���ѴX}�Z�"y��@h�����e���#y��іhZ�:M!`�M�V��0����2<1�e�gQe8%,[�s?rF$�  `�N֙�(��0Cʄ���|ѳ�X�_&��TE꼋�QeƲ���AҌ��5�>��
K¬L�V��m<�u����p){{{agggƥ����iʯ�^��lz�0�v{�tIy��ĵ���RF�~���ϫ�/eHe�MaFu�͍���֌�ϟ73��`��	��A=P����21,0'�>�)�Lck�Y�M���0#̘J���-˚��)�;˅&sa� %�=0c�h~��,'t.Fέ�vzc��:X�E���2���p�ꌦ�>f��c<�{C��:x,��)�3���5�ɂ0��>m����dfb�q�ڦ��X�Mɧ+��Z.�r��WtKFMSv���ޞ�'�7�TZ���8k���iA��0�BvM�o�c��W][�����MT�1aI�A����[[[���ŋ�u�%M@ˌx�!9]8xVL���N�
j�[.T���Ӛ0��G�~C����&̬��`y%2a�x���c����I=58X�E,�Ժ}s�⒔]����:���N�K��%�c�����	C�)�YnĖT����\�|>V~L;�L����������<�Ȅ��S�c�3�2n�E�I,�+B�1�c�� s�lnn��5M��«�K���?������'�I�u�z45�Lv	�*��~�mS}���F�	i&o	�����"�Xb
KYI����#�l^��-�XF�然�\ �iL�h�e�k�#�z�S�Y�+���h`�Wt���c��+�1f�Е�8am��P}fC�X��=޲�QBM+U�ʎ��Ʉ�s�X�i�A{�tP�d�0��-�e4[��Rw���QB���q�%X�E�	֊�R�7b��s���$u�.a���s]��ԭG	��cs]�}^�ڠ��J]�2	%K�ٞ�HX�C���d�'j��<��뢀9�"e��$��,�,��H_A	3�b��V4�<t�r��B:E�*��:
�~�$a��Q�$���28U�[�g��8�D�����}y���a���]ai�`��Y�yS�[�,�kl�k�e^�NĶ`����Y;2m������ү=�ͪ�c�u>3-�u���d����[��wmqJ����?�x���o����
�gqN'�.�[��D����� ���&�5�E��lh��*���PX
V~�񂹭ˠ�Dm<*X<
�#(ˎ*Y�zA"y��	��CP�A�!��:�>��Q/k�K�l|c �9��窱�1�k^g�%�H�Y/"��Be0���h5�v&m���<�-r��̭�4�&�`��hxj�x��W_�\3���ܩi1�c�V���с����!����?�]3t����m�隗��F�չ���l��΢J�b�ZWF���)1ԦZ�+��1GSW�E��Ԣ������o��Mْ����aq��N���g7��*�(�I������)C��ו�-'\KC;�
K�g�����XJ�^g�ߢ�lQ�����Px�~C�U׵�?k����7%����e���hkx���  ���i�ѱ���@k���S\&2�b��Zw�����<�N(<�`���:���qj�f�4j�Otq<`����0�"V��8�1�<�s��@�R��T[y7�:뵜ufAy�*�w�R�o�{L��uUǇi���;'ʵ�ϓ�q���0�&�V��{ޚq�"��fpœW�������L���u�}���32��x����h�0�� P7���S�Ӗ��C��s�����"򮯲z���G��+&��]���fGGG[q4�
2�`jo`YZ1�����Ba陚�G���\g mڸ��wQ�=zj{DQ���g��:B�}�X��0ψ��ѥ�r�y^O��24y6��^���2�Y�l�>�Qu�[cb��r���@����g	�u��oىa��*�f^�#�R�r/�OŻ�ż��������!q��2��@�ej;� �"�2�E6fd,�H����QVy�A��"�e����npA��E�Ǻ��*I��m��&ɺ��=�(#-XE(,�����.Cj��r��"! ��cR��=�g�<M6�"����Y&&��c�b.&&�X�zJ�M&������=�.�(,�A�z��6��,���B�(���]�b���׍Y�e���T�b��)����"Ke�����EW�iy�b�����H�Y#�~Z, Fܶ^H$��C�s����iե�U��(R%�Px$-��wh$�5�by�4�G�[-��U��XT<%̎�����	%���:R�a]�ϩnW��,������RSG�NԌf��	k�����>��T�g���X�6�T�@^�C�bTG)���Hc�^$��q�GT铩<g*}���7<E��X�ey�i�R˯ë��m|1�61��c�lG�)a��Nq��-��H:(P�K|h\Ù*X�1r��d�(�s�h���H3V^˾x��W˽��D����j�*�m�<-��q���,X���+눏�j0��Ǩ�����H��7o�.�#Ӣpou0�x���z�-s�X�2�k�y��oY�L��:(�e���#���1�N	�ifk�p|�Z\�:x5.�!cf3�?3#md�)#c�P&�2҇GY=�O��T�9t�a��وn�<����Ө��u�v��Q�Л�~����[�-B,v���=]�U���n
��HX��J2���"�<��ʽ�ޥ��{]�Y|�b����k�R�a�*+�V�u őe�+w挌�����eE��.��>���s���`�Ȳl0x3R5��}%c ,��%�<�]���Rv&��7���-�T�q\��r�} ձP>�,�⣸�x�S�����/����x<e�~�ϟ�}�ж��hsP,rZ��9���(�����3�fܠRwz�6nS=Xo󈶝�<.�� ��!j��<$-)SS��̺r�[���
9��h�<�OO�����ݾ}��j�Dǹ��1�2!��%�e�n�����k�2�c���y���q���;mڍ�^wa���E�y�c�1hyX��~��i�2mf=�j�c�ǲ%��	�ݔ<��P�~zM�r�@�D��C�jB_򵮌���ʺ��u�;��b]�:�sP=b�y9?f�c�XE�2���i��C���9)�"�T��������6�{�uNP�����$��a	C�6#��z뭭��ËZ���.���rY�W�^�:)3����--�q�7�[y���.����gfL�i]=��S�`��G�.'$��Λ�,���Xf·R��h_a��xlߢHW�2	O���7�j�t����d�5�[,�<��:���IC�tR��G 頄҇�ye"BZ��\��T����mN��6��e>���.2c�6��#1�L�,�'RJ�.%�W���)=t׿6�<#�&�����ÿ��N|6�@�Ц���V�W�[YX�c�A��ߥL�7P=�����N]�`� �XN�<��a���X��}�i�bz�e4�M=1HX� ���ч	�N'^a�bmL�攰�}��9���������~7�׷<�C�ǔ�,��i�gى��5�i@F�)<�����竻�e�E�^a�Q���M0	3&,�-�vA��>��R�a�y
4�W_ʿ��a[�3�.��'���	��+�1��~�#����L��ϸ�č(��}���ig���͚pۤci�d*KU{�V	rF��}Ų�Y{�!�H�tXc����b�����袎���q!�"���=�Oz�w��O�:`Yb����>ˮ�xtd*�X7�w�1�B��M&���Ŵ�X�8k^Ky`팈��-��:���ٲj�Ze;d9�X�r0����x(�}6&��d����$�H2�H�(a&���4M%�,��)�L��0����`��@qVEl�#�t�E����9�<�Lf/�4�����çB����D:<z�#z5�!`z����	lO�&x$�#2�E�s(����Hǔ�|�3�Vaf^�]�$��#`Ei��G��y�S^uf��G�5��m�Y�Z�+�6�x��`YvKא����v�yi���X<F2�C�l��%m�d�wB`!e*G�T��ˉ�(�r>Z�e����u��\��J|�i�#�bF��:0;88�(��`���AjZ��%!�ʤz_|�4e@����=�N�oll��R�5!�䷦��:oF T���6�+�R����v<�fֆ�21]�z�!������ϟ��!�i�A�A��p��XG�ٺ1p��2,�h���-��lc @*�M@uN�1����ѠbMN�Fg[�SX	C�sV�d��TI�!`�v(Xg����z0B�0Ǟ���z}�v~D�d�O�}�2��uyu9r��L(y���=:���,���L]IQ&б�(����[����*��<��7y�5q�V�3�ْQ
���7(s�d+�M�|����ʠ�6��+�3�J�loo�s�΅����~�:^__o,7��xSR�	!Ր���S�Yik��CU�"��RΆ�Fc����`��,y� ��(�<��S�9���ΖH����aH:�L�q:kXGw��T�Yi7��2?L��#a&`y}[c���XG��rz%�+`�u�0B�		�~�Ǚ0�`-��sB�X�y�u�L!S9Մ���)ڬ)Ϧ� A]���Зl��w�'<�vZL�L�S[�n�((�W���8+�g}ȼYI��(TBH�l%�F3f�}�Ύf���F�3}i�Y9"O�1!�._�<�gww7��Ջ�EXfͯ)O!A��NӤ7�k<m��R���.�OL�l�F`��D�Rr����o�:���H�73J�Yz)[�9��Yn� �Q��	��&�6H�3�tJ-�L������hX�OV�3��h$>���$���Pʃ�Q�&9Lb���M���f�Z�K4W�o�qŊ0C#���AU~H:}��]P&)���㺉hmGaډ�'Q�L c_^ڷ5�L�5����W��J6-�X����˂e�Y4�6y��.�2T]�
�֑�S�r�K���>>�N�%�,�����h��
��UP�$��64�Ff����,�ka��c�[vo�T	3��!��
�Ǳ���}k�e7 #H�٘NZ�V��'AW�sx3�hZ,X:1�j�b֘���5af]������,s�{����ݘ�w!�Ǫ���ǖ2�����̎ʃ6;�0섩����G��u!E=�1h:��)��R�L_�s��f��T�H��X}�a�-�H��+��Cy\H6AI�rš�U��ĘԑD���o�W�lB��yoo"̺��O0�f��o�X��RA�ZM`�k�����O����by��H@z������q�f���[���-�D!�t@k�i���byǣi0�#����F3�]���!�s�<�=�Qt��}{�[3�Fm�u��a-�X�GC�[HٙQ.H����8�h��#�zJ�"�1��&�Y����G�T��f�vra�i\�!TsҾ��j[7L��Z����Ӆ4p+�-ޕ&�6U.&�y��^�h��,�{stt�%�	C�YS^f�~��B�q�^�5�8~���h��քs�e\��Ǆ���2ih	D>x$��b�Qk#:z��%�u0:C�[FNe�(Ѷ��Ne�W�S����:G�,��F_o}�z�Af��L��ix�^�1ѶO�5���X�3e�3�o^�X��E2��K)��c�O-�V��5�:R�m=�2ߒ0c�e�����:��&�u�.�ro�߬��>�k�������Vq9q�Y�N]��u��O�;��]�5� f���֖m�J��՗~׿U5���e<��E�P��h*C��v'C,Yy��{�/M�o��-�,���ǭ��?o���+`z�<�<�9_y�fs;��c�kR�(��2��d;{Kق�|$?T/c �?�vA�PB� `�<�QR՗�� Pg %�@�&S�f���F�EO��r�5q���1ţ</���XE�u���I���Y�&ެ��u���CE�4d�X�0����m!˫�NU]h�S��:neQ�68%�b�����d�8¬�ڔ9f1��,�OܘUm�e)z�����e��eԉ���g���T�eB�)U2>U��i���u_�T��`�DK�YO,#z��m0Ѿ����I��
��hzFİ/�-�X�����<��K�'d�u��-#��X@��Z�헪<G�$ ��$J<:\�Y�7w,���\�X�D�rW��g�1�$K�>ӎ�*��iU�K[!��������_-u}�����c����$s�c�	=.�K}V�[-U���R�:g�q�PWq`S|�߼ .��_�������Q�*��5ׅ0+���3��=3�8��R˂,����	kr�	h�hA�5b�1�#-S�xy����7����j�~P��i�D�*L�ZF�P0e��׷G��G+d�3�\�.0�s���=��C�!��
a�BHæ����E������h~ֆCokG&�m������z�U�3�f,��i��۔�F�@��w!�x�%Y	�NomI�E#$��ת�لs�#Xv�͋]�\Ò-���k����]W��;B1���.�nj�/��H �����N������^����e���,d�){gV�؛�żr��ڄ��7�4�6�\/�EH�?x����D��k��$xXFm��@�1#�6�y���s!�8�qѣ!ȣ�s�VX�Ś�M�y3��|���.T�>��Y�1	3�Sӑ�)-��B��Z C�.�b���,G�!�z�D�5X�L';�y6�u�e�jC�����n��?�����h~m˴(�!���2ͻ�a��M�Yf�6v�Em��fm�D�N<��"+-�.�Z��� ]4�I�!�b�kc3�7���q�Xm�:[6��
ݎQ�S�Dy{���Ț$��d�V�\�*��T=W[��`�Fy��:��	y���3cJ��
���TK��d*g=%Y�,ZO�Y̅�W+�k��`�k�b-�ǋ5�Ąe�Yc�����ְܖ�z�b�Yv���$�Xf(Y� Y�2�3�~��w�SkH&,�a&YmV�b�́��eY��k�E��ʃ�f}3������T����2a��lֺT�ݘ�Kݠ�$�%����vlL�0ksg2f�Y������|]�0C�����VvV���S}5>ުLB�e({>V<a?�P�E�,�V`��cHZM��|�!��RYR%̶��fd٥K����*7��ey�Xz*	<*��2���lB�	^�9C(�,�.�ta�5����97�0Z�y��R��(,�)�X����������r�C�B�4��� ��'뾂��΢���z��S���"Qv)f��^-�U߲�k�Y�;k�j��P0�9s�֕��z�"��O}��#4���cr��9�HZ�s��E'��M���1����]�1}�3��cj���e}חF�Udm�@�	,R~eR��m�׃4���꧜���V�2y!��ϗ��{a[{�!�hp��pa]�Y����{� C��蠓j?����5i��Yc�J:�9��d�Ek���f�ZN3*��,���}�Z�iz����a.�4��贉��Ly��h���"M=��u,X:?�`�fL�>&�Y�#h3�1�s�\�r>b��֤}�1:o�G#̬��>�^�w�Y��(���ӡ,1���]!�o�G�R<Q��MJk�L�U�,�K�<���o�}�{}��+)N"L0-K1A�
uo�b�ɣ!���9�%:�	�^�����C�Q0��ȡ\D�"�=<(�q��s���L0��iȳ�+��Xc�����A0�N�Ƅ&0�-0�Ik"����PYǔ�ֺ"���1� ��&X;|���o�jߙW�6e�^�H}[�{��)���� �+eCt]�}�O�+��F�X��Z�0�,bq�H�y�B�yt�X4�8�Iv��$�PPގ1�[�XӶ�#��������dT�L�J����4yy��e���P.':�j��pBIO�1��˄$�&u&e������pv�ܧ��yT����� `*9LX�!����Z�0�fֲ�cTqa����wL��#e�6NyE����\$��[�n�w)-�� s� mlM2ѧ������e�{\[FY`����q\�N�6e��E�%�dE�Z�t�&��O�F���Z�N�h�%d����x+���9��ߐP��\�bʯ�D��)1�]:�+����@9��u�P�<"��r��j���>����a�(��vRm���.����3222R�-����������|Fk��W������k�ǰ4��K����=�eC�h�e��=��kZU@�.u�7�祯9�
��ǲ�E�!�4�#�,pJ�)����>��1�eRV�
ufMaz��Cޫʐp{x���h��U��>�e_�g���gF��}�'��f0�WO��d���}����U6��i01�|��c��W'���������w��k2�%�۠�:@�uPG��IV��|U����I�{��`��Djyl�rE�+�+Yn��G�e,r�M�⬍w�7X�م�~P侙AF����qM��1{6��2�CDnX�eE��*eCeQ,��w=�Y�}�.ք�5��̯)�:{g_Q�UF�4�ց�`�e��+�[z��zS,��'��������k���x�'��Ňg���H�Swx�J.�o�G9O}?�^rC,�,�(&ˎ�Џ�a�6�\����(��q�e����i �q��X�y�8�z�Y@��Ƅ.�þ�c�Y�.]�Cg��3���!@�Ð�Bޡ�M�ov�XvZ���4y/R^�uZ[ԍ���+�9���htvl����ݫ�$��hV��0[__�����֞"��\2��T���4��ۤS��.���٫a�u��6.r����YO�8H��y�B�����/E�c�����L��lِ�3?���蜾mO}:��u�)�yH���{�ء�����|����uˬo	R/?
��6o������fkkk{�����I��~���b����B�U����(M�Y��}�c�e� 㬡Θ�qk���-�<�&���/����`E��mJ}�S"ˆ�5��1/���3�E�x�I<�\^ǋuF���87nQ"�}ܦ��"�����6��U��Aԍ�6�L��K8�2����!�f�0�s̄�	3tBF�����5B�	"�N�F��Lfg��>Zr#���
E����v��ǃOd'�t����L�,+�喛)t-�i}:�!��e�ǵ��s'����L���--۸���y�T�0k]�X�9;ti�2Q&/|2ےquuu"�eQGM!�cZ�y�^�5��ic��UfH�E�^x}ã7SF�Y��{UTY_�?eE(�Č�s�m��������}��I}D�Y!��d�V,�؛Gl��XW�e�<ʰޖҺL��M_���m�ޢ�jm�>�Fݸeh�"�S �ROm"C��DɲB^�a%�����*�^E�{�9Ϋx��1#̮]����ׯ������D�3�8���	����dXՃ��&d���������$rN�����gy>4�r�����ьH����(٨Qz��\/��{S�G	+��	���'�{�HT`3�LEIt����������M�ގ��<G��E�c�Z�,��r#�`4J� h�����6�E�k�MkdH~h�CJH~��,X�+��a٧��L �d�kޔ�d��C�ȃE�U�t��F�Cv�a��r���-�|�u��9���j{���!�ݼ>�ֶՔ��o��T�_��=n�k=��6Nd���8�`=�P;��]_�u��g��#i��)��t�@�'kNC���UGdi9Ն+/B��_3���(L��0*f��xm5��J(Nӗ������bF������0��8������f��+��2��{ZИы	��A�����m��g�C��װ�&�h����h�
ko�e�d2�����
��M@��T�K&�2�`�K z�({Xr1U�2#�~�lX�L�	�#<��ظ�bGA�y��~e]O�țy�Y�al��y��U�wV=��TG� �<��P}�I��1��}E�y��/��,	3�ў	�,�&��]�X3�>��m��IK�L��M� i�\�2	X�R��w	�iJG�Y� �g�x���M`�1V����>������>�X���<�_Қ^_��"�{5���3���ic���\J,����ͧXa��X�ҁ�[Ut�I�y�1����2�H�r=�e:��e����2hi���5a汞���X/4�~��ѫE{�����k(!�L�.�!".XZ��2�{ե�E���|g�W���U�	�YTU���I�`����n��L�&J��+�>䏥�=�yF��7�9�q
���I�!@�S��������|�̷tB�E)����y% Y`}}���4�L�V����Q.��m�8ծf$ٌӐ�B"Ɏ�o�7�r���(��퓝f��xW
�[��R8Q��s�����Trd�Īkc2K�D��:Rr���*�Uʌt�&�,��	�̏	�Ʈ�]�!ȄYg��Q}�I�#�h��87��b�u���~��D�GX�L���E�x�g��Cm�hjY�&�:0	3&��.o�7C�|�(�&�A�x!���k��He���
V���㔥�c�2��b�UY�jܲh:�uL��"2��ˌ��ք���0%�X+�pP���ĉ�d���l�E}E�ٌ,�U{L���V�at�s+�fGJ��mŬ�<��[�T�Tr��B��$�<賩�,h9zL��r$��.�V���A{}��F�L����s�����L��l� U��t��fC�c�a)�R�wLoQE���C��u��k��B,ƿY�aVu]U~m����q�Ɥ�3�W�#����0Nu\8��V�"̆(G_`�j���N̵�G"ӺL,0m�,��hc�l�u�E�G����k�4�g�<��=�<!�FOȲ'��&$faV|ʌ�=��Ҟ\ׁ4{jKFyW�W�=)����SZ��C4NSǑ�K4W9�|�$ґ�1t�m�(�Xq��1JR�J�YGXY�����n��m�s�̑SeuF��!`.���<�҅u_A�Uw�4 �
����ms
�蕔Qe�*�����"�Z� �U�V��:�v~D�`hǍ>���l�������̚�g�7(�e�*
���w�m��$�X��l����ɏ���G�#��ye���yT��������	Q&i�(Y���H8���o�Ϟ�+���1�d#%��=�)a6-�Dޥ��%�Y򾻻{��hCGU-
�Gi�[K#��%��E�N-{)a����1Y��H�� �ݹs' z�t�*ְnk�r`f>����2���� �=ԗ��`}hz	3�LֆC4r�QW�64�%��Q�fP�̺﹞>��r������4�!�7�1��,����v��HI�0k[0�(ҳ�	��ֺ	Y눽�l���QB�Eޠ�]����~o�7�L���9�O9��hZ�;ĺ��Y�9fޫ��.{=ͅ��'���Qf�'����5����giA�#�KPɥ:�L�� l�َ���9�eՆh�M�>��/�ń�.n4}����677gg�I=j�������̽ǅ-���f ��2a�Ǩ5R.�7�j@F}�r�ч���Ӆ�h.�LL�D�6�l�ǕW�1�y��Q��P�j��>a���/�"�1t!N�Z&�uP��LGgfZP�b����[oy�aV׏��F��c�.r_״�ub�G�C��5}�`�7�Ȳ&�O�,Cm���<�~��;�Α9�e��u}�i��P�P�SNE��O��4��x�����/6��ьT�j�����bպ<�ST�V�F��d����V�P��#�s(�����7�^���0��%�?>loo��/��3�d�`MZ�	�-!�(F	%��a֦}��a��=��(Ѷ��+,oJ��^�?��V휺�<���mX`ꀣ%ש��G��R}��"�>	3�zq�E˴(��\��3�X�e�}��1�+q��m�-2�4�`t�`f���6��6�H:�XG#�X�u�Zn�LJ$�& ��)�����8Z�,,�9p2�4����M���L¬N�ƿ+O�[�nqZ�1C�$�lo��`�㈲�f�Oo/����)av����Ν���ÇPl[ /$ "ר���+�S�f���J=�@�<666N#��]���%_�~4Z^c��M`y8x���P���x������ަ��h �b�\���ץ�zl?&���^X�oM�6���F{{>���~`-X���"�# PE��ӱ�������"<PCP]���c��6X�/{t�c�������um�>�o^Y��ꌖ\��b����u�$x��W&q��<0w,`��y���U��y�e��r���\/�ż�=��'e�B�M�4����Q8)��}�w���jNfg�Ͷj\��4��8��L�����s�VW�3�N	�g�y��˗/��ݒ�LY ��bftb��Ӵ^?�m��*i&!������r=���C��MH�T����XE{��x�̱>��<�A�F��(�X˅�u~hߴ�����X���N�Lg��G���L㛷��Ѯ]Xr�a�̏���e3�s�G��ŸEU�c�<,��ǹ�Xr�ƃL�B�1bې�H�N�����:{#�zNf�6�"Ṙ972ׅM�=��r����;�kkk��H�y����䲰�$bl�^kv<�"}vǘ�H'r~��,�l%����>)�c>gV_01sJ�]�x�k׮}�ҥK�r���S��ڟ-zp!z�v��H,oͨ�Ƥ�F��=<��nb��
Aֶ�hs1��ړУ�u�&ht��lA`饳��S)/�Rk�r������荏�啈�?C��T�7��ҁ���$7R�+ְ��(B���<��ze��ѱJ`m̴�G�ay�3��6�ԑfma�ox��g�c���^�R͇��k9�r�wo@ʆڻ���ղf��\ls�>XE���kW
�E:�5=)���O����<&�VW��K�(�i�M�AűD��fdYQL/,>݋q���u:f�a{\��0��W�z�ڵk?�p�¯HBB�Hx��6�PPT�hJ��0ӲJc�bUI1M��)S�(7��,��y���	���4�\�R�\�{5T65�!2�I`5]��5�bE�>�9͚8e�<�7�r��ȃ�#x�CQB�)ϭ�Tv�ve]jt��G���e���MZ,#Ko�hc�,<�5)��@Ί4d:��v�\�J�/��;�(���P0��4��A�LC0��D���R��7չ��Ms����*;X�i)�|�7�Ȳr9�zB���g#�]�c����g�IrN�����keV%m�2�|2+����Ō0���0��cV6ұW<9�lF��k�q�e{{�#9PV�²:k�����F�XjȉP�Wo�(��ԧ���lL�,��udQ��¬	H�h,�E� �9�IG�n}-�xf0FY}
����Uu�����t٣�<������Y�8�c/U��c֑"���m���ȼ�̳�3��\<�D��H
��1��-IK_�v�az�K�K1�I�m��`�x]�5m�}�:z��6ml5o����>Ye�������g��ʋ�x̴� @�`��|Ѵ�X�E6�4C�j��U�Ҿ�<�>�����IO��������z��VFѽaT6�.=	G+��F��u���������x�'Z�ϟ?O�2��f
��,+w�x�X��F1�wS_b��^��%��̬�p677�aJ��H:,C�<��	U�P�5M�Jm�M@=��F����D-�O���j�P�r��X��fC YhZ.�FNǔ�H;��ZW�Qz:�Y �����֗���|�<��o�񨡋�z�~�Y�a�Q���'Q��'�B
T��z�ܖ�!���]���q����t�m���f�VX:s��,�`�9FQ�����Ѐ�Q�K)s/��j�\���Q�X[	�r>�8?)����ã���d��P���9+N�f��d����r���[[[�Ϻ(TƎ�D�$ �k���<4�L!�E���-ף=ї�3<U0���]�NZB$3ʆ.�������|2P�
�����u^i��Mi1I5kY�*�k���M$�y����D�X����M�����0C�a.��gS H��Yú����5���e����g��AX`�,мX��.�j�h�4��YH�L}fu}����4���}�$-��
�~n=֙y��,��i����:J��\��ѣ����ٻpŎ�c9�L��V$R�8�I'A0]e�"��(�;���8#��������l��G�S��+W��d��Z
��!˂j�M�P/+���؉����;;;��dkFy�:���C���R�P<�őG#�e:hZL�x�6L��e
�"����^�H����4�[������e�k��c�i��F��ܺXf���9m��7�303p�M`m�e��y=�ԩ�͚���U:H�:j�c�3
;�l�af9?ZG���$�P�}]q�~1$�U��7��o��<�(��W�}��<+����,�Hɲ6�Ȳ��V�G�	�b�I�'�89
�R���s�f�:-�>!B�1�U���o�)��ҥKo^�zuo{{{K3��B�}H�����ɯ+��YCg�ѥ���,BB�K"���*e+˳6%AT�G�����$����R623��:G��N��:0��T#%XH(��n4�!�����,c7���Au���&�<,�>��(#����#��"2��x�4ȳ׎g�vq�nsoW0�x�'��y<��o��R��\�'jj�:2�c?���5b�ﴐ�=�;uQ�vu�ײ>�:��c+�+a<����Z8�v�������N���W�����]aƗ��B�}[��)a�-���_����?����z���}��'�̞@�J��h�Ȣ@TZ^e9�!�F��u�w�l�{�!�F���0�x��g�YUvoI�"+��=3OD�ANy$j-p��,UE�I@2~����k?`�c�w����XegT�Q��s,T͍L�xV�Q#s����E��y�il��d�Y.�A�^�!���s��1��<�ё��<��1��l9�:q�fٛ�k�������0c�[G�yG*F������	,�\m�SE��yd���,��)O���G't,��l�:>����'�d������O����n8>����p��zx����hn߹=�	Bk�J��={��A�@vi�L�?:�� ���px2�~8M�`r]����v��/}y��9>s�+�����⋿��o>Ua����
c �R�%'�E	)3�Bf!iŝ9� +��i|y	�}{{��%�����G,�0ca��dEs����r�e�x�j�jBU�t�,c
k����\et�b��<E���O������Xf]�Te��{��bdcz�<�SֱY�ū>�3�2�٧<J,X�ɫ����×7gD��rhRt���Y�>ڸ��{��=���0���{��﻽��g-��E�߽:7�9�{%�,�.��㱯M��?��c�v�,���� L��h�0l_8>�����W_
G�I�xovw����x��z�����Mǳ�eFY"��6��x5�O�x�~x����W��_}��w��O?�����o�������[��g?������K�~�c-�g�k׮����χ.��Έ�����L^�8���=!�,��G'd%��%ę6�2��a[O�Qȷ8d��� SY%h�a/
/AF:}�ܖ�N����4�p=J�������7���ܷ�R��>�-�\���~����y�i>Kc���g�e��e7��(���Y׵��,ë����u��P�zk}���Q!�����sh�0�lC��*��V�{�;�S$����x%\�z%|�k��_�B�!��"�.?s)\�.g'ӌ�ý��½��������*<��p��Q��;�n�������_���?x��/��{w£{��{?�g���?�w���}����7���}�/�|�0���?�������^����۷o��O�0&�쟼[+��`�C����V��X"�s	٦�Ȼܧ�i�U�ϲ�	�^��^&]���y�iy\���/^�t���r�]I�F�x�k�c̷����UE���D�5o=�^�ֈ�Y�<�8��,�����dy��9�,`����|�-����ǲ���i����(�[� h�m�	���u��aY�k/�[����ɹ�(�<g��±�R7V��x$��(+�b��`�������w×���l;F����v�p�\X��{w��͵��������iz{amm%����t'Av<>�}�w>
����'���Ã{w�dr��|;������7o����W���������~�?�a��/}i��k���7���������^B4ɻL�FV��V���7D�jt��k�aR^��c���/򀇑���蜂� ��kJ�zK��[�.�n^ۺ���E���C�sO��6�P����cE�zF�<�Ї�D�#I�4�mg�2��rʛ�,U��+Xr�X�9����>�^�><o�ޮN�����T�-��	]�*;Y��D�t����}Ȼ:g��:u�=}�Ϊ��~�Ģu`�pa���x�B��>���6F=,x�q-GGa��vx�ë����/���a�X[�6�h���A�xi;ll����{�g�޽�0^ݟ|��8\}���yp�F��6�CX��ǿ�w���㓰wXL���G/����7�z��_������W�����\�죏>
7n�|��4�{3�L�}KB5�K�(�%�LJ��cM�Aɰr4��jD�b��"�2������H���I���,����Q�M:�}IV�M�ܩ����j��W9r��x���Ӱ�r=U�yd�GCW_i�=�QrΒ�,���Ʋ��e�XbYm�z�'�jX�VU�]�m�Xִ<�b�|��%���.��by��>t_뱳�����u�վ����TQ^��D���ݭ�g�����P�qX]����¹K��d2�f%���'����=��ʕ���W�/�x1|�v�^��m���W�;��/^�E����wg��_[[����>�h'|�ʹp��+���I?
��C%a���}��������Nܛ�������z���w���[�n�"�4\n���6�G�~8���g�	�g�=�쳍�IJ
�{kJL���7e#d�NQY�����4b1���%/�2�v���o9ʮ��e'J�cHo��c�Rn��T�S}�!�u�$m��#�6iU�g�PS����>��}}�� �HE���%���+��XC�D&,���uNfڅc��Q�+��fot�C��2�:�H��"]]��Z�E��za&�q{������wo�����>acmz��q8>��{��h/���/����_t!�����3���O>	�o��}�+�٫��[?�<�q^z�p�ʵ��<�͛�^~5<�ů�O��b�|�ܵ�Մ��[��֛O>���_����'?��;w�|}gg�'$�D5����x+8´�'O"�֤�o�����}���o�=����ښE��q��5i�6��c�ͣ�s��� g��P�C&�����-u�sz:a��`^��N�y�"݅Ԣ}�o�����.���&A0��ҕ�����/�����g�5���T�zQ,�.Ui����y�cf�e����:$�e�9���0t�TH�>�,�u����'�b��F�(�tu��O�'��c��s���Z�]vw�w~�f����7������k�p��z�����^XG��W����o~)���vx����>�l�������˯<^|���ܕ�Yԙl���υ�W6������_�Fx��­���^�]�2�0+��_���ӷ�C�x�������ƿ���w�ܙ�d���3�F�It�D�������g�U�1�=�a!�����4K�Sih��Yt�'����o�YoŒ+��:@��5]�e�bú�[��</ch���6�2i�2��}ޘ�z~O�<���}|��w��$)�i�����P�^;�b����	�xq�ik�&�Z���Yvv?oZgXa�>UW���D�*C]?�s�U���������Z�y�����7�w/������s[�asmzoq��G�赗���F�|q&��¹��pac/L��G[�a-��p!��<�;a4��d-lL?��8[k������8Mu�n+�,e<�������^���?����=1���iK�X��At�5y�gM��Pe��u�1���H)�a�fʰ^�u9+�k~}+ө �4C���.��z�Zc�<���,��2�2�b��5��$�"�i��w/qa�b	�b�yuMߒ�g�!o2|:x��I6�>�ֺ����M�c�����F�R�����8;�]VW���f�zy#<�����K/��u!����a8:|N�v��h/���F���������������a��������h�n�y�V�u�v�w�p���u�Ax��'a2	��� <����\x��óC����+��}�{KcL&�YT�((7�F�iC�l��h�ѵ��޽����"�i$��{xT8д��>8C���Hc2g-V��[ޣx ���,�e�<0坵|�Z�J�E���HJ��.72�.:��A��)[�=��`1�.��`F��c?Gʴ��J�	�s�W}����1RuA�$]�3��)�-��icG@���L�Sg�V0�+��@�q� `�1+���`꥖2_�C��8�Jֲ��KTN�d�u?_�:@����9�2�%	�"����kx�~gg'l����/�~�?������Z�}t7L�,�	���� l�M�9��oO?���_����ڍՓ���.M�-���$\�t>�U��:
׮=�&����;�de3��_��ͮ?3��`Z駡dm;K�0-P�`�_u�9�� :Az|�E�ˌa)d���9퇩.0XP���`*����]R"̖	H�{����Z��x��=fTfF3�k�@ɰ&x4ڏ�\d����GR����ClanI�1"<ږ��&S6�����9eY��i
�(�Q��ti1I.&�h�&�r���"@e"��� Sas�&�����@ӌ�3}ŶN>�{Ŏ?9<��k���ac}m��� =���vX��F'��j8��A�}x6V.���IXM�;ۛ���O£���dr676�4�p�ܹ�8\��4���CX�:	��^'�a�x3lo�;[��t�Q6k��d�*{<�}�d"e��HU��
�~���1����h���$#�R%E-��Y���%���<S�0<D?`�ѼR�먎���:��`>?ә��|��4�ۖ��H��k=��!�.��Ƕa���D�\�1#�YeG窦`T泂�N������Ƨv�Xבߥ�K���Aw䓿y�:���G�On�w�y/�M����p~{=����x7���Q8��K�k��F��+�(l��������0��8�M���2}Mӟ�}kz����/��A�O�xU�YG�"e¬%�MNUQf���~&�|}֑Z,����#��Q����G���2�B��
q6����^vx�Rf���u�3-o��C���:�"��d�M�!�"�� ��c�A[��l]&@�$Ġ�5��눡e��<F����ea��%ˬ#)-�|(��q#Hy���+LB9�,�-�H�.�F������o�]�p�ν���v��Ͱ�3��c��sg:a�g.n��={-l��	ӻ�Jq�9�VF'a��&G'��Ͽ�&��k��4�+QV��aq!lg���]z.L�Vo]΄���Ro��8��v҆�p[i|���� �m�=�� (R]�e�,]�'����B&��a�[/4-a]�GyN3ǲ{yE���e��:N�JQ��ߣ�*�줦ˌ�`�Hx�e�̞0�>
�#��5?���̶cn�Ӊ����o�H\�q�Y���.|�L4�,�-H
���¥k�ʳυk׿&��akkVWN���v��a�8��\W��r������amT��sa�{o}N���}�a}r�Ɲ�u�u�z+�d�n�xP����b�|���2���b3f(�H��h�����AM1��Z�2�$e���������mH}�Id���fmұ|>�6��YW���K��sq��Q_.�l�`�U�T��}ʫ,c��ݮi����̨04�0UX�}��b�ga��S�eT��u:�(f�S1�Fێ���h����a&P�+�yO�D��v�q��f�o�C��̥��^�ڷ���|8�����=�Q8:ܝ��W�Ɨ�	���pp�0���0^�4;�lr�����v�&�Ga�x3�q�<ژ�5
�Gk�`ڍO֧׌��h#��[�0k�y[2�A_�`���;�oss�Rp{����4��3e��md���y3e�,��T~��2#Udݾ��

=x���{�x���j}��.���]�1EE�O{��Z���".м�2�.B�!�D��*ϋ�:���ˍ�u�N���h��F�U�u��M`},�b$iJk���Y �-�g��;�it{�����wy_[[;=/O�c��>>�܋��^
�~.�auE�Ɍ4#yɘ�^�nx���ƻ?�7���kW�����E8���_�]�'��[Az�Ov���Q���O���qx���p��υ��N?1f]QE�����(��Px���Si �z����ޗ��T��F�L��k	�����/��Z�C.��C�����S2ext�a��K�1<e��*���HU�b�u�u�eT8sG�y����>2)�(�i0���2�d<�m��aVt'���`@����M@)��&���`��51�0c�g�gb�YY7(�������p�ac�>��� D���!٤���8�����;�����Ux�o�:��Xׯ]���(|��������~/�M���,��/����p�ƇO���֥��_
��[��	3Ty�pz8�T�?�4�l�����<�r�1�G0�N�9FK��yTP����ѩ��(��t��\Fy\Q��
�-��X����P=�E��:R4���G���:��l�l`M,�Jd��5���6�al#��u�sZ�_q֔��m�V`���ؑ>����q�5&X�[3�n=:��u�����a�|�(��UL�P��b�L�U~D����$�������5^]kk[ӵ����iZ��k��K��Ǒeű��W�wq+�񣟇��ݰ>>
�._
��$<���7W�[<
����;am�W�l�������pR�{7ù���v�z8>Ÿ́Y�	)�^ﯩ�HcK#��/__�������D���� 6�kQ���VE���V@�(<F�0�=*���M��X�Le��B�����(걆 ���m��c�hyX�,�ɔ?�D�u�����<ȽF�,;��Q&Xz����yO��^���[�YºΙ�m-�P��1��rֶ+��k���d=�q,���m��6�*c�8qX���6F��W�܉��-��U����j8><
�n�	���0���a}��kڇ����� L'��ݝ�чwÝ���i�Ǜ�ރ�i�p,���Z�y�n��.>~��~-����}�Qx�?�<s%��_����>����r��^~��?=�Y���1[��L�2y�~�̲0�4ŋ�*�L`�~֕X&�x>o^�l��]�֣L�7˰�q��`G�1����B�hg)���ҜCP�)K�Y�k/lf:LX��T�J������	�r�b�s��G'�!�QFY;�Z�7崪�E�F6�� �(�=�a&R��"�~��U,�f��$W��Kb�z�k�'�_S�֎�():/]�ә���b$*\�4�V�S�s�������;������5��n�8�����k5��8�L���Q<�	o������x��,2�$��i�!ȵ+����^X�~1���_��;�O~�W~��}���_~�'��ʕ+?���_��_{��Z�L�P���4aF���g���㙑>�`@=�QXzĠ&���x*uiI�0��[]
���T�@��b�zk<Ve���u�k6�>�5qjI�3�΍,�g��f��̯��Kt�"�uŐ�E�A�Q�Q&�3"US�ɩ>�:����hM�!�H�!�r�<ǰ`=�1�c��k�.�9ƚĳ$��df^)�EH�GX�1��@��#/!��x+���.���۷ÿ��������嫗�d�VV��%�\$��09<	o��n������0^]��a��<�^7���q��k/�_��������7��9�j����/��/����l�	��P�w!��`; �'�@��3-�U:]W�Hl�V���`��.3�Üج	A�j,bm7�R�жc����}c� a	�~��~H�[��E˅�WR�c~�Lxm�pU{�-��,3-f��Y����& N'Lc��>���[/-�;Zrݔ��A���0�W�s<:n0�m,X}J�
�0C�ł̍�d���L����E��Z�0�`̵��5�0cmo���љ�v|��@��i������ݿv��Wã�A�N>?&քl[�f�vw����(��7B�2
��iz��8�f�ҥ����v�v\םg�^�^^R��HQ�mIeY�lɖe�qb�#6� ���1@�a���_���t?�<~H?�a�` �O��Ďe)��S�(�u)~\�K�9��Eo���W��Z������:�����k���'?����O������9��2!3uʩP�`&0��-��
/�k'��e
Ѕ��1{�
�:l����k�)����yc�X����7#���0�|�E�0�q, �Xk��XF�{��X�6�˼�s)X�^Ά�&�xK/����Eσ�e+++�y��q1X�Ԇ\kL����+�~�יִ�r�c�V���L��&������е ��3�!���}����$*�*�U�9�D+`�ˎ0��4�L�����I1-��[+���9e;����ť˗�=+�R0�L��2Bm�x��dVg���W�HD����{�:[&<+��o�<�H������g��_��=C0I�j�T�~J�
i(��2����m��C=�>S�5�X�a3�-�h�b�,�ک[P�0������Q0C=�=n=��Ћ`J��.s�a-�y�x5�7��n����>��#�XT�)���IB�S��o�p���ypS��Y�6=;:�G�I�|���h� ����s�gz�c(���fZh=���[G�Xއ�y����ի�� �9��<"N!0�]c[:���g5͌�cF����7��A�s��6(�Pˢ����������>hcc���e�'I�������Q�]3-n��{���"��-E0��=����8��\w��ؾqK3)DP�y��;��#G�w��7�w��#�9�T閌�Z[[+8P�߿����e�ޟq��i!��2�&�'q�Hi	S�C�Z4J��s��q�������[	h��ޢN��-��6���Ј��0,=J���\�=���d���<'ӟ�����5jt�u�m�uݴ��0=�Ygi#m���3�}���(���|B�R���[b-*��*�!�@��:@ 0��Y�AD<ݺ�
����Їb}t�P����;��T���n�%#��h֤�?�vo�TT_���3k�7�H3��=����ط�RL���y��y�g��#o��)�*���[n�X�7{��׋׷�w7/����ϒ�.�=C0[�j8�t�e�`2q����Wm�=�����
Ө�4T�� ��k�D�- �\��]1�:r/�tqϊ�b��2F�)˶�yXm� d�S�-Z�2F��!DC��\EԹ��"�[�k�<��0�w�	e�a���G�pNi"�(�&��	�x\����h�6�XG����n��D��a��C�LϺ]�6K�����=V�[��W�żϰ�[(֎jmǘy�&׉^"���/_.�\�Ri%���h����bg[��z���jE��3��7Dky�<�l2�S�?�7f/9�l���b�ޕBb�JN�n���#g���~�̖D;N��QuT
]�����k�A�����2���v��l�����@<.�
��sA��M0c����c�)�0EQ,o-�c�[��m"���,aX0�OK�����~����� X�
��k�>���{�i!g,�`����3�3�v����������8ŞK��˵�a2uZ7��0h��L1潘}'���cz�׵�O�}��}?S0c���}��DԊ@&;�h&�K����2-	+����c��,�ٯ��������=��Za�rs&�0�Y-���/af��-Q޳�Md�%��d�v�k�6�V+ƼmtQ��_��T��D%�-UTK�P�4���ZTC�؍�L<���kk��D��9�����+^��R�nZ.���L� �-��A����6�L2�;<���CB۶�^�C�خ�n���.?Ӽk+�M��ZǺ#�k|6]#�<F�X;���+��E��r]Ȏ(a��`�q-��'���"j�'��"��a�p��l�c�Ok4-��Y�^�����"��y�"��5"��{r���V�җ�-3�+����bZ�h7����ٵ��)�3��E��N$"rZ�d��/�;��.�V0�U�E�O���S�
h��*�]���Y^�w�B�3���6�h�!�,ӳ6f"af`-Ԏ�NY�Mk��c�z���;kϯ\A<Ç���hW&��>�h���O"x?�����Lۧ�A>�y�7�p�X��х���z}&�|��[M��=������1�	X�vv�$���uz^�#��J�����QL�:��1�(�߯�9P_i�X���[��Qu� "ݡO��Dv�K������b����g&+�d�l�8��?���[Q\�1-�d�Nnn�([/��&���}E<���]��i�O��ﰫ3�:���h"�K+���$�1U]O��,<zE3�)sl�cg��\�M�ə5̭N��<���_�D��麶����1G(#�s�!�)X�ɦϠ祢}�4���J]����n9Wd�o�^�~Y��,���i_Ƹ������W�"����Y?,�L1ʹ����@L�#��<0�>T,�L�}O�y��\I�R)�Mno�X��׭�n޵(
Mkϭ�ͫ+��/����@�f�su�T˴��頒V&t@��F�\�!�$��������Y�����Fc>� ?c?���������p�2I��<���>����G�Y��zL���v�Q<©I��^�3��:�m"QX�,�fh۟/#�tM�O��,u�g�"��7B0[�&����`��� �"[[�Gᔙ�t4=斚�3_���F���<_�V
f7n����3�nF��|�5����k�~�[�ݼӭߦ�k�yZA���T+�N��3�]R5@�	f�{��Z�S�[XXb-�Y��*S�(#��������0��,���k�d��о�j��˘���$x\��%��������Y��5�����0R"�׮�U��VPrѷ���g��.]���)U�f=��[�yM����bY��y:UǤ>��E0�f��e�Cֶ��#��<g9�Tw����}�����n�*&itY��D絷��}�馀V^U�1�T־>�`֒���dlJ���y�l�,Mx\�z4 Ȣ��[a�=��ܐ{y˃&p��L�kW���%�~=O�ҋ��D���,g,�=�o�:���3�S��3! "������%,ֱ������z����%ބ�!{V吰("
}.k��m.�a��Of�S��¨=�1Oj�PӗPY�Ҵ���i+{W��{��[Y0�y�MM�+7k,ߜ���f�Oo^��n�8�;L���YGP�lQ'U�,z�y�[��VL.��\5�D�e��0�@<F��c��G&/�s}vģ�3���ް�P��@\���^�u�՟�@a�#��/��bnS�,�V��H�h�C���Z&���t�|��5�x�<>�`�U��`��H���E�3��󵿇|d��Q�c�;�X����}F�U�r�G�f�3����;��)�1�v��0)�a6��~��$}Mo�n��̖`���*��wgU<��hS9�w�}��=vڹ�=a]��I:�`�u�5f��o�,�nF�����c���^z�~�����m{m���m�l�]���#S�A�3,Ј~K������V���y�4����6�T��z£��d�sS�xt�f;#�Iσ�����n<��9�mX�,�!��ٟ�s�_�1=GvϞ�m=L_�$v["������tR���9��/�0kCfA�Z��fu�$U/������5�<����[�x Y]��C�ǐ�4�z�y�us:��Ia��u?�ʅ�������c���y,����F�T��c�d�2fXm�ݮ�d���\�X���2n2,�s�X����3ϙXo�k�V�:��z��yu*Vrs����i GUȟN�1�d�fKB��i���묷������yAG���p���n�Mn��F�iL�/$�D�M�[bY�ZE�?����Z�i$Yz��D-�Ɠ���3��}�{y4�z�j�-=�D�i�����M[�Ӊ�=��U4��F۞G�5�y�+LÌ�e�����.��+&��/�xS7�쫬P��f�����v�C�_V=@aE���X��C̃-�\w^a�#����#;���볼���P��ɢ�-ۃ�3�YGdz,vz����M�_���t:�{$2LU�Bߟ�"���狛��'�г�Qg�[��l�5-E�m�{�z���@rgg�V�_]]-�_�~�=\d",?�����1ʵ���sEXg-� �i=!��Xzp<z]0ӳ6�YJބt�����7�S�3Y�=f�u����t�u�<�O��X�m�xl�H]a���>���]��Ft�d���ƍ��XG�;$ ώ`-`�=�\a3�������9�s�M�����l�{��׹b�y�\0���^�3�[�-��e9vGb�(�gb����ԃ\wdh���k�s�ni#:E�~i����KHu��+{1��=%��|��AI�?����l�}c����w���7f��Q�Fڹ�fx������2h�K��+���/���$ }&ot��n���b]ϙ0D�6��XԱ#�����!ʅ�0`;�D��db0B���3��w��f:��B��:Y�5~Q#���Z�5��9HH�7!�P҄�Ȣ.��^;z_���m�e�\__���uϸ��Myv�s�����񼉪]��s��%?-a�;�/2�C���5���VFz�v��ٖ��B�S�,,{�P�L����^L�s u������w���-V�yݭH��oit�}�n�U6Ր��HN3��v�����.zt¤�UP�UK������\i�5e!��$��;��1��\0c���Ȅ���m�;�0��x.k��v�k�A�k<noͺ�-�ZΙ�E�����#s��5�:��YH�%s��\[x��(��i�߿�����'�xF>0�LdE�2��Y�8PX��s��%���J��g	t"V�ڕ�HX�3f���v;f�Q��㪪�j�j٪F"�mq��7#�~��_������!� �T����bsss�P��6f�Uk���G�R�c����d��f���L,�����ɵ�x4yt�h8�7�5�<�n/cj��[I{��A������Z���Y��vv��/L��ܧz�<C�0���fλ�9С0�V��n�(�6m�1~0�C�(����-}n�>�㚗y/os;��Iǆy��D"<%�H&�%b��$�X�hT�-۴�i��?��R�S�4�W~n̬=t=.B�.
.���0�;�gDN��2�[�a�dF�14�h��T��f��� [2�׿�j�k��+�6X�\�3ZXs)�㬵�m��k�h]W���b0��fM�2x\;Z�ӆ��[F��u�`�2�D`��c��Ta���1�)g���T����﭂�F��`��3*���8����hK����]�����.x�������!�o>���`��w*˭��C�&c6.Z��B�E�X,>�T�L����{� Ј&���X�U�>�Y��u�5���ݢ�Cf��"�NZ�
 ��G���QŹ�k�c�e4)������z�Ѧ_�&,��f"����8�����\��j�Zc��������YgT�3�l�p���D��նȵ-X��F	���Zv� �ţX(9<��4�Ep�>��1�/�m|z��<�bh�u���ɀ)����B��t�1��x���\��ͧ�H��H3����V�����������)\����8�����g���!�]0c1�m�z]=��f"��V��F��e7i�rMz����\��&3"iE�����u�}	fm�e�ӢyLx��{zcƫX����/��f��|�oA�d���5�e�ݴ}��ͭ�f��Z�k�A�6��<��5�doC����&�|�4kX[�yt�J�[j��l)3#�������'�m�u/4�����/3�\A�l��9G`�S,<������C�<�����V�"���"��&�M�KM��<����9hX}*��k߾}���{�N�z�&�&�ޔ^���C��2�陰�=�۔�e>���~�g�-�����ko/3t_�5(֓t�7�%^����sk���>^}����	���[SY:a�B���Uzm֗��i�efE����E��#
�r�mX�m��;�Ў�`i_��w�5,����� �A*���VU�d|_]]������/uI����fWfh���I����WU7���or��t]���/��z��ࡓ��}��'^#<X�5�x�����"�v�l/��yL�=�V��eTb���t�v6�hҼ���4 0~��c[`=*���pV{Н1�����o���$l,���_˶��_d:˲A�C��y ��mGf��˃�;!Ch#Q5�S��f}?�M�~}�{�l��u�帎:�uI��3���rPb�f,�.����Z��kh�kz.نQ�"�PtL��eNw�ڵ��n�k=�*R�gTMF�Uv~h�O�V0kS9SESNE.�t�Y
I�R(���Rj��`m\Day��5T��}6�`���Ǜ��W����"�.}VtSp�8�A��4 �`.�,bւ}�}����@��3r�R�(�2A��Ɉ�Lq
%<���e{h��,Q4��!ː����M[��Ms�0�뵱��S�e�9S��^��9�W�k�B��5=D8�Kk��C�q-�b9ǵvFX� _�a<ׁ��D/��
\��ا�˼��K�p\�]+�-K��R�L��toM)������r�թ�j4K0[���IDNx���za���u�3=�XԵ�4OR��&�<�3'�y3�Ø�)f�a)8�*����5�{�Ϝ�b��k!GWXώFޠ[7�<ȝ�Ll,�@Pr�'�},TL�����N�d���zݣ�`�\�F$0ϒ�X_�vʨK����q��G_6O(C�\f��B���
:E`�bu��b�Ω��C�F���D+��~��-�4�i,;����җ�a��T�������gNю�/#d��2�����:ek��hl����ã��m<�	*�0�|v�u��z/�B�ȃ�Q0��9�'�h��ulh��'z��\~��Aa�W,��Wv;���W�m����u�5�b��٫Cn8�N�LGnV~vmW�D���:�u�K��y�x,'	4�X�˄yO��bae������f!�2^�~��PD �m�gݲQ��u��>�`�D:��FUq�LB>|[1��%�5L�E�F��`�-
$wr����L�y�sժ�W��\�,�y��aF|Y���(z� ��sS<���h'�]0�ji/h���f�5�9�τ�5*�:��	�`�4� 0#���cֳ���7X�@C�Hz����Eh	�|�!�e"���B�s4�5~t����O�#pӳ3������l��&k�I�i����W�>����:�"j�C��If Z������KH�a<z�ha�瘉B�m�8Td�"�"A��"#��zq(x3�0?KOIt2�Q0�H[+�ë�1�1��Sr����5�ϵ��u�ۼM��n�^��x3�1a ���f�g�x����&D{L�)`���]k�%I�B�EH���Z+X���e�%�I��~�z@�K��v�B`�ǎ,j�t2/���F�e�P�w�q�ٗ��a�cQ�z�6x��ma�Y���>3]���	|��K����E�l �ǩ�Z�0�-=n�dmC�H@&^]'�D�y����#�XL�hk��&�������\#}_�zN��2,A&��ӂW�ң�Β!�)�`��L���C���`��w̅�5�s��;yv���`X��)��뙐HC�K斾H$�3�e�C�kkkн���Z0c�9RWX�7h.N�M ��o�jJ/�3��zn)���m�s��1�uֺ�3XsD0C�C�;�9gM�Y�{��	��,�Q,�����uK�U1L�����;}���y�����eL���dDZ��Z�[[[ŕ+Wn�Z��"	ӰVg����-'�h�|�n	�&<�:I�̤/kjW�H�s�f!˰fm0C���-#J&N�Po�ŪLQ&"��nCg����^P��r3J�yH��,���%֎�	��B@�x���*��_��_K'Iٝ��!A����ѵ�G�/t-�ދ�2z�s֎0L��a#A�i����y�}kG�>�]tfĞ�5:�g���Ĩ�w���F�I9�e�sz�٢��T�fZ����*�:)��E<����(�|&�ĺi�_ט�͌gbc9I�X/��<�5��n@�b�0j��Z�=z���(�B��`�=�m~��^^�hK<F� �ޢQ,�L�9��;k�z�a��L#3�>
�,�wC8iYG���v�b�V��:��c�Cb�؇cX���N�r}���Mg�&����y����]��}=����*?nQ�Dıt�E��:q�j�\�]%�ifJ!�������﫪-�b-\5����w����sySۅ.gM��q!�]�`=��sx�)}N��|�͢���L1E�ǠN���	�i?�,H����c-���L(�Va����^ƈ����^}`m�F�f<s��
���󘞅ѥ��A��2����op�K�����@�8�K5�6xV��}����)�������sa�/�|[;���1]�̼v?��ћ��%�����)�i;��X��'�)��n��ډF���"�ez]�����5��1���}X�U��,Ӷ� n�{ h!hhp��H����Ȇl��g����:�>��uײ��R�t���k���(֞X�Bs��B�F_0v�����5󓅇g�2�U�����gB��s�y�>��ocB�iN&>�,���Q��x�σ53=�=
o,cz���^���4�{��,�f��Θ�\�\�X�TX��!�'�K{���-2��E����c˶ǎ�C��x/&�c$ہ.��k��AG*��e���&�}�zW	f��N3	U��:U6%�%r��=obAA�Z,��s`�vAA>I��4�H�ӟ�KH���[��T��[i�Ϸ��(��** ��i��F���ӑ{�AA6�X!�AAA>T#�R�,}ա�1�5�{W	f{��)�!~(խE(K_uA�+ad
� �˂�u�Y85��� � X�T�R��5�I_��������I�W������:��ݻ��/��ݪ�/Qe�WWWK�,���h�I�K�#�L�K�vu ~���3�s�1=&��� � v����,��b�墼��M]ԙj;U��nGA�qbK�9H��
fm#�-0������bkk��9� � D�Y4�$� � �#�Ҡ�T4��,t��������scc�X[[;�>ۮ�VVV��fmS��*��=��+W�W�^-.]�T\�~�҂ r��o�Ȇ �~	 � �N�� � X�j�X�$�_�kee�D�Eg����9R:t�U��v�`&[2��^�!�^3��{�bss��$�,� v�X}��MB,���6�A`z�E�� � ��6�Y�Ţ
hy�Gd	�`V�A�n+F�����/<x��|�J0۷o�����ˌuR2M�!KC��=/���i�Jt��e�(�����y�Ο���|��;���&�L0>�l��wV䱌'N�]�x��l�}ԟ���n&gq�r���a�uָ9���L�{���|:��!�*>�M��2!�2Sa-���b�\[=VK����V�8q���~x}�]%��q��=z�;����r� Qa�T���������=�$P"�Ο?_\�x�˪�eUu��of���kp��`�\�`Q��]��ϹޱZp��=�L�g�	�w3�ɸ�1�ShZH���X/2P����3c��y`�:�K�Lb�ܼ�Ű�K���|^f	�n��]���y�[&��po����+��}��~��6٘���2�Z7�k��ҟ�¹T�tKE�3�V�T_�#�D,ӣ�4�)E�2�{��E�ψ�s�ĉ⡇��6Ϸ���{��~���Y[[��Ν��+%��@)��R�0&|�ڵ�w��5v�VAAAA�47�  I}IDATAA�S�]Ҡ��g	���EXQM4�QP�?v�l��j��w�`&<����:y������R�2�P� ���T,�@���ZA����MA����ł ���]��m9��yҔ7�������P�%�F���G�-y���ӟ~����:��駟~������/���b�:���"�Ię�)�>������"���e���AAAAA��T(��h�/�[4�11i^����S��j3�$������x��'���yv�`&<��#�����{��og�`���d��.B� � �t�Ry~�m���fT� � � � � hGD�A06�zA��Rm��	z���/f��:�ۜ<y�8}��_�җ����v�`���}�;/�����7��aY�
�d�fZ��=�*���,_��-�&� � � � � � �l�S�$�#=�L��]�t+F�Jߓ�(�1�#�H4���v�`&|�����~��������>���g��g��K~�|����2ٖQ5!� � �Jx�AA����A�C���!��2�c���j3�R�-=K#���2�]�b|�'���#���.v�`&���={�?���?����N5���^�c��§�e���V�͂ � � � � �`wS�c�f�̋4�����-�X���x-�_�뮻�ܲ��k������z��3�Z�L��������/�ۿ��~�ܹs����C�}@��̖��"�����A��Q"�'�qAAA`A�f*��ޒ
f��ȫ�����3���w�]<������g����ϰ�3�w�w���Ç�����ՙ3g�-�=Z��+�b�L�K�K9�L�o��Ј4ٲQ"�Dtӂ�M#��:Ԁ�k�*�B]%gcm�<�KW��h�c>����%��˽)�6��0��ߵ��<S�'�'�g�-�^�-�v��O�y�s�0�؏��}�<<��9����<灜�2y��J�m~�]��v�lz�@�c�����w��/}�U}��ٛ�fz���;R_�}vH�m�U��s]Xs�.e��u9�y״�مS�x�]�c�'z��-'ۤ������@$��\4�I�9u�T1&ڌ��ӟ��x��o2��JM�g�)���/��W��K����}�cg����Ӭ0��������f��nyV��d�l�(�$���Q�q��r�vJi�_Ty���$�A�+��A�#�_����A�2,Y�P������<m&�+�������I��3���ů�ʯ����"z�7]�v�<^K��m��R,�����X&�z�Lx�'^^__�?N�<�7?����_|�QQ&�$jL
@UT�,;r�H1��<�L
lgg��x�bYXNN�mXY��"�~0Q���L&QW�D��vD��Oݙ6N��,����u4��%�f�1Mw�K�$����"AL>�`��O~�`��$���ٳ��r�h4'N�(>��l~�_�_�~�0�[f���G?z~���ɓ'���~�'?��W_��;f��ʥ���ʖ�(�f�7Q2�����euLb�����井[7��A0^"��_"�y��[����*�Uw�K����%9�����Ł�w�y�x饗�����ޣ�>*Qe���'?����z�����Y��|�3ߕ�_��_~����[[[_�-E�QL�_�LD3Q:�w)(�?�`�e9"�,#Q�� ��;1�A�b$�E0	a"p@]=������or�X�FU ����+����w�С�رc��"z��/Qh��|�������MA&T�9|�����'N<����G���We�EAL)�;��>Ox_��9�l��-/QO��7�F&Q��e�[�m@��:�l�DoD;�I�j�y��n�kyl{h?=d~VE3�0�4�RME~��U4�Ev����c������K���X�@f8}���s������Ͽ���/�)��Ię�)[1^�|��?S�p�yBY�Ƕ6��@��n2�6�����k:r��$�o�L&1�
��D_���{A�<�8�w��f����ܔ�e~�ŉb�3�D����e*�齮]�V�;w�x��׋�W���e�x��h�����B0k`kk��ƭ�
�8�B�L4)8Q9�f�,�AA�<t�� � � �B��*��(�-�'�&/9
K������k��.�e�k~�ӟ�B������u���
���Y!���B�=2���W�)☞i&�X���0� � � vu�a<g��K��x�^��1M>�}��f��,AJ?��ϋ���2�I��x�RH�+W��,z �f�D�I��ޘr��ɓ'�{ｷ���(C�z�b{{��$���V=�L�Iã���A!�����u��<�<��W�x/fXoyk]~���D�I�i,=�s[@�����ȧ�6Üw��}v]����]ⱞ�\�}�<�e�;��������{՝kV���X�'3���UM��߬>w�>r�2��sϢkLK��"�i`��t�E}��"�b�6������΁�B0k`V(�"xI��@v�ĉ���p����!�kkk�?��?������?�V�	u�����A
k�N'A�{�djD�djd�uJ=Ә�A`�$����e�Du�7W����1�L��7�>�dDy>�쾈����(V��\�9R�D4�x,�4�nܸ���+��>��������Y�y$�q���2�lV��ӧ��%P
N
Q�n� ����!6�`�x����F�E����� |3�yhtT}O�d��%pIv���%�L��z����om��h��YZPRQ5�L3�.^�X
fr�YfAA0�L��@���Q�%?	�,�!��� �4*<���:ȝ1��tG�T<KE3�$pIv��]��_�^�k��믗y�g��Af�
iU�[YY):T�u�]�H&��r�����o�AAО\��0DC�=�&Q̉<��ʅy�yAA�*���X&/�a�;V*�.w�qG��
f��&�Ha�{i�{�X�A=cM�L»�J���6��A�:��+��9�M&y���"
��D�σ ��e�)�4����mQL5-&�f����I!I��;�S�/��իWK�S
/� �2��m������ܢ�.D�s�ꖌ�/󘄡=Ȝ��>�<��<ȝ1�a�n�0�[677�.��^��\�r�Н E��k��YU&!�,��k����v�gϞ-o{{�� ���Il�8vƞW!J�2����[b�͐�%͏͂ � kv�Z�1V�D0�x�bq�ܹ��w�-�������W!�50���gg�T3�z���W_-E������2��ڵkEAA��Lv�X�V[�$TMB4� � :��WU�K��K�.�f�ϟ/�&ڌ-ݺ�L����l�(f"�I����F�r��"��ߥp�@:!ݢQ���AV��7���;���ϼ\����c���޻z�b]�C��om�c�su�!+Xm�+H~"�.Ȗ�9�>3k��4d�z��Y�LZ̾�W�:ӵ����2��Fd������3���&��I�`��c�C]�)M�*4���A�~�rLc���q�9�w���5������ٮX��(�>���c��^���[�������	d݄�+��τ�Ŷ�u�k۷,���O����!נ�U�x���O�vC9�j�K �\���z[Xӝ o]���з����Y�H�H�]�~�ʹ��3	���P&�-���tZ���s��V���j,b�@a5���́������ւ�������!τ0OD���	j_�y�d�Y"O��u�E��&dl�N-��#i�/��>W�6�^��)�-=��s,��e�f�	u�e�"����-�������Y��_]�����$��JL���L�gJ��yu��uE�X
f^��*��R�����3��n�L�#�z�	�?h����m�Rw��q�Z��s����̘0�u�����o-�!��V'ºz����-Mi���J�LM�m�{ڎ{���Jo�؉T4K덖��'���ŉ'�{ｷ�f��۟ΟVWW�=�Y��� ���(�>|�,\)<�6��<'����f"���Svj8lΚ@D3��޼��tY�-��E$s���LH��z���Z0k�T˥�ޡ�˅�Z��t-'��"�e��h���:7�M����@�e����(�eA���&��ϩ�Ϣ~(u0Aӛ��Hn�o�9²�B�@@�M���2c����~�g��3�����e�K�s�5Fӳ���v�4O�j[.��� �zF.�G���c\�ߑ>��h�6�����
T�G@���	����uF@V^!�k�5Dz����.�Euװ�ܣ�m�y�lf?��0�ƽ���U!��)�z�A�ӈ�����M���MI�ж��Qw_$�t��E�̼t�>�ܻI�lJGi+,z̘��"� [.Jp�$8p��X&b�ɓ'�ӧO,�H����^{�5���=�Yg�)H��첻ﾻ��R�RPr��fR�Rh�ɉXv�С�=t��ļ�\g�D@&B�� �isK�K�	sQP7AC:z�>},5˘�&����w����1��Ь�˘�Tꞡ�X����-8�q���A��`^~ �:f}�˙��e�`Ā]����y�<Kާs���~yo�3-+t��m��:A�r�'�%,��F�6x�suuL�r/�0�Y��X�x��іE�5C�l3�J��YoM���P�E���U���O�ȑe�C`;$��C�qv�F�4=ۢ����ѐQ�Pе㢵�>3k|D��9n�>Q;E�[[¼{����1u�k�yn_�zkLqL�~������K�D_� $�z��رce�o��V��h���oD���^�K�4 )УG��N�*QO�9w�\�)`�$�z�N�P��6�eD�yt5�+]'�]\�	8r��=���=��>�Y�Ff4��Qu�}���g^uxX�.��6�1�L;��U,�
Z�u��̙������N��Um�e�q�sV���b�_�Wu�����>i*�~��l���M}�6,,�E�sw����5�Q0c9�F�y'¼z��g����e�c{2��1,�>�L]��y��fXb
S�B���Y.,P����U�Z/YN���#τ
JHzlqcY���'h��g|�[OTa:����s[{�V�{m��E��$����u`	f�z ډ�_�&�}����Od?4�P��\�zAti����\���͢B0k����/���%&aRXU&j��Б#Gʟ�,3�����9)TːEV��u,2��{LO;�:֖�,��6��̘�ҫ�g^]c�EC�fMT��^�+=DL`�g)�0�Ӳ�\m�f�R�,�SF�[Ԯ��O]`,*�0��CYm)��:���<_Fa�K�u���|&f�W�m��3m�{�:�Ѥ]�C���n3oa\�<��5-?��s!t��x 1ȣ��uT���g�2�B_��2�Y;x��Ve�)ބ�jzm�V��g[��d��JS�q���u~�^��fލ.m��mҚw��X�n�r�u�tYc/���[�����Q0q���˥n"�����*�W!?�u��r������~���x��G�=z����GE0���ڵk�&E
Q1),�T����l]EﺀO;�E�`yb�)(y.,TL+r~W���4��`�&�&�#��j��B�d��A�/CpC׼�e�ߺ���,c�����s����wy.K�y�6ױ�D$z��L}���ϱ")����{�f]��`=/E@�)�g1򪍣aS]b;-Z݋i0D�K΂�e�K�\����gb�)�2֢��R�@a�-T�dD?
�g����|��ѴX[��C�i���=M�qͼ4��eF�������Z����(V٠�˾��}��x�H-�cH��۴c�3�ڨh*o��v���b�Y�Y�2�W�o���9�D��{�����3E�`p�ȑ�g�������3gΔ�e�����{��&�%����	�\'�-ږ��Y�	��������sm�e-� �X�gf]a]ׇ���#=�>%����{u1�w�_���>3=�y��}Ku2�g��Zϭ��.y���ϰ�M�1�1��A�kf��e8]�ˢr��e
��V$=��V�-o����Kĳ>��c=�8P�2����Z �A�:�֑�֣h0��d܇%�轐� rk��������1h3�-}���N1�1� �$��b���B�R~u���-���]����]����'M�	V�b���o�Q\�x��d7?=Q"�DKE4M_4	b�v"[5>|�բB0��)$Q0777�������"��{��j��N���R����;���_3��5� X�}��xcm(`y��8�����Ϧ�XN��b��SXީ]�¼�������z���2�`& ۹1������,cߢH4�LY�����Rց�E�1��H��<�e@n�Om����l����5rXv׶��|yY�5@���6��qE�a���wz]� ���JO���b܇y/f��"nt���0�M�ۧ����͚�bE;1��d�xm���D�>׎u��]�rA�?m�`MQR�]�,+ʴ|��X�9]��"A��=b�3-�����-�:FZ��uql\�SD+�������}���2yO��]6	\�,	r*z 3������lJ����7�,N
S�D��v�(����iR	���� �)k�����m���}�rB���|� �������vׄ�{�F%��(kqNhۮ�֦��}BӳX{@J�k26=s1wQ:lP��u���;lY1��9V��4�is/�>�q��qM��Ƽggoɸ(�.,ۗ#X���l�h�jP�t�)�jf��-���4h�%����������P�,��<̹*�ZLq�%���(Хφ�ה^״��9�C�F;5��d��W��F;n#� ��6�Ģk�|B@�i�5���>;�%��[��?#鵝�/���ٲ6�4�L���2?d�>���+@���ٳ���w�dDcD0;|��?=��G>�o���?�x�uي��W_-I�L
PM
M
QH	�Sޓ��h�F'�RY��0Ifz�YL,�̺ߖ���}{�t5�&=����0ɜ�f�1�l�3����A`���@�=�m�zq߇�Ā)V3��+���|B�u(kJ��ߡsEƼ;��y�dK��Ͻ9��y`}^��ڊ96���|2W�ߏe#�v�EH����M�G�R��
�)ue����8+,�D����ٷ0�����+ϙ0���Ƹ"�1���y)��t���tl����r����=	ND�D����[~���Z˝w�Y�+��[��ԩS�c�=�͏����B0x�駟�嗿��/����z�ܒQ
X�i��{��w�H2Y�K���)��%�L�3�ʹh#F����h��^��#k�Ǵu�hk	��F����>��ּ���a�S�`.�r�,�hQ��q�㞀~?V����yq
��P�&XX������k��`)V��&�޵I�
�������c��<R�����2��eި
fu�6��w^tH���u�Lڦ�b�L��%	��Z"y��ّ{!��,�s�!��k��w�{�X&e�Qc�$G_��r��W^)2�F4����g�g�<�Hq���������?��3g�|~V����9w�\y �D��&ʨ�)�/�Ie�������L��N���3������g�鄀%��9zT�i��]̬�֑��2�4�O&�6�y����h�+^�.9?S��n�'2�b�<-��CoX�v},�e]��˺}Z���΁�3��#���9Dz�X9������k���>h�X�v�����X6�v��ѫ��XG2y����z]h���n��m��{�5���`�F��V� �N�-��,"��6����'��}�s_;}��7��!��H�߬p�ݬ#�����>��/�>�L^RЪ���h%�����j@P�et��#�RK`uD��j�ͼ�p�4���Ҡ�H��S$=og$���o�҄u?����̀����["�
*<!��x4�%n�ۏx;/�sx���QM0�$��1օ�nC�KK��������*ర�~�X�1��D�>�"�̋0Kf�#�o�av�`�c�C&k\@��f:~XoS��9��N$y�kǴޤ���t�E	2�L4:�k��K�.���p�ر⩧�*~�7~�?>�����n��=B0k�l͸�����9��~�����e�
*�3�ک�a�� 5��ӊ�
f�ƕ����d���:�:�H;��@�P����W]��� L&��3'���B��H[G���3k1�y]֓�1�(�a��W�h�tѳ�}ֹc���	�+z40�Z�ߏ�� �+c���`�s��A�V����=c�}bW�x�h�H�cwfg��Z�iC`�Qm��V��]��cb-�����G�#��=�����r�(;���Sv��E뺜w��Oz����߾��/~����YK��W����݅=w�ܧ�<�T%ME/�Z9u�?ݞQ=_�Ύ��f\�ok���Z��fV��ǰ}K���u����Y��cE�Q.m�d\��0챮������`.f���N�!"`U���@��d9N1眖�CtY�hZhD"3MO��}�F�hD4=�>cSra�A������tD�]� ��Qtm���O�?��,ˑ��t�f�S>�^M�߂�S*��k}_����U�hr�
��N�*�}���h!�	!�uࡇ�*g�}�{��#9pNB�2�����M�LR�4�P*	�V��^D��1ޖ�0��:�j'��k=ba�ͨ��(�&�����w��Hg�L,��c�+̅�}�"��[�0�k�g�=�m"���\�2�I��hXoe(���qkR'��t6�.mx^t�yn�;;1�#�������`�b}��%�N��V�Z�5�,cu�J#����!�K���=2J������������#w�u��:T�,��y+�oj��CE��%�L^Bz��V
K�v��'�'Oӽ���E����~��)k������;=�޷9� ����[l�֟{�/�3Y�˅���<`T�0�3r��.
�gB"�P�����u0a��z��sVLF>oc3ǜWM��<�(��G�����c��C�Y��=��b�Q�M0�6^#���kU�S�#�k%�D;�m�%Z��(���鵚�����v���s���|��
#B0����Jy✊]����T,ӂNQ�vss��]�.
�^�nو����m�F� 5� ��{4�!T�y���Z����Y��6�z�SL��c �)�eL���輂^�\��Xu��ٙ^�L ��M3�O
�^��uӫ�c���B`�Ĳ�0�6�z�̃\�5�>�c���4O {��<��B�;-cD<\6=k�)&�f����/�;;�ڱ�}���Z�	�Ei��LG �z��Ym��Xv�ڵR(��{no˘�k�������p����C�ПZ~��:"��o��o��C=��.\��))��������v�R!~��/��B![9�{"�iȡ~ І�4
��)�k��!�]f>1Y}���k�Q�\8��a��\�L�����\��� ���<P�)Kѐ=Vy3F3���ͣ���1�~t�e���\�����s�s�4M�5(�DC�z��&V3aF|Y:�1���,�6f0���22.��+�X��<�uxQ=h��t�܆Q7�|�\��<����t���k=��o-Բ��`�U,��9Ob;s���������'�K4�e������c�=V<����=x���眕���Ύ�>/����/�:u껧O��faHfK�|�k?����{��7+�յ���ܙu��J����*Ǳ�G��ѥK�>�R)M#д�[��ض���O}
f��\�6�)������(_F����K���,�7�>�m=g�>^!X��L<-� ������C�(D���6/e�������6��_(,��<b�f9e�25M9;[�`�H��O{�ۤ���?�x~�v�kF��8��O1��ڈ�}
dm��&N��Yd@$�9r�x��G	@���>����l�=^y��Y�\�}����3���IfK��C�֌/��u�o���{饗>?���,=�L�c�E��>���LCx�3=�-�d:�c>7��Z0��h��'/B�=;3ϭ�D���`N��(;v���8k�M�(��Q8e���8�\�r�����q���>O�~�a�E4�ר>���������z���t��N(��j��m3�:�Bw�A��閉��o-V[;1M����i��p�?��Y�Wc̬�b&}����2�bo�-u,���.~�C*�z�o>����<�=���&���@�`f�s�=���}�{����_F�pԳ�tG�P�!�������RL����.�b�V_a��ìSL������m�[}a	fm�łU��m���4&X/���P�n�czV=G�	�w�6mM0ۺ��]���G�zo���Yc�����v<�3�ǹ):Y
X#x��x�d4�϶f�1z�ڱ-;Vz�3����H�وޫ	ɧ6��*��c+rkK�6_M���\���R�Э�����zM~��E4���;%���e^�l �?�������;��KB[� ƚ!F4=�fM����+h�Ek"��s�:�<@���;�i(�N%�am\B�k�u��yɊ�`��`mE��\#�s5���/��QA�5w�=����F������$�6c	�<���7�/�ѐ��)�y���Шpk�y��b}~���@,C�E}�!3�鱄����	A�(�&ڈȽ��'O[nߢ�e������;4z����ʝ)��A�T���ի�T�f,j�!����l8p���S�R)e`c+�T��Rґ���,��"���;�ɘ�e< �Vz�ɠ����U��b:$��|&�p�������^L/:����)�rn��r�������d���d��(���m�IX�0�h K,4"��L��<����s��ƜŔ>��m}�gb�q��s�w6Q�3��km+c��m��.߯O��Y�o�}���1�u��ޭg�	���}��'�2~j�ַ�`6 8{�С��ڠt�@<��F8D�����0�̼"��p�ѻ�u/��S���d�`��{�����:3=���W���^�xt�`�5Xb5Z.Hz�k��C�q�j�)�1��
��y��GX� ��2�������iЕu��1=��Zĳ̬�̶�j{H=X��h�Ko���Nh�L���{Wf�+X��r���!����kдX������6^F8e�E���~W	��l�x�Ȁ�`uuusmm�E��#H&���b�PA�l�=�2!X{<���t�ޒq��
��-'�^�C��%#�e�Ɇe|C�C,���[f�H԰���B��Ggֶbh[�y,b `���9�mo�������O�Hukc&���駐�#��Cʸ��2��XG��u� � ��c�`:��c?k���s�W�f���p�e��'Y���Ov�W��Y���y.�wHz��"��n}�t.�������r�8_��� ���K��J�1�@�~C�d�8�
}g�aLo-o�}��i�!�	?[�e��Ft�zgmC�
jdfE1Y��Y� ��X��d\���'�[x!0�:b\D`�?k��P��a�1��g�Lc�u�/zk.�T~^�C��!���[o=j����Ƭ/�3!0�CE���� `���3;��d�#���q[�{V�o)�3�C�2�9��CB:��W,�w�uȸ�e�Z��7�/�GB0�k׮���,�%J����@K��T"Đ'�k̰R�A�����Fo�qL����VL� ��m91a�M�nRW���c-s�`�X˸�.���D�=����,�b4=Ԙ�r���@���Yoǌ`-R"��e!�۸[�y�?`~ֹh�:�Y�^��i+%���g�gF����V�a�X0����k�<�"�z�gb
��s�<�x����Y�0�z]��k���.'�9�~��=ۦa-�Y�m�L�i/�>���R�W������^��-�%�l�:_d@f���u�����ٳgK�L��L��D&�B�Fd��s�n���--#������K�(���J�c[��w��"�B�q/kG�yπ��J�K��Хi.b��!�Rĳn{�¢�0� �|f�	K$��-�!"��	Ěy�<}�-�[�nX}>��� X:I���^(�ve=O��54�
f��4�����m��*�x���v&��KۛW_�B	�>s�Xw�.e5����G�I-�;�,���x��2����'��I^2GS�C������l �{�R0��&{xJ�F��fc�m�L�e\�{஻ƛHɜ(H�gER2��X�C�6�&-��+���~�ڳ�����yn� ]�$B�?D��uvL�E�<�\X�y�5˺��o�s�P�6c�b�G,S��G#:�u�!�L�3>��R����Ϫ�H~2EJd��Uī�X��z-��k��]�5d�!��#�B����4부���h�&���-��i���)d"�!�;Y3 ���vj���aY�Ʈ��\�k�JKH��4��`����Lg ֜�Z�c湥s�bn�<j'�g� !m�����E�`6 R9�]�rE�g,'�2i����26�r�	��g?�i��J&M�$��Y�t+%�A�]&�x�<>S�떥�d	i�, ��6ImXV4�7b�*L�"��an���(���,����'�߯	԰ς���'*��;��
tM���fz/�3�=CW�?o�Ú<w����������k�m=�X��mD	+�gZ$J �m�%l�g�{�G�̋zO���H�Eb.����}O�6�\�yL/W��)�[�9sΉ���-�8-�K�Jt�}��'���"B0�;��ջ���{�J#g���@�G�G���L/�\'CR�XXO��k�)3T;�a��H���^E<��*�3=�=p�����N��J�b�协���-�tj��v�f�DaE21%�f�]����bݮX�	d�`�Uz/�!�z>��>S]�!�q3�B����>8g�P�ǙԵ��k�>{��+x97n(�g����E��6�x�
f�>��:�uS@�,d�g=:Z���[k���i�g9���ի��Ɔfϟ8q��"B0�����.D4�
$g��{z�t(,+������1XX0�L��!�I��j��Ud�((1���Y���s�w*��J�ע��ϖrh�c���\ ��2V��y�<.�Y��tҲ^�"XG�3�6P��u��u�h{�G�8���f�1�9ר֗:A�[�B�T�4�t��f��1ζqY6�M�ᴀ�a�|�Z��M~.��m��i��+��	kgD4M暉i�c�c֙i�(��a�Z��)S�<�}H�ّ#G^��G?z�Ȁ�����w�v�r��T ���h#F!���E�Gþ`�\^=�{y���r:Tpa��}�G,�^aF簌oLoQ��eW5D2�&9�Yxm��F��$oс�eD�X�Ѥ�(BV۳6���A�p��C�	�6f[F#��`�GY;$亦�Z�F�1a�?�y7��g��=���-��M_�e"�Pt��(Mk,���a�+��"^���y���"��. ���cǊ�������?��C�e�l .]�t߹s�3gΔgmm�|_��h�Lo2��m��m ��9�)Jx̘0'��<`���m��4f2�B���3����1�ޢ��0�����Ggk�u��tº�|��t�֮к���降�"��(t����gZA��m�%�:�g�9-�Dt��J�I΂�����67k�uѺM?#�A���}
fuiZ3u6o��5�A�W��Y6h�|�H[�L�V�%����,x��g.]����O/�	�l �����*Hq���r/�}���V]��Z0C��$�C��-���P�4�h����<>�W���^�L� 䙘�15 ����$��n��u1���S{����y��k�I��#sL�u~��g�x�z�!��]F0CA�#�>�k�%V�����)m�c���H�#�&<FV{��1�h��i^�W��;�##����W����X�'Y�^�J��n��2�k���ڵk�{.\(�\�r��,�cVIv���_x'��`��Dk�=M�ՠ=��2� ���%kO,�h ���3�쿟ǉ6:Ae�Y0��G�2���t]�����i���"@ӳ�����#0�F�>�R�`F\0��h5�܍;�+�o5����GѶ�<�� �w]Ӛ�'=�cr�̻&���帇��k�/cG"��9#�rfٱ�k\��s�.ѺUڌ��D�y��b���Yf��%�"�G���8�c<�יi�\Q�e�^�k{{[3��`6 �Jr���pq������K�1�=>GS�f.~��r�^Aa.�X���y�^,�X?��ߣ ��s���mŘ�Lg�,�w�Q��uV�a-��\��S�48�Ft4�\�2�aF`Y
fhZ����y&����^�m'�13����Y�)(L�/om�=�2��g�l�̲����|���s@o�L���&�:�Yڠ��y&��{��X�0mR����V$$Bٕ+W���~\�|9������U&G�/�l�	5�ᠠ�ޔ��	hٱꔤ�xpX�y�;]� x̄��u����^�]��m�A�>#�)6���\Ԅx�y3!�1V�W�1=�Z�m�)$0�4��m�Rn�9Ʋ�
��c���n��[��s[c�̾ӣ33���1�i�`��f�p��������WM�s\֜�~�w�|o&Y��PXb�G���>��'�'�q�>���{��w�u��w�Ȁ�@�0����x�buu�̤�==��{�∥l�(��<Fٱ�(��a�֋m&���"��z�`-\X
X�S녶��{��A�2BzWQXN��PfZ����:���Pr~�&�~�etA�0k�BT̕5�L�h�]�n�?�6�b�U.��/��6k�EY���@̨,Q�ZLa�.��Cm�Hݴ��Ds����YfR7d�;{o�Ȁ�`VYV堻W^y��8���e��~�z�?k�u+��k�C�X(�4<Y.�s���/�HC&C��C��ւ�-0�(RZ�2
2��Ɉ�1*��㬵�ͺ+���G�*v4�>�-��Z���㖷�5�yaȽXyV�c�Qo�o����W�E�2A��ۘyd�y�ǾE�Z��o��+XF{��իp�`=�zǙ{�(I�y+`A�.�e�%� �f ���Q��T�>���3!����l_�z��L*�(�Z�d�FQb��Zo13��c��!<8<�X©Ǻ���z3趹�?g1�'��Ek���x��$߱!��Ns[�����Q��ƣ�8����:������b<Z��r��d�c6k�6��l-X
�C���=�M=�-#o��v�F��Ð�C����zϣX&X�-R�Dې� ��q�:u�����ƙ"B0�}��]��2y��*�G^R�D<C�Ee��^�,�F��u"�bM1�3��7��xۯ�q�7����3&�q/�|�^l[G�[އ}/��+�F`3���!�k2��,���\�:WdX���#orݖ���,��������v�m�Λs���ޣ@ǊPB���g��� ��O1����#
Z_�����ŋ��r����/"��Ç��^��� 9r�~��2<�w�)�;w�\q���r�lId�I8�$=W�����5 Z�=T��w{�,�z\�y�Z(A���^��<n��\#K�Y�X~G��LA����]��c�!Xu��w�3��W��n팀�5<Fwzź�𘟬v�[�����rtV�XFN��l=6��FZL�鱶���:ϙ��w�qGUv���bmm�܎������G?���E�`6 _���Ǭ���O�����|�̙3�������/����ay�."Y��.ox5xZF��C�Q��S�ο���E,��k�$"�����-����:�]/Y�5�E]��*\X�9:�f�#���3�wH��[�4�n�?�������ۤ�b�;0����;�:�fD�ǈT(a��i����:ly����<nъ�Ǻm�M��ΥP�$��9�{s~�8_Fa�;dN-u�c�X��3�l�Hv���2����V�	!��s�=����*^z����s�=r��W%�L*+b��Y����	��Α�s �\�"��6�k�b�3�-fr^l[z	��G/�\k֠�v�պnZ���2A񸵈%C�p�2���1o����NH�1�S�6ILP�6fzMx\�0a:���M���㭐���Y��b�F�՚@����b������1���J/W�7�}X΁�8׹"s���ZN`=w���'�x����?��o�f6"YJf�pğ��'�ߏ~����$H��L+��.����� Ӡdҍb=����g���!��τ��+����'���ڇ�m)0kޜrƺ����.G�����X[f0����n#�#�;��o"���G7�����u��:Wģ@ǌ,��*��<:������z�0���G���eߒk�3۞u=G�c��X��:SU��s�2f1̺���K���������&?��!/q���oO<���U,B0s¬��s�~�(+��d*��v:�F��6*!�<�PC4�Go�yi-�x�z�U�@A�嶔m��X�Q�^�F@x�����ɂ�Ӡª/L����m<��*�Y��!����uL���<
��_h��}�u�2z/�Z���$���|�f#A�c��<:n��6�3�����s����(�1��(�&�tl@�e�e�y&�O�MȚ@fR�B�
W�\q��nCfN�U�َ��7�,+�T2����/?_�v��^���yx���^���H���=Wc�G�������'�4�E�形O���!ڧe�X��Ltak-�xl3�L�P�",�sx����}rf�c�$�x�L35
F���5��D�Y~G�hR�u��|�U�IXbsM��q�-B{�4d��!|kk��+$�G�
y�]~c}}]�j�Ș̜p���=����իW��/��w�}�eܷo_Y�_�~[D�F��)�=?����Y�4�����Û� s��6i2@�ڿ"Q�����
�E;1�-��<
��b
���1��c��s�:����zl���XG��j̴��L�]\���̭$-a��7�?D��j�I��TH���y�}ZGN1۱�����,X�A΂��a2�J���gkkk�V!=z�|?~����{��^QdLfN���>��˗/����z�So������}������eC�V^�n�Ȃ9 ��X��iH�"P����<
f�WA`����- ,VIG��E0۞������L<>�8���,Xgдq�����Ǭ���s_ǈG���^3�/Ӹ�{��3JX�9���P��)N1�i�Ck��l�Ş����hZ�L����Ɉ�Q^�Ո�f�;K,w�a�e�z�՟[;wX;3����c);�O	����w�ԩ��'�<������Ǐ�p�������g��Ș��/}����U�ɟ��W���o���ٟo��vY%�Q�k�
*�g�pV�<j8D��Eu^'�����qq���GC�%*�5���`�l,�(��u�ۏ0A�Z��Z�QD�o���\M���,ga삙%Cx���s���s��L�%�9�5LOm�z�,�`�
},<�;��Τ�\�	S0c]g�L9f��=:R䚗�1�y��;�_M��I���w$��sd���@�n=�s&h��X+��Yeu���_����_��_�N1B0sʑ#G^>t�������"�I%��2A*'�M����#:2gu��\Mx�G�|&�I����z�<&�3�"S%���)Xo����a�j����N�"%+-���gb�am���B$G�� ]�[�E�q�ɵ���	�\��z/kG
�@�0ujxb�h=hg��e���Z��k9k�У0���� �)J�`��q�`�Ԅ�ӭ�`��&Xs�!�Q��k�u�\�Myn�'�Xz��������+++W���S>��O}kk�_>��c_��|}}������Y�\�M��o�ggq�kVfn�lwVٷ��DMύr�sl�ڃy�x/�{o��  ��8�7���W8C����Ŭ-��&�����k��Hz��v���e}A�	�~�%H�����Gкb��� �w�8k�uy뺕��7�������<
�ҡͷ�o��	�-�ϴ3�K��\��<G��8W��+�rac�n�q�[�bͻ��C��7n�#�w�h�Y0�Jz:Vy�S�LVz��j����ڌ{�M�꣠�ya��u`��&���;��{k�Jyv�2���¿�׎��M�~J�����U�������<��g�}6�3˪�_t2��8s���+� � � � � � ��*�AAAAAAA���,����I
    IEND�B`�PK
     uK\>B�	  	  /   images/687e948c-dc0a-4fdc-b588-e952ae529de1.png�PNG

   IHDR   d   2   �5~�   	pHYs  �  ��+  �IDATx��\]h\E>w�f7�ɦI���4%�Pk��
���>�m��!��`|R���**R�/*����Ӽ))RZ�*�b�(�n�bZ������u�vg;�ܙ��1+�	��9sf���9g��ܘ����q�������D"Z�e���"�:Yn������/cu2y>��`iCC�p,;��f!����ŋ��������|2��Jv�s�RvC:
vJU<1�_2� �0������dzzFGGaffZZZ�����-�:�I�?�s�|:�B@�,H�ӱ�N�G��ǻ��B�ϟ?d
����;��ē�]�2��� d
���ʅ�dJ�=�Lq�����֜���777?�k׮wm@H�`r/,..�w�WU�%S��:}c��)N�t�����j�(��0��$�ۃ�x<��>�/�؍��	�:� s/�v9��B,�/ˬA&C�p8�@��|����я��#V}}�Fz��K6�y�qk���L�qO�wR"�D�Vt�10M��f&���\��ve>z���!��@]]��l*�t�:��>��Ů�d
�x�);���ME`M��y*��#U��z_]d��F�bW2�������|����:�CS�L�N�n�\���2��S>#����<��y�D��,��(X�X�N� &'�����TI�����H�>�4C*�����@��&[S>?��C�@��0�$*S�(S�=xҙ��.����x2k��0�D���im���%7�ٌ�֩���݊�8[Et�P=�N��$�5�yDKc2f8�~3�Ll5�F�zS�#��Uw�"QH�R�����̵`�Q�*�*�|�,�� ���#^���G�7����{ߏ����o��O�;uY��yWU�kLFw"�D�x��N��E+�i[[�G�`p�x�u�$�0y������d�>K_,R3���w��'�W���W�0e���"�1�.��������=�,=z�/,�����H$�jgggޯ�Z����F*b3YT�sR���rM�x�]�tnܸq����)<P���76mڔd5�+)���B����z^ZZ�s���0����^��Qje�����m!r�r1�n�&Th�H�J��H��
@��n�\�b!eD4�؀�/�*V���$G4֐�1X6 ��\+TZ�a`�c��K�
���nU�z��H�
H�m��w� ʇ*��2���*km�Fe�UN��!�˲�R��_��[�V�s����S=s�?Uـ�S���d2���իw�MXC���l��s�/v������ݜ,q��~�eG�R�=�;���~4���ajj
N�<	�w� B5�P�S��b���ܙEQ��vXY�wj�s���<� #�� �Y�!J�o�<����k׮}k���ٍ��ۡ��c���˯��H��9��s�D�/,㰬⿪*�ϣB��KMMM�]]]���}�.q�̙{�~���U봉8 l�ۓ_�P�FgE���ɗe�����a�L�D�[	�H�0顸v*D����QSSC�
i��32�ae�����Q)�?	y9�/N&n�2���S�a4��87�tf����e�ŬO,Pb��Ո|��N���l�\��bYTX�@Г���dJ¨���#�+��nݎl˔+k禎^�+�3Y�,�������ȤHEqU��_�R�E3J��t�ҵ1Ս:��x����ۡ��xԼt��S�p���חݹs�d������
a���qMn�R���k!,U�邨rU�2���h���T��g�طo_����*&K�C��e���tWMNub�R�L�Nr:1�ϗ0��ħ��ϧg���|b�:u
�?�����dG�����/D����<VvCll2�XY�N��G'<������~uKA �}$y�~MQ�m�����<q,ʪ6�X�n��<Oei*W�Y�Q0%^��Ute����Lt��}�E8q�ı���W���� �S���u.Jn�� RY�]�T��1���}��˓!�������ڀ�߿8 �������	�=D��4p'^!�:�6�rW��a��.�J�x�����#j6�7o����6�'K�Al����+ç�ub^$E�Y���N��YY1��cMɾ�3�}��T�F���7�W'_�X2@�)�E����g������`��}�
g}۩П�r��u[��KD���Y�v+ds)�a�%�ķ��x�$� �t����ϭ�5    IEND�B`�PK
     uK\�c��f  �f  /   images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.png�PNG

   IHDR  �  �   ��ߊ  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  a�IDATx���|SU���M�M��ޣ {��Dq�����~�V*�~���(���(�"{�Q6-�-�M�{�'I�M������K��{onn���cU{�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!����(0�� t""���NDDЉ��B :Q`@'""
�DDD!@��-[a츱�aC�5?�q8�^ݺ"���0�
�"���l�a���>C��p���Oo��vn����"��mE�9F�1\���?ۛ�����(:���c�X���_wlP(�ʔ{���=��|+��#}�Y��mo�w��k��]�o�������?�O�0�?���'�Q���W?s��3��"Sڶo�dՊ�}�I���i�f����gf^�t8Z������^d�g`���>�n�q�0K���k|=Ϗ���5�1��}���I0�p]�y��U��'3r��~'_{���G���ߢ��h������1o��v�#�����޵{�I��z�}Պ�ged��x0'""��!;;�߁�������t8�ADDDՎ��4���N����E�l4"""��L�����QQ���ԿTP�UK���	���sn������BDDDՓ}����{�������H/�=��|!'""�c�4a��sh׮ݔ�#F���u�}�?_+.q��p8PPP��o�O���m+�p���DDDG�}ǎ툯0;+k����C���PA܉��\��+z��I#<r䑓�\y���O5�Q�?�^D��R]�]R<�5k����q֦=11Q�s�*Yǖ�Ull,���0�C�Y6'"�`V|֠g�HKKS�o����T���Ύr���������GXd$���(T�:����=3+Y*��D�~2+3K��H�h#"���sx���_����`:͈�����O��;r��"""
f����6.��p�)�ggg��oDDD�����R�7Mgx�'�����"""
n�Cii����p:M{�'��]��QP3��SSѼE�8���,�3�:gOݟ�F��:�������y�
�DDD���";+;ơzI2�kff&���(��j����H�4�L��at""�`&��:���K@/3�^�a�Љ����nC����E��J膻��0���(���*w�^���(@VV���(���*����:��D^^>���(����p�Yo`� ��;w@/;�����FDDD�Mr�0��mPP�ϵЉ����iB��'ԭiՆ.������Q�V�%""�Qt/w���^J�&�΀NDD����m6È𶁴�{+�Qp�/^�T���t""��g߾m�*���6�Q𲧤�H������]��1�'���i��*w""��g����m*`��r���/��Ä�m�����NDD���3��G@g�;Q�S%�Æ����˝��(��3�����G����ΐNDD�Lس23��i�I��S��)U�ge���'{�3{NN�
����%�;Ճ������zdDD�i��K�DDDA�T=&&Ff��Н*�;Y�NDD�L{xD�t�S�:M�~Q��l6;|T�;�&L�Љ����=L��*w�Su"""
^v�a�ax�&�܉�����0�QN	�U�DDDA�T�\J�׉e���U�DDD��.K�|tV�3�|�i�̽t�U�DDDA��%���F��8tV��rK��U�DDDǀ�����t�K���˝��(���K�z���X���(��E�{	��7���t�,��ʝ��(�ٝO	�:��:űʝ��(hI����4�r��YB'""
fv��a�iz	�n?7�)���(�ٝ�sm��NDD��r���SQ�n��^�n��GDD�쐕�L��T07Љ����)U�J8|�r�Nq�DDDA�n+/�K�g@����<����@=?""�F��0;�*��乸ҵ033ii��k�.$'�@jj*>�����9	�QQ��S�ѨQC4k��6���\���1%>�|��%rpq��+�*3��?V�Y�?���Eb��-طo/<���<W�C=��,|��\`�!6&u��C�V�ЫWO0 }��A�&�f�1�Qȑ��i[�I@���p�{�W�܌���X�z5���;�:��V�ޯJ��(��Q�w�{�>)ͧ�Ė���/s0i�$t8�#�=�\|���ܹ��v��D$<�����pU���Ʉi7`��r��s�C��\�U�^�x1�����n�n٬��E�ۆ�)����`�E���Oq��W���GR���yv"��\�g.~��w|��g���;п_?�i`7нN��¹�}�\�-[�b����Gcǎ�p�W�����=轢������i�O��P\p���������O���u����拓�'�S��o�T!����>���2>�͘����3������_��p���T�Y���tf������ذq#��nԉ�cP'��'������ix뭷�|�2]�Y�^�z���'��2���V�{!�Pz^�0���*RS�µ��Gݷg��g'a��Mw���������{���#R�۟���#G���x䑇Ѡ~}u"
Zy���7o&��f͚���8��yHo���;�1��&��ޔ�y~&M�\�f��`�
���hܸZ�h�:�E˖z8Z�*UGGG#7'�z8ۆ�n�:lݲU�TU�[�Z�QV�a����HOKǨQ#� 1�A������K�,��߁�����Qi�tn��lC�C�����g�><����!??�oF׵kԸ1����3���&M��v�ڈ�{o���b�ʕ�a�:�~�:w���Gf ?/~�$��'�@LT�:�Ca�^��,���eʐ�0���or�gf��_�G*��`���9Q'>�>n��V=��v�Z�ϖ�|/C:�5i�H?�~n��L�<S>�\��S�5��s���[h׮n��z�~Y�(�2+&K�"��n�f9U��W\�Á�U	x���s���Űa�p�9�v\-�_+Ƴ�L�׭Kg�;��|2��֮�ù�J������ѱc�ؿ?K�DD!Nt�s����!�{Μ_���~�2�M�!����#г[7�_+O���/�	u�b��aX�l)�36�6��ѥK�� "�P�c�i7���*w]-̀^�n�ꫯb�d�z��L����p�Wb���hռy�Kƞ��u�@����~�H޶�����{�	�_xK�DD!ɕ�۝�i���q����0��)���_Q����p�����FTI0/N�}�Yg�����ǟ@���(�/3p�@*�y�m�4` ��cP'"
9�����rg��#���,F�9Y�.;ѵ[�G�M�VG%p��,2����/�L񲕁?���?���%]""
I�L�곛�k�Ԛ]B����i_c�jo��L������ރ^=z�R�'�N݃~�os�o�X��3��0s�L�{�DFDT��y�"X�X���x�����X]��:Ne��.��� ״������͞�}���[8�2{�u@|�ٸ��K�ɲ'8�w�{���O��������m=�c���xbP�p�ٟrss�����f��u&"B=�ߞ��y�v����y���Cn^���OV}���a+���N�[�8r��!�1�(ǲ��V�Nq�|����EFxȹʵ)p�>[u�rm��ץ���u}]�����OC��:����9�?���"��\}��ˌ���^��Пc�{�hU��)}>޶�R�5RT�y�s�C~J�@~�V�,�[9C�����57"��_@��U�?ϙ��+V�ۭ%cͯ��zԍ�?�7�/&:�^v	�M��C�0���-lطo�-_���Y"v���X�vV�Y��6`��]f��S�P�,�B�Z�ШQ#�n��:u�q�uD�����JZF233��]ۺ		:�*�>��)�f���X�x֩��s�N�I�##"�{hѲ:v�^�{����k�}^ŏ�r�*,Z�k�5۵k���t@����36o��{�@��]о];Ԋ�����u�8��W�3K��t�	�H��r��!���Q�X������u���lչ5m��}ջW/���u�9��a��5X�p�>Ύ;�q$C�����M�4E��ѭ[7$%��k U��{2��3-=[�l�K!�9n۶�))�����C��(�OL�3A��E�ΝѦMk�V���~�:��.�����MIJ�)���+T���6mB�>y��zK�D��f͛��,�u���㐘X��ZT��gVvv���}<p����_�X�����)�T��21g�(��t���k�8t�(���S_om�&���O<�R�>}�]}�������֊����m����ޭ{w�P��螛�J|���f̘����[�nEzz�����u^��t ���x�s�98��S�P%���w���x���٧��U8r%���5l�/��2ڵiS���C�o������
+T�g��>އ�";4h����õ�^�A�����8;U��n�����/�l�2���w/�k����(u�p�)����N>�$�R�ؑ^�/���<iR��r]d��_��*Hz����ᇙ��/�x�b��>>_�͎z�����5�\�s�g[O��J��`��F�ܰdrd�$���q�#T�T�9���u�	�$xUU��\�M���5�'���X�d����Hp�uT�.�6P�]O�ё"��*�W6�{�U�~1#G�ҁ�0��j�L�#�<Rbd�<������ս>Uw�MNNF���zoR����Z�.�1�sp��#�}{���� ���'��o��H׌2*��ґ��,X6�����?��v��#����.�С�)��^��C�`�l�R������;�ޱ�A.ǭ���*�4h�=z�K1�tP���>��U�ɫ3U[����{����z�g����t��.��c�JXd:ܛo�Y�ʮ'� ��%�ϕ�X��$�9[�
y���N��r��z�8�ޭ2�|��~��^v)U�gR�ve�]�b���ٳ����:���q�*w{�6|���0�Ǚ�Zɇ�J�͎��T%���_��u���<�+�ȿ����_�sGvv�_�+�lʾ��5�����y��ǟxݺv-���I�����B��Z�'_�.w�ځi_}�9?��ŗ\��{I����'g�k�|���z9ϕ+W�i���-�����nՏg�T���p�������KGb�*����?�{���K���Uk���̾R�����'[[��>'�dIAa����G��o֙)��L��M�����Z[j�֬^�u��T&��ge�ԯ���(g�pKU0߽[� �=�%~�q�I�������5�گ�GZ����[=�m؀�^{��9N;{$�6%������/�E]�r�Z����5�m��֩��,ǘz� ^U��7����}(���\�;=���}lٲ�����]J������7'��^��=�ܯ��5sm�?5o���ά���:v���)푆V*4u��p����N����|���f�?c�u�!�_L�[�n����|��"�>� /���]ŏ��VJx�n�\��cǢo�^��r&�9�UeXe�sU�-//��<{s][ɠIFsŊ�駟�裏�_����2��-�S�-��⟩��]x��gT@��&��̊ٵ�̮Z��?���H,���>��I����6��x���r�#����D�Х�2���>���:wB��m�Ӗ���[*J>�9*Q{z���믿�^�)��2�J(2���ч�R�J�H<�!C�v'T�%���'�x����d�k����~����@?���B����3�{5j��4dee��2?E�q80��oUf-�Ox�<�$�*�9
o��ffT�|ſ���Gzo�3�up��8���J�/�_R���>������O���$}�+S%57�F���Ƕ-��f�x��r��0��iذ~=�}�\tᅺ�_�SXO���/�£�<Zl�)��m[6]��������۶n�NjA@�����:lM.��t�t�2[�зO�׉�:�\jf���C����໻����m���WJ�Y��d��bX�w��_�h!��^�����_���*ڋ�	Z�1�w����a�B^���t|߁�'U
�4q�Q��-,���1a�J�=U�9�����NJ��= �r]���1��W0��	�ζʼ�������yx�����K/�Nco��^;i(��?��@���u�ȑ#�h�#!����F����9�[f��zH��������|���ū��s��z�
���zg㪫�
�gYڌ�3K�b�c���+�������Ǚ?⥗�cܸ�������eR:����ǝ�Tk��g��Ѝ�bz͹xť��`Ϟ�^����B�.]t5o(]!OR4��Y:t6o� ��ê ^�~��8ӻw4k�u���UT�h��]z���˖��]	��=gö����Ï�k{�E��T�ק�~��%���#"Ѵi3�B]Su���7';�R��Ҕ�n���VS�JЎ||�ɧ8���|�
_/�]	hLl��h��m�"11QG����uo�;v�;�Yg|�T�H��E_�.�W����=u�4LU%9W{y���D�=M�4Vץ�>o�$��RSS�a�l޴I��[_W�2L�:_r�
��0�L0w]���u�4G����u��n2�Jz��]�V]�dx_�X����(��N8�_�������ȑ��v� ���N��B��I��K�.�3�����Qڵ7oެ۶�'|��C�.Fq6=���=�;�^�I�$��t�2L�<����\ރ|O۴i�{�K�HG�C��r�򹦧�y9w��LӁ��}s���c��A>�G���}��/��\=�7mܨ�[�d��%�ף�t�S�֭[6+��)s���2>�����ak2�H!�ک��H 5��_�|9�?5��`�Db���T%�W^y��#פtu���ԗW��M�:����k�Nx�;�oÓO<�F�h�8Ce�Ru tu�+
�R��ۯ/���J�v�ih�����̈;)q�P�9����oM�R�1�f�Ϟ{n֫���]7�
�u0��3p�:N�޽Ѥq#=��s9���6�k\�����}{���#Ìf��:��^��"�>R�s�v.
�a*A�ޣ7�P���[�j�;W���W�dΤcۤI�����e�	�34t�x̘�طgRS���v":�N9�\}�U�qӦMu	�s]dH�֭��ݷ�����W`���"C�O���}zW����3�ǘ����yp'��o�駝����,���!�1�S��߅�����Y�,2K�s�{]VN����y"����}��ΕΠի� g�u&.��b=�q�ƺ7���zA~>RTfm��%�����H�Qِ�o�}�]�pB=����m곸��{p�-7���]���;u������gj��Q#1��u?�Lɐİ��?��kf@�R�+���D6Х�P������*p_Ub'�|*~�a�q�@Ĩ���'9��x��W�������6g�l��X��mX�z%�W	�۪�Ѩa�J't�P�\��T%���;q뭷��JPQ�L�p))�҅<������>V��t�Q%�����[���x��Gq�E��P��8R"�ݳ�w�'��?��*SeyUR��N�m\�а�8T`�*�G��"�*�ȃ�Եi�Jp�+c�\��-[��u-q�
�R��
�e��B�u��l�kޢ�=4LW97�_��K�jת���ҹ���N�ñ��?��IUb���{�͚4���^֬߀ѣ�ww����'�n��s�mh�2c��:��&������Izʿ8�E/�(ٰr�r�S�O|�Mԫ�P�{]�냅�Q������O�Ї���멈s�m�y2��|�q��aʔ)5r�:�����$C�j�9��nE�Bf��Gq��Յ���2����4��>A�I	��zg�'�q��ϬH�Zž�b���u���1}��qc�}˻C<��&g<�[��c�=�i_M��8B�)�|�ɧx���T�V�6j�Q�G��7�Ꜽ���R%����믿�vxz���T��^��K�DwZ�VaoǑ`0d�`]���۱g�.��lܸIWG׫�$.֊�K|ݺ��8����I����[Ǥ$<���X�n}���H&�ƽ8�{��1ͅ-���?U�1c���nƖ�-�c`��d=#�t���a�ĉX��[�թJ��1b�H]����ɞ�V_]O�II��V�	V��3f`�*9ߦ2��Q��J��u�_��T�3�9?o��!�Ho��]Z��~oSKK��|��:��^��X锸��Zzj|j^�9bz.w��멚�)N:rI��+�['P2�HL%&�6�i�ܵ��.2K5�u7p� =L+�]�#z�����J��t5���H{�|�ǨK/��\gW{�C���]����ݯl'��I�ᤷ�*wk�.=��`^ѡ���:^t�:�D�g=6X�z�J�+��;�w�q��ů"ץW������1F�t}��H�[O<�.8�����{��N��T`�>��C�aݺu8EmW���]���-��V�e��O>����+0��g���L{����t�{�+6��hˬ��z(��g֥〥)�|��a�葅����h*�I��K/�K�,յVs�H��c��	�N���Ց]���g��m�vM_d�p/SfVWs~��ŋ�[0�j��숃���V�ǞxLw[�'�([)�l~��ttx�� u��8��tӍ�ڸ��A�L�������mE��ύ7݄s�����9IIpР���O�x���1t�=iK'��֝�RʖL�ۓ�Fj�>x���J\~�e>k,���*�O�4��C("7JG+����S�#S�Ju�Ν�U���|�M�A�n+̋�Ƌ/�Pw}a����$C}��1�����Nt�p�Zb���W^#�j�G�)S�m�U��y�f�?p $k,��Ͱ�۳�&��KG���l[�V��P�i)��~��7�Y��~i�'�T.��SN�|;�����}�}�a���k�������s7�p�n���qM=%�u�]W���:w�&M���`��G'Z�l��.��2:$�~b}��f���A]�&"#�����)�Oj�V�Z�:�y�xm�>C�u�Ǒ���w�5)P����蒤�NS�*	����2��:wŭ�ݪ�D��.���o���f��.�+K��e:��^�\���0��$��a�k׮���B�{��]��Cꚻ:�ѱbJ��M&a.GMkC�_:Qe����B�+�ۄ�y���$\q���L��OI�.��=��?�:�X�b��5hr�9�<����uĀJ�엨J;�u@_�u�SO;�U��� �p��z���L��U-��V�[a���+���ؼE/S|��s��ǣg��*�JB����m�uQ��^�s��Uj+�2�aa�ͼC��z\�ަuk�{޹z� ��ҿ�.�M���[�5h�Hw@�L�kO@�*yw��	�M�n����̬��б�>k��]/�jb�db��[J�6�`�=D���3�:�[�
h��Kz��w�y�c�UU����0�!�^}UB)=g+P"UF�a��^����r�#��.N����72C��- �>=z�@�J���u��$��ye�лO�J��/���KH��uY�C:�z��(���3o�<����^v��F���,u��x�	i�8p &�5�G��ۇ*�"�Kf�c����(�;YAN'���*s��"1tL�v���u9�����M�>f��ܵL�*�W�L�b���:2ɔ���B�F�4i}�7\�c,XY�K�}9���B:]�t��{��_�׶BSO��1 �Ԇ���qb�>/A+�g��IV�mV�5�ef�U������U+Cw2S׿V-�m��zQ_v�ك��Vx}�k�nh߾j�Hr7M<����J&ϑ9�s�n��^r�ש�������"B���VMcNgH��Ւ����yU��n��sTt�ϭ$G*������٧�`)Î��z�Y���j��ڷw���n٪�l.=����� �+KWT��{�ԓ�4k��e�����H:�1u"ݮ]�J��}]t3���A�?�l��%ǩlgTڶ�ː@���;�`0���I����K[7o�|�y�w53+���m�Fe
7O�d�$3lU�.�Ռot4�_˫r����$ш�Yb1��4W�Ȕ���ɬ�i�u}TsV��]R�����<�b�0��;v�eJ��(qq�t'�ʒ�k�')=���y?�u*�픡��&ޛD\%t9Ve�U��쨌M�7##����=\��[Uj�_��d`�e|v�ڭgᓀ~dLDFE�q��Nz%�*ڼ-��b��/�$t���g���3�I�!���*s�I[]%�Ƃ��͝��Y��4C��I�oU�	��!+�Ig$�6:�t����W+N=j��IЊ�=�Z��k\�V2TU-Zer�t��*S)&	�nݢ�}�H&j��=���_�HaS��L�*�Y��?x�S�W�8��A�@L:TD������YCg&~U���JJ2��M�����۷O�U�w��`���4�eɼ޲�CU/BӴi]��(�8��;��[��.�?G��X�(U:�N�H���Q��H�������܇�}޷G��YO�����Ǐ�믿T�o��ѽ��z�����d�1�F��(8I	�^4o�L��]KJ����MWz]=��i�suj);�7�����/�yJ�99e�2�:Oα2w�T�JG��&�;F5J�$�v42 R"=��M��R�&��x#�k2��q6e�&5��؏�d����j�k�#�\m�5�m�Q�ƈ�]���:�i{�w��`&��[�M�*>
U��1���Idsr+7,�nS�+�����]M��W���e<���X�����z�Uѩ��jH	���n����dLm�zu�o���.;�Ɂ������O���V��G��*@Ib���C���l5s��J.�J�*��<�f"W]HG���e��@u�*��d�;Y����r{��jh@o�X퓒�F�3^�kv$Y6P��7o�3e5o��u�`>?��>�P`��+\��U���Q�*��SNUC�1G9��qk%�Nӽ�0���pk���a��򎥚�gϞ�V�;���˗/׳N�`��ʒ�F^}�5|��7�бz��޽{��%�KOfo3_IU��`)�hf��0HR��g=9�!c��5>�'
��L���C�v�\�3G�f3u���@T1�Yn���5��^*�K`?�a=fu��eض-�:f��#%g�/%EO��c�6����l��ZĐ�3z��K/����)�N�p"	��(�H�`)�W5�s����OT͝Oǎs��
M�?��$&�?f��:U0��8ӟznC�u:N�n[`��(�mHNކ�9�]�]��7�B<�*=Ʒmݬ���ڷo�zi����A�p~PzȘ*�gdT}�_��Z+�و���Ы��`^+�{'O�0J�\h�8��TT�Mu�H�ʽRU}'�zY����?���_�e��]	؇���%����t򓕮�ԫ[O�Ѷ��(��Ν;u�۪v�59���v��1̍f63�٤������Y����mT�:1������]޵Ls������U���v���_�d�R8�rF[�nÌ߫�J�̭>RS�v*���� Q�������*K:ffe!.6�J����]�N�L*Svq9������m�2��Uږ����۷��~�]���R����ft���;�-^��k���Æ�;vbʔ/зO�c6C��gb����|�z���#q֠Az-i�O�^�zhּ6m�^�e�Mz�}\_s-������6��u2;�$x�����BNN�I�d�����K.�Z�%yd^�#��n�Ն^3'��%k�r�U)}���^��u��]vN9i�Q�b��yr2>��s���d6�����mZ���O�܇gq����1��_,�"��u�֣e��
[�n�ƍ��mXY�֭u��(ڨ�^�nv�*��|#d	S�z������H���.���R� 'AIa�������������t�m6\~�e��/�q�:��ٰ=y^z�%t萄���G�)�L@1y��X��?�7��s���0{;�������`�1�Х��Qe
N+LtE�i�쟱{��>���٫�^~��ߊ �y���T@�a񬁕+WaŊ�8픓z\��������s�~��*cQ6@�&MФqc�h���:�����N~3u�	[yU�5��]�}�Νqɥ�`��qz&'+�&M������ȣ�e�i�l���{((��L&�hּ��'A��9���[q۱}�f�*���]wމvm����ٻ3�NG>���ckšO�����}'R �=$�����s����>uON�2����.\�_���Ԕ�أ�d/:��]�>�p�'�se6s����巽BL��:/l�
�W]}��6�[��e����+HHH��s"�ë얔m�*�?�̳ػ�[�z"��.��{�*w�R��ۯ�;��f����0u�T64`S�����|K/���ŤI��úw>ё����3�w��S8�����^ݗ�^���k ��r�ÙY���U0���;��2�UI=�S]�h�����z�I�YN�l2����~�m�a�S��p���؟��}N_��o����W�|�^�/��,^���dNt��7�|�.e�:ݎ^��?�|UZ����&m�'N���N9�J�/9�e+V���^Cf�� ({+JO�s�=͛5�B
$��ڧo�4�GX�1�=9/�8mޜ����W|e�Q���o�nW;g�uV��i��ЭÏ4�y�d����Ə:sJ"\݀7� ��*O��+/��6]���O�^<p?ڵi��	D ����3Ĩ��x��`����E�.]�>�Yg���y�υU_��[6���c�L%rmZ�:���j߇^��*�[�V�hѪ.��|]�
���O��UW_�y��!+Ӻs܌�CR�x��'sd�Lxz��^�cǎՙ~o��N���5ADd�^��j1���<�Kܒ%�ωe@p�v�����ª���n�{�X6d��a�oa��ŸM��SZ������6�I]6mقw�yWW��L���NJ�W_}���
�۞eY
��oT���*�;�����J4�0t�0�ya:�kW�DN��c�.<��p|�ŗ��l�$,,�^{-�w��`NU��s��_���V�z~~�|��G������n|���ҫ�ɧ��?{�j�v��|��hP�~���ccbi�?��}���3rM����t�SB7ٖQ��XRU7��0l�CؽSz�Z}A}����O=���'�����y��'�u�V��c^r9��,lܸ�~����5V�Ҭ����X�W<s }����}���~��3>��S��e%��_���}��GqҀ�^�&��Zi..Z�J*���7��/�p��	'���E�������{J��}��WGw��.:s�����q�
�����"G%_��Q����g��Y::{�ٺ�����w����<k�̾t�����z�T��n_���N�e�U�Zn	ݕ蒇L6q�嗫l�	��jއ��Ds~�	���;Z�j�~���G�����84i�1��:�K)\������{�`ٲ�X�d�.�oS9��Y�|��LO��1ϣm����}݄x�Y�իWc��%�J䤏��ٳ�f�\}�5�����!)Ig ��N:mڼ	ӿ��>�[6m.�WYN�l��?��^�`NUi����{���#��]z���eMM����q���~-[�@���}f��`��ǧ�->��l\���8ѵ{<��Cz\zM����j�ɢ֭�z���];q�}`��i�ԩ���9����ߥ�q�1��+�ak�r���6`�ZD����_�uz���F`�~�+odC��v�����٧vĨĠN|��)�H@�ǲT@Vw�����}�߳|�I'�ŗơO�^���ӫWO�5��s�^��[-Į�;0�����T/5+��e<�L#����g��)Y�p!�'o��᫆����`��0���@T��b-*(�y�ر};�y�/C@��z���xRe�'O���w��4j�	ut'���=m�r����زe�*I�.��{�F���SO���WMIg�}Ʃz+U��s�^�ru2���4���as��2q�i������G��T@/�#�蚢*\����$��z��c\r�˗-��Jg�[��d!�Çӽl��J���0���{�y1�Yt��9 7�9C�F���裏b��M�ԥ��k�v��~�=�UxD�c����<��Ư��M�5�SÇ��T����hеR*0H&2?� ���C�v�m�#遽i�z���˯��uהφ������3#��y�&x��q�X���d������u2
���X|�\������{�a���HP����z�Q^���ß�Rsx��e�^�6mZc��Q�q��ɖ��\+o�:W�L�ÿ��[q��w�I�FKdH��a�����ß��E���^)z����I���ʕ[�ҵ�J܆�63���&%ntlɽ�X}wF??J��ߞ�6�I/k�Mi�W��*�+�[^F���mݦ-�����
�\�����G��X����f
�))ػo��Ŧj�
��k����={b�ĉ��������H�|=�ze��W��SO;��s7�W���$��;g�^Fv�8���-2����U�9�s��:�	���K����ݺu�Čp�3���^��:�=��Ӻ���W^����aZ� X�E�ʻ���=22��q�}�����DU�]N_�#�=���{?v�H��A����HNN>f+\)���ˣ�����?��ުґCf�[�j5������G���!O�[OO[y�5W��s��OH�۽kL��:��x������,l.�H�M���O���O9�]w�^�F&�����^!N����5Z��W�������@�S�Z4���q��^��z�Ksp�	�>����*�e���G~y]lt4n��z=c�dοV���7��~?3��C���
�Q1�ر��Tw���6jРR���Ɏ�{��^�Z���bu<��qD��Is�|��F��}\(oi���9nӦ��=Opv�A�Н�����Ti����õ�K�L���m.���lݲUw�������HH�G�vmq�	'b��A�ӻ7��M�[�*Ty_҃]ޓ�������3�`�?ر}������К�fG�
�mU�\f�2dN:i �={+}��^�[�e�v:�zᜰ��Wmʾ���t�ֽ�LWr��I�V�!5r���֭[�kWu���Ǒ��S�Jur��=�d�%�v��!`��ʔ��{�,�w9���� ̋.׿Es�믎Ӷm�A�Hy�:��2r�sz����9?��ʕ+�����ɽe\
Oa���Eb�D����w.NS%r����Vi�٣�
n9% ��e��/=���tb릮yZڡ��/Sjk���W�\i^�fK��|���i�Oزy3���c��B��Zj3dTP||�����K����]],�J���մNG�s��gC�t�8�3t�;v"y{�^&TƖ������Y���HH�ڵ�PO���5k�\y�W]�fw���[�9��&w���ur�v�Y�F�N�e��Y%#=]�Ws�$*�j��^f��ر:w�W��#d����׫�	Z2���$�뮻���V"""W��+�I���>����QQQ~�ŕ��qϊ]�#>@���S�/�r�p��}e�#������-7�d��|b��+}lԵ�N����6m�ڵk�z��}�����lnn���bս.�=˒��ڵC'��v�{�Z�Z�
��s;��S��w�-kO�\�����S�|��/-�%� _��C�:�����Sqݮ

�����~%'�:u�ѨQC4i�T��1�2�S�
Ԭr�"�W݌�*ˣg����ِ\���5���@$��A)J%J2�Qj�����_��%�o��>�]� C��2w�zߒ ��� ��Ë����}�u�Dӓp�:�ʪ���qU{�o�VD�=��������"�LU}��qq�Q��)�/�I���&=ⳳ���ס�}��$�(:yHf˰�O�H/����r�;P�7��aUu<O�Tc��Q�9��k������΀^)f�K)C�\����b?�w,��#��L�im/��;�hݥ��8��|��8ގ)�ňp�z�����<��58��0K���0�~L��6�@;�\{u�yy�PM����Ni��f7����YB'""
f�S\�[y:�Q�ѝ8�)������^����3�-ӯ6�|v�#""
b���������(�ٝN��ֈ���7=S\�[�,HN�Љ������W~	]�9:����T:v���3M�r'"":�����,�Tn�7+�O"""
�K�ݯ8-%tFt""��d��m�::QPR1����DDDAKW��UBg�8""��e��˝Et""��U�:#:QP���U��8t""�`&U�~lU�?"""
F��ΈNDD�̊��3�)݆ι܉���;��~e/w""�����,�NDD�L��YB'""
jXm�m�DDD��"���������r�z�DDD՞S�r�5""����U*�}�k�r'""
ZR���VN�f,'""
fz�5?7eX'""
V�ߋ�0�'��,�U{�˧2�5?�r�܉�����m�r'""
b��U��DDDA��Nq�����(��~W�Q�b�;Q�Ǚ∈�B g�#""
~�C�˧2�+��^��DDDA���2DDD�ʏ�\�L��NDD���ΨNDD�����*w""���*w""�`�ʝ��(p�8""����kb=S+'�܉��B ;�U\m������K�p.w""�����\�DDD���X�U�DDDA��Q��LqDDD!����,DDD�*�˝m�DDDA�ɉe�������CgX'""
R�
T�Q�͉e���B��m�&�܉������6t"""
F�U��Gk��DDD����܉����
t�#""�`���WЉ����Dh�m��(񃈈���aT$��UBw8�HKK�!�p���� �`PS
Q���c�=�l����j���둓��ז�n��0l�C��Wæ�5�������]8
�������p����*�&6���e��-�8\yS~U��^�t1����h2�g�.��6��sDDDt�I��f4��&��� ""��JJ�:�烈���+UB7��͖n:�� ""��Hfsأ��ege�U;6�-3:::�^�n��������{�g��0=""�I&������K���;w$�Өqӻ<�t^^^/�4cTD��u�ƪ�3*8���c:1ϑ��g�#|���g��OF��x���$�����jժ�y�����W�<l��k�ŧ�O����;v����LP�F��]mn�G���E��l6�&m�v��0�æ�`ap�4�����rd��ϫXf��Ta���
�+����ſ�F�_JoWl����l�	�Q�k1׉x����󇢿B�8*�g�J����b{/���}����(:f��Qxn(���.u��{�`[�~���0T�.b�ҥ�{v�
/���G���NC�&M�T�^n7TWr�֬Y����[f�������=��ILl�o�Nɟ�f��MX�<[Q��}y�~����1�\4%�Y�wϮ�����,�{������vW��3K���yxv�c?%�l�Kb�R��\��W���)|q9��,q%��[����ĮK��}���n�a���{��_�]�r)�'�z_/)���N�l�b+��(�-6-�Y�b����J�-��ڨ�9��G�}{ΧԖ����t��pJ�e���%���-:�b�G�J�JM����.rџ�ݠ��:IϹ��\�������0̘�hg|BvIIs�����Saw���ʇ���G4�΅�Ϡ ?W?j"�gY"P������Ӑ@�p��ÐB�l�S�t8W pr�����T$u:�Õ��p?����w���&���\]$�b��$�o�^ܙ���kѾ����m6�����u�]o�ٽ�ً\t�Ÿ��[Bnn�;z��͸�λt"Q���N���on���'�<�������OOL�<O�EyUw�g��&�%�f�L������õ�Y�I�?\���u����hY<u���	S�,�;u):/��s�]6
ӛb�r�����
_��G���R�����̰�^����kc��4�ͦs�6Wy��-5�0�\�����6�]^cs[�e�._�CA��o��0RB�zHٿo��>�S?�� O�l٪UH��7�

���Vtx�is8t��4��J4�m�j��m�w��/�(5�_�O!_ega2�J%J��#��X�]<�g�إ{�i�'6�^�٧�Lexb�Y��Z�;�'���|��������Jl��2y�.�-�܌Ȉ��Zu#WD ��x���\���j�ژ��~̯s~Y߿}���E���[_a��p�2�mW|�ҥ�R��(�P�F�s+��(��/��(]�*��2�M��x�k�9��?ós�t�<�t�B�{��#�?=�Og^�{Tx6�k��F��'�����ܙ��r����w��=��M\�C���x�y0e[��|�}������vU��2��pU"R��Ɂ�
��c8�Զ��r���گ�S������r�Jt�ܹ�ug����e�,���o��� ����W;����"�#

�eF���e���سgZ6o�/S�T婌���o�c��-]:�mҬ�ks�u���'`��u���+AD,Щ���T<�$$$����J��ʬWr[�l���kt@�`.�;���*CS���f�^��?�>��t��6��{�Q0a@�2ڷh�ǞxR�����v��V&����a�?�`��A�>������_<��sػG��R���Jn߱ø���vh�] "
F�d�q�&�ݧw�_|�^�ڵ����������:��m;����x�駱j�
������f͚���/s�~y��6�w�� "
6�d)-��p|n���V���]*�J[�j5�nۊݺ�:ҝ���1f��y�l�i80ԫW��O>��/��Lꐄ�cǂ�(1���N�#:&f�
�y*�G��¦;�-Y��������λ����(�	N����h׾ݘO?�$%'�0���:Y�6�6m�ʔ���#���5*�M^n6����\s"��Q����{���K���@��0�=�Q��o��}�'�?�fM��;�"�`ŀN�.��b\{��6�#""|Wf��Ȫ/���K����^�jӎ.�bي�1b$��މ��\�����g��w�;��>�Y'>�G<"�`ƀN^����۴9�����U��Uv[�n����t@�$������ѣ�d�b�	�JtTTr��-�L�655/;DD�:y����`r�ڴi�Ff�*;ͫ��b�e8���Q���㭉1��o`5���W��k�.���� �n��O?"�`ǀN^}�~.����j���s�yyQ��q8�p�"���"*22��g��oLx��ٰ*�׊��ѭG��Np�����޻o���:`@'��M�ݺ�@TT�&e~^nS�v�U+Wb_J
Z4k�`�i75r����`��y���ϛ�����C��޻Љ��`@'��z�\vŕ��Ď�QQ۳27-���m۶bÆ�A�u��~w��b�vs�ݞݰA��+W,[8��G�Գ;n��jU��S߾}p�ק�<{�Z〭�%�:tK�.����`$����˒�����|�)�ߓ���mxi� "�N�ɧ����
���e�Ͷ��뻗�t`ѢE��ɑ�AՎ.'+��'�h7���]ٮ}����-c��� "���ɧ_�͚�D�:�W���g��^�j;iG߻oZ�h�`�״����p���n7���hܴ�����)_}��K�aԨ "�n�ɧ��.B�=l˚ի����Xt��۱~���	��SRS1z��^Ǜ6�,����\�պ�k0�|���K "��Щ\	uиq�ݪ�%=-�M�-����y��y�5�fϓv�I����v��:uz��/�ʱ���)�����b@�ru��I��9�U�a�Q�c�t`������Flt�1oG�v�7&L���[��#���7o�r�/?��y���ؽsN?�tUW�T.w�8�{�^�򚣠� �j�U+Wa�޽hӪ��x�#Gc��vsy6���s�͜�����O��3O���:c@�r͚5]��@|B����������e���ؾ�֭?f��<�`�E���_{�����/���w'OQuǀN�:��q�7�t:��/]�+++�n٭����v��:��(���y�EtL̎�mڌ�����0 ��Qv;"����_�z����/��?x�`�mLӡ�S���BlL�QoG�����7����`n���7i������3#����`ND!���Ҹi�rӍ��:���l��]y�e���ػwڴnu��MB�Ju\�j߻w,�����P��'�<��AC�1۶m��oL Q�`@'�<��Ø��iG_�J�9y+�Ihݹs'�o�p��������`���n��]�v�g�������q��_3�QHa@'�HǸ�I���Y����J,�v�e˖��AgU�9I0�/(��＋iS�I�?����#�7i����[2���ѳ[Q#��ÀN~��q=��t"۵�߅�2�3,�V3��ѳ��sƣ�4�g���k��΄U����s/�`J��]�v�Z<x߽ "
5���m����n94��S��`5��X�z��KA�U3�g��u6�y�w��˪vUX��]��Ν;��釙Y���� "
E����Cҹ�ٳW��av�� ?�2��x�M7VY@��JO�ر�������n�ڢeˑsf��)�a��_����Q(b@'�=8t(>��+ԩS{UDDxFA~^�	f��Ұt�2�y��*9��~�?|���0M'���e6���Mz��W�r�x���0⹧AD���o���Z�i���M��ѻ�23�Xm�׽*�G����ܹxy����̀uU���s���Mxz�3�5�[��ND!���ֿ�?^Ƥ����/������m�5�Wc_J
Z6o��K0߲u+F��m[7���m�ڷ����{�r���_���?Q(c@�
9����1))�s�n+m6���Hޖ�M�6,�K0����K/��彩�-�����4m�t��?��9���дi\q� "
u�T!��ɨ];			K#""rsrr"�n�jG_�l�vj@��0M|��g���>���U��a��~�ĩ���K/3���1�Y��Q���N2��3q�"22r}dT�����&V������%K�������J������k>^�"2��[���ۻ��*�<��?�����n4$kBGMk׭�bv�r�s'k7��f�v�Y�j^Rlk�Uh3#l[��dE!0�&"��*'8��e7��s�[�<|?3g8����w��9���L����ܶ�3� ���~�>*J���k������%��8m�F�Y�Dz򃴘מ���5k��\���G�|}[Ǎ�� ���T�|~�3y��' ���~�6�f��ҥm�3�t��_`�Kjj���ٳ
����Z:;e}F��������zWxDĎ�~����
� ?_�n� �pB��oK�zJ[`ƞp�m%��e����A�%-�-RRR"���;�jQ��y_v��]v�����	:���cGW@@���1��v:��Ç%.>ABCCK||}�m6k�����V)*:!]6�x�}:��W���Xa��MY+��f�����	�����Z�N��M*{��:�m������gŠ7T;v��J{{���_�|%M�&�w����74HRR��*+�^Q���ᆌ=|��W^����አc@�B�d��Sr?ʭ���0�Ӹ��*����	z_h1���ƍ�$���<��
�?w�?����/�k� W29�$��ϲ.%��*�~���p3J�su^ZZ*�Ϝ��s�ݷW�l�"6�U<͛�Un���o�ަ��RXX(��� �pE�1 ?��DG��M�'����X-���q6[�?^$֧�b4��禥�Dq�$'�H���t�����=>�Ճ���; �.\���x�ጠc@���f�~��������k�X:�=]Mk����-�q];��,)�k�d�	����N'QQQ{�WO�?c��v����+ �;��������L1u�
�k/{�$?w��������&[�n�?�#�}��Z!�!E3�e���hjn�m��  A� ����c�>bޙ�uZ���{ڨ���(��e2c�t���ҝ��'37HW�7ڢ�r�K�Z~:yrʮ���t�3R[^..  A� DDE�,0��_�Sl��~�����(/���EEb�Q����{W���%yM����Iϭv7��Fo׍��;�צ~x�;��Ȋ�� �_6w�,���Hxxx�ȑ#-�W�~�o�����XZ��亠����F6��Jj�:���/�Ӽ���ZdT�;�ߙ�>����%9�� �w:L�"uz\����-��dn�����R[S��o����)ٻ����i��%A����3��^{�g5���*� �C�1`�G����>Ѿ^��Ω����t��_� {��S�Iz}O���]��.�X����s����s�bc7�d��ߕ�P�1���y� ��:eF|��
h	)3��6���8m]��۷K��Y2g�,�8wN��$u_�WK/��i���_�Т7W�|�.�,~H  �"���ks��y��t����ߔNj��%=-]���$c}�=rD<=��]�GFF��=gv�ƍ�N����
 �cP^߲E��#gΜ)�;엺�����򤪲J*����Ԗ�u?o8j��֙�fnX���g�!�>yR  �t��%�n�Nʻ�|\z��t~�)�'��MR�e���i�L�]���훶lq���ɯ�<)  �:�d2ɒ����������ں��tz�~���w'L�X}Ͻ��ݺu���ݻD�d;A��tZ��J�:m��/>q����ā��%�GZܽ s�����j��u�̝@t�'��˧G���;�x�iʦ���X�V����`0J\|\ުU�v,8䊈���� �aC��?��{\Ǝ���?���b}�.�K��`4��W�Ǜ��j����pF�1$��^��:f츎�G������q���>��K:�n[xT��i�ؤ���[� �Cf�Ν��ޮm�r�������T����C�i�+��<�����-�  ����2˖,��/���s�J�ط���w���-���*<!!��]wߕ|������� }G�1���ِ������l�X��m�I=��������3>m�^9��ŕ���*/���  ���cH͙3Gv��-oeeɁ��"_�$�ݑ�]�Qn���z�;f�y��g�9��ӈ9 Aǐ[�x��d2���D����t:&8�UN���|�����`4�1��Eǋ���ʤ��V  C��8UZ*:�QBCB�'LL375�X::��lA:�����'wtp��u��wZ,�z�j1M�$ ��!���86ih��^��������dn�:V: `�:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
 �  (�� � � �:  
�O��Ր���    IEND�B`�PK
     uK\��EM  M  /   images/d3694a2e-5bba-40c3-8069-8db85c4c9209.png�PNG

   IHDR   d   d   p�T  TiCCPICC Profile  x�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D������d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c���Ԋ�_PY���Q���Tϼd=#CsP�CT�%���X�}�����ߍ�������k'BLÂ�A�����΂ĢD�33��10|Z����� |�'�8��,������z����j��N��������.j���p  !e�2���   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK 
     uK\���v� �                  cirkitFile.jsonPK 
     uK\                        ' jsons/PK 
     uK\����  ��               K jsons/user_defined.jsonPK 
     uK\                        � images/PK 
     uK\���)G )G /             �� images/ab296a80-256f-428c-a4e8-e177cdc61bff.pngPK 
     uK\���@  �@  /              images/c19b89aa-68d9-4a98-b509-123aa1ab0169.pngPK 
     uK\}�?`X X /             Z images/f6e2a5fb-4294-42a3-957b-9521668fdddb.pngPK 
     uK\�6�P�L  �L  /             �\ images/8fef4bdb-224a-4a07-91a3-222e74c30575.pngPK 
     uK\c0��T� T� /             � images/2b856d38-88e4-4759-8ee8-6b01c1d6fb9d.pngPK 
     uK\�����a  �a  /             �u images/9aa3d03b-0c22-4f62-98c6-f5f844a0dc7c.pngPK 
     uK\zn���1  �1  /             g� images/245bc533-66be-4bb3-b22a-43c007a581bd.pngPK 
     uK\qyဲ=  �=  /             �	 images/51c64262-e188-46ba-9658-f0d60e053320.pngPK 
     uK\��92\ 2\ /             �G images/7fb2f62e-2fb5-47b1-9980-8ec272392bae.pngPK 
     uK\y�ݥ�  �  /             �  images/2db9ecad-5c51-4c64-ac4d-4ae785eb4e5c.pngPK 
     uK\�$<�ʏ  ʏ  /             f)! images/cb669bd1-12cf-42eb-9243-39a8a80a0435.pngPK 
     uK\�T�'}  }  /             }�! images/1be29400-b52e-43b8-b531-83e2df2121b6.pngPK 
     uK\�}���) �) /             G�! images/146a6d58-0553-42c9-b8c7-03425202d69a.pngPK 
     uK\��C�I  I  /             ��" images/d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.pngPK 
     uK\��e e /             # images/48caf11c-09fe-45e4-9b76-5b0bfa123a56.pngPK 
     uK\���'  �'  /             }s( images/16bd2965-d7b7-4d97-b402-ac1747e7568c.pngPK 
     uK\�d)e�Y  �Y  /             ]�( images/ae99f124-1aaf-4a6e-8177-44087bd956ce.pngPK 
     uK\hyXe  e  /             ��( images/f7e3f572-2cc7-414e-8b58-58f37a09912a.pngPK 
     uK\P��ޮ  ޮ  /             5) images/98bdfb38-4044-46ed-976e-d2b53bff2879.pngPK 
     uK\_����<  �<  /             `�) images/1a257b89-3953-41e9-990a-6c271080df8c.pngPK 
     uK\G�BN��  ��  /             ��) images/d6a4f4f6-fe0f-43ac-893b-20774d3ea628.pngPK 
     uK\�4%2P  P  /             ��* images/c7b8e0ca-67ed-4237-9266-7527aa3ce92a.pngPK 
     uK\�|��*  *  /             1�* images/fe816bc3-a1ac-4496-aca2-7e46c72bb630.pngPK 
     uK\�|3�  �  /             ��* images/559c8cb2-c573-4147-bde4-a0b817dc20ed.pngPK 
     uK\ә�CJK  JK  /             ��* images/a0bdb5a7-9945-4126-87cb-dac9f24142ab.pngPK 
     uK\;b�i�  �  /             IH+ images/68998569-73de-4f26-b1b3-0b6c45f8499f.pngPK 
     uK\1y1�? �? /             =e+ images/a003a845-706b-4c0a-bac4-0f60a60b44e4.pngPK 
     uK\�l��P� P� /             R�. images/8a348e4e-00a9-420c-8c54-2da977db0968.pngPK 
     uK\+B�<r <r /             �P1 images/9d915518-60ad-41a3-8ee2-5a1cc2d88e80.pngPK 
     uK\z?�A�  �  /             x�2 images/a652ce68-b987-46e6-8408-d5645582d4d7.pngPK 
     uK\�u`�) �) /             G�2 images/a27a8979-5023-407e-b6b7-e8628572ca80.pngPK 
     uK\QQΒ�!  �!  /              5 images/5441ee9b-7343-4a92-92bb-e3ea11bfaf7c.pngPK 
     uK\J�-E�I �I /             A*5 images/10aa979f-dd42-43c7-9c2f-b8fbfcd42f21.pngPK 
     uK\>B�	  	  /             ot7 images/687e948c-dc0a-4fdc-b588-e952ae529de1.pngPK 
     uK\�c��f  �f  /             �}7 images/c88b2895-5e8b-4a57-9f9a-b80dd50058b1.pngPK 
     uK\��EM  M  /             ��7 images/d3694a2e-5bba-40c3-8069-8db85c4c9209.pngPK    ( ( �  ��7   